

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771;

  BUF_X1 U376 ( .A(n643), .Z(n355) );
  XNOR2_X1 U377 ( .A(n397), .B(KEYINPUT71), .ZN(n595) );
  OR2_X1 U378 ( .A1(n635), .A2(G902), .ZN(n482) );
  XNOR2_X1 U379 ( .A(n527), .B(n425), .ZN(n496) );
  XNOR2_X1 U380 ( .A(n366), .B(G143), .ZN(n527) );
  XNOR2_X1 U381 ( .A(G128), .B(KEYINPUT84), .ZN(n366) );
  XNOR2_X2 U382 ( .A(n354), .B(n431), .ZN(n430) );
  NAND2_X2 U383 ( .A1(n626), .A2(n625), .ZN(n354) );
  NOR2_X1 U384 ( .A1(G953), .A2(G237), .ZN(n510) );
  XNOR2_X1 U385 ( .A(n543), .B(n542), .ZN(n677) );
  INV_X1 U386 ( .A(n536), .ZN(n584) );
  AND2_X2 U387 ( .A1(n361), .A2(n591), .ZN(n598) );
  XNOR2_X2 U388 ( .A(n567), .B(KEYINPUT45), .ZN(n750) );
  NOR2_X2 U389 ( .A1(n643), .A2(n770), .ZN(n593) );
  XNOR2_X2 U390 ( .A(n428), .B(n427), .ZN(n770) );
  XNOR2_X2 U391 ( .A(n755), .B(n458), .ZN(n730) );
  XNOR2_X2 U392 ( .A(n496), .B(n451), .ZN(n755) );
  XNOR2_X1 U393 ( .A(n508), .B(KEYINPUT0), .ZN(n534) );
  INV_X1 U394 ( .A(n623), .ZN(n607) );
  NOR2_X1 U395 ( .A1(n552), .A2(n551), .ZN(n555) );
  XNOR2_X1 U396 ( .A(n541), .B(n399), .ZN(n704) );
  NOR2_X1 U397 ( .A1(n534), .A2(n357), .ZN(n535) );
  XNOR2_X1 U398 ( .A(n415), .B(n520), .ZN(n408) );
  NAND2_X2 U399 ( .A1(n371), .A2(n367), .ZN(n424) );
  XNOR2_X1 U400 ( .A(n646), .B(n645), .ZN(n647) );
  AND2_X1 U401 ( .A1(n373), .A2(n372), .ZN(n371) );
  XNOR2_X1 U402 ( .A(n413), .B(G104), .ZN(n514) );
  XNOR2_X1 U403 ( .A(n426), .B(KEYINPUT64), .ZN(n425) );
  XNOR2_X1 U404 ( .A(n412), .B(G107), .ZN(n525) );
  INV_X2 U405 ( .A(G953), .ZN(n761) );
  XNOR2_X1 U406 ( .A(KEYINPUT70), .B(G131), .ZN(n512) );
  XNOR2_X1 U407 ( .A(KEYINPUT4), .B(G146), .ZN(n426) );
  XNOR2_X1 U408 ( .A(KEYINPUT15), .B(G902), .ZN(n629) );
  NOR2_X1 U409 ( .A1(n592), .A2(n672), .ZN(n429) );
  AND2_X2 U410 ( .A1(n615), .A2(n767), .ZN(n616) );
  XNOR2_X2 U411 ( .A(n424), .B(n461), .ZN(n693) );
  INV_X1 U412 ( .A(G116), .ZN(n412) );
  INV_X1 U413 ( .A(G137), .ZN(n449) );
  XNOR2_X1 U414 ( .A(n423), .B(KEYINPUT77), .ZN(n410) );
  NAND2_X1 U415 ( .A1(n393), .A2(n374), .ZN(n423) );
  NAND2_X1 U416 ( .A1(n730), .A2(n460), .ZN(n373) );
  XNOR2_X1 U417 ( .A(n500), .B(n499), .ZN(n744) );
  XNOR2_X1 U418 ( .A(n411), .B(n358), .ZN(n500) );
  NOR2_X1 U419 ( .A1(n614), .A2(n613), .ZN(n395) );
  XNOR2_X1 U420 ( .A(n470), .B(KEYINPUT20), .ZN(n472) );
  NOR2_X1 U421 ( .A1(n771), .A2(n644), .ZN(n562) );
  AND2_X1 U422 ( .A1(n586), .A2(n585), .ZN(n587) );
  INV_X1 U423 ( .A(n629), .ZN(n389) );
  INV_X1 U424 ( .A(n460), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n574), .B(KEYINPUT6), .ZN(n594) );
  INV_X1 U426 ( .A(KEYINPUT104), .ZN(n521) );
  AND2_X1 U427 ( .A1(n526), .A2(G217), .ZN(n422) );
  XOR2_X1 U428 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n523) );
  INV_X1 U429 ( .A(G122), .ZN(n413) );
  XOR2_X1 U430 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n516) );
  XNOR2_X1 U431 ( .A(G143), .B(G113), .ZN(n515) );
  AND2_X1 U432 ( .A1(n633), .A2(KEYINPUT65), .ZN(n385) );
  NAND2_X1 U433 ( .A1(n378), .A2(n377), .ZN(n380) );
  NAND2_X1 U434 ( .A1(KEYINPUT2), .A2(n381), .ZN(n377) );
  INV_X1 U435 ( .A(n388), .ZN(n382) );
  XNOR2_X1 U436 ( .A(n744), .B(n501), .ZN(n653) );
  XNOR2_X1 U437 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U438 ( .A(n580), .B(n579), .ZN(n592) );
  XNOR2_X1 U439 ( .A(n392), .B(n391), .ZN(n438) );
  INV_X1 U440 ( .A(KEYINPUT36), .ZN(n391) );
  INV_X1 U441 ( .A(G478), .ZN(n416) );
  NAND2_X1 U442 ( .A1(n646), .A2(n369), .ZN(n415) );
  NAND2_X1 U443 ( .A1(n417), .A2(n376), .ZN(n694) );
  NAND2_X1 U444 ( .A1(G234), .A2(G237), .ZN(n485) );
  XNOR2_X1 U445 ( .A(n433), .B(n473), .ZN(n695) );
  NAND2_X1 U446 ( .A1(n472), .A2(G221), .ZN(n433) );
  XNOR2_X1 U447 ( .A(G119), .B(G116), .ZN(n475) );
  XNOR2_X1 U448 ( .A(KEYINPUT3), .B(G113), .ZN(n479) );
  XNOR2_X1 U449 ( .A(n514), .B(n525), .ZN(n411) );
  INV_X1 U450 ( .A(KEYINPUT65), .ZN(n381) );
  XOR2_X1 U451 ( .A(KEYINPUT80), .B(G140), .Z(n455) );
  XNOR2_X1 U452 ( .A(G110), .B(G107), .ZN(n454) );
  XOR2_X1 U453 ( .A(G101), .B(G104), .Z(n453) );
  INV_X1 U454 ( .A(G125), .ZN(n492) );
  XOR2_X1 U455 ( .A(KEYINPUT18), .B(KEYINPUT81), .Z(n491) );
  INV_X1 U456 ( .A(KEYINPUT90), .ZN(n431) );
  AND2_X1 U457 ( .A1(n550), .A2(n549), .ZN(n561) );
  BUF_X1 U458 ( .A(n691), .Z(n714) );
  OR2_X1 U459 ( .A1(G237), .A2(G902), .ZN(n503) );
  AND2_X1 U460 ( .A1(n583), .A2(n596), .ZN(n688) );
  XNOR2_X1 U461 ( .A(n445), .B(n444), .ZN(n409) );
  NOR2_X1 U462 ( .A1(n594), .A2(n672), .ZN(n446) );
  XNOR2_X1 U463 ( .A(n695), .B(n432), .ZN(n532) );
  INV_X1 U464 ( .A(KEYINPUT100), .ZN(n432) );
  XNOR2_X1 U465 ( .A(n441), .B(n440), .ZN(n439) );
  XNOR2_X1 U466 ( .A(n471), .B(KEYINPUT98), .ZN(n440) );
  XNOR2_X1 U467 ( .A(G128), .B(G137), .ZN(n462) );
  AND2_X1 U468 ( .A1(n409), .A2(n596), .ZN(n418) );
  AND2_X1 U469 ( .A1(n405), .A2(n528), .ZN(n402) );
  INV_X1 U470 ( .A(KEYINPUT102), .ZN(n399) );
  OR2_X1 U471 ( .A1(n730), .A2(n368), .ZN(n367) );
  NAND2_X1 U472 ( .A1(n370), .A2(n369), .ZN(n368) );
  XNOR2_X1 U473 ( .A(n527), .B(n524), .ZN(n419) );
  XNOR2_X1 U474 ( .A(n422), .B(n421), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n519), .B(n518), .ZN(n646) );
  NAND2_X2 U476 ( .A1(n383), .A2(n379), .ZN(n736) );
  NAND2_X1 U477 ( .A1(n382), .A2(n380), .ZN(n379) );
  XNOR2_X1 U478 ( .A(n653), .B(n652), .ZN(n654) );
  AND2_X1 U479 ( .A1(n638), .A2(G953), .ZN(n743) );
  INV_X1 U480 ( .A(KEYINPUT42), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n429), .B(KEYINPUT40), .ZN(n643) );
  INV_X1 U482 ( .A(KEYINPUT111), .ZN(n435) );
  INV_X1 U483 ( .A(n597), .ZN(n437) );
  XNOR2_X1 U484 ( .A(n553), .B(KEYINPUT83), .ZN(n554) );
  NAND2_X1 U485 ( .A1(n407), .A2(n538), .ZN(n667) );
  INV_X1 U486 ( .A(n672), .ZN(n674) );
  NAND2_X1 U487 ( .A1(n408), .A2(n539), .ZN(n672) );
  INV_X1 U488 ( .A(n584), .ZN(n588) );
  OR2_X1 U489 ( .A1(n737), .A2(G902), .ZN(n356) );
  XOR2_X1 U490 ( .A(KEYINPUT105), .B(n533), .Z(n357) );
  XNOR2_X1 U491 ( .A(KEYINPUT16), .B(KEYINPUT75), .ZN(n358) );
  XNOR2_X1 U492 ( .A(n356), .B(n416), .ZN(n539) );
  XOR2_X1 U493 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n359) );
  XOR2_X1 U494 ( .A(G125), .B(G140), .Z(n360) );
  XOR2_X1 U495 ( .A(n424), .B(KEYINPUT108), .Z(n361) );
  AND2_X1 U496 ( .A1(n631), .A2(n381), .ZN(n362) );
  AND2_X1 U497 ( .A1(n623), .A2(n596), .ZN(n363) );
  AND2_X1 U498 ( .A1(G210), .A2(n503), .ZN(n364) );
  NOR2_X1 U499 ( .A1(n424), .A2(n573), .ZN(n365) );
  XNOR2_X1 U500 ( .A(n436), .B(n435), .ZN(n767) );
  INV_X1 U501 ( .A(G902), .ZN(n369) );
  INV_X1 U502 ( .A(KEYINPUT2), .ZN(n633) );
  AND2_X2 U503 ( .A1(n386), .A2(n384), .ZN(n383) );
  NAND2_X2 U504 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U505 ( .A1(n460), .A2(G902), .ZN(n372) );
  INV_X1 U506 ( .A(n693), .ZN(n374) );
  AND2_X1 U507 ( .A1(n393), .A2(n375), .ZN(n545) );
  INV_X1 U508 ( .A(n424), .ZN(n375) );
  INV_X1 U509 ( .A(n393), .ZN(n376) );
  XNOR2_X2 U510 ( .A(n396), .B(KEYINPUT68), .ZN(n393) );
  NAND2_X1 U511 ( .A1(n632), .A2(n631), .ZN(n387) );
  NAND2_X1 U512 ( .A1(n632), .A2(n362), .ZN(n378) );
  NAND2_X1 U513 ( .A1(n387), .A2(n385), .ZN(n384) );
  NAND2_X1 U514 ( .A1(n388), .A2(KEYINPUT65), .ZN(n386) );
  OR2_X2 U515 ( .A1(n750), .A2(n628), .ZN(n390) );
  INV_X1 U516 ( .A(n390), .ZN(n682) );
  XNOR2_X2 U517 ( .A(n607), .B(KEYINPUT38), .ZN(n583) );
  XNOR2_X1 U518 ( .A(n517), .B(n447), .ZN(n519) );
  NAND2_X1 U519 ( .A1(n595), .A2(n446), .ZN(n445) );
  NAND2_X1 U520 ( .A1(n409), .A2(n363), .ZN(n392) );
  XNOR2_X1 U521 ( .A(n420), .B(n419), .ZN(n737) );
  XNOR2_X1 U522 ( .A(n555), .B(n554), .ZN(n771) );
  INV_X1 U523 ( .A(n539), .ZN(n538) );
  NAND2_X1 U524 ( .A1(n393), .A2(n365), .ZN(n577) );
  AND2_X2 U525 ( .A1(n395), .A2(n394), .ZN(n615) );
  NAND2_X1 U526 ( .A1(n602), .A2(KEYINPUT47), .ZN(n394) );
  INV_X2 U527 ( .A(G119), .ZN(n434) );
  NOR2_X2 U528 ( .A1(n536), .A2(n474), .ZN(n396) );
  XNOR2_X2 U529 ( .A(n482), .B(G472), .ZN(n574) );
  NAND2_X1 U530 ( .A1(n588), .A2(n587), .ZN(n397) );
  NAND2_X1 U531 ( .A1(n623), .A2(n596), .ZN(n506) );
  XNOR2_X2 U532 ( .A(n502), .B(n364), .ZN(n623) );
  NAND2_X1 U533 ( .A1(n410), .A2(n483), .ZN(n484) );
  NAND2_X2 U534 ( .A1(n398), .A2(n403), .ZN(n529) );
  AND2_X2 U535 ( .A1(n401), .A2(n402), .ZN(n398) );
  NAND2_X1 U536 ( .A1(n704), .A2(n544), .ZN(n542) );
  NAND2_X1 U537 ( .A1(n691), .A2(n400), .ZN(n401) );
  AND2_X1 U538 ( .A1(n544), .A2(n509), .ZN(n400) );
  XNOR2_X2 U539 ( .A(n484), .B(KEYINPUT33), .ZN(n691) );
  NAND2_X1 U540 ( .A1(n404), .A2(n406), .ZN(n403) );
  INV_X1 U541 ( .A(n691), .ZN(n404) );
  NAND2_X1 U542 ( .A1(n534), .A2(n406), .ZN(n405) );
  INV_X1 U543 ( .A(n509), .ZN(n406) );
  NOR2_X1 U544 ( .A1(n408), .A2(n538), .ZN(n685) );
  INV_X1 U545 ( .A(n408), .ZN(n407) );
  NAND2_X1 U546 ( .A1(n538), .A2(n408), .ZN(n606) );
  NAND2_X1 U547 ( .A1(n410), .A2(n700), .ZN(n541) );
  INV_X1 U548 ( .A(n583), .ZN(n684) );
  XNOR2_X2 U549 ( .A(n414), .B(n448), .ZN(n715) );
  NAND2_X1 U550 ( .A1(n688), .A2(n685), .ZN(n414) );
  NAND2_X1 U551 ( .A1(n418), .A2(n417), .ZN(n622) );
  INV_X1 U552 ( .A(n620), .ZN(n417) );
  XNOR2_X1 U553 ( .A(n525), .B(n523), .ZN(n421) );
  XNOR2_X1 U554 ( .A(n498), .B(n462), .ZN(n465) );
  NOR2_X2 U555 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U556 ( .A1(n715), .A2(n598), .ZN(n428) );
  NAND2_X1 U557 ( .A1(n430), .A2(n765), .ZN(n720) );
  NAND2_X1 U558 ( .A1(n430), .A2(n721), .ZN(n628) );
  XNOR2_X2 U559 ( .A(n434), .B(G110), .ZN(n498) );
  NAND2_X1 U560 ( .A1(n438), .A2(n437), .ZN(n436) );
  XNOR2_X2 U561 ( .A(n442), .B(n439), .ZN(n536) );
  NAND2_X1 U562 ( .A1(n472), .A2(G217), .ZN(n441) );
  OR2_X2 U563 ( .A1(n740), .A2(G902), .ZN(n442) );
  XNOR2_X1 U564 ( .A(n443), .B(n518), .ZN(n740) );
  XNOR2_X1 U565 ( .A(n469), .B(n468), .ZN(n443) );
  INV_X1 U566 ( .A(KEYINPUT106), .ZN(n444) );
  BUF_X1 U567 ( .A(n720), .Z(n760) );
  XOR2_X1 U568 ( .A(n516), .B(n515), .Z(n447) );
  XNOR2_X1 U569 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n448) );
  INV_X1 U570 ( .A(KEYINPUT78), .ZN(n630) );
  XNOR2_X1 U571 ( .A(n492), .B(KEYINPUT17), .ZN(n493) );
  XNOR2_X1 U572 ( .A(n522), .B(n521), .ZN(n524) );
  INV_X1 U573 ( .A(n534), .ZN(n544) );
  INV_X1 U574 ( .A(KEYINPUT32), .ZN(n553) );
  XNOR2_X1 U575 ( .A(n449), .B(G134), .ZN(n450) );
  XNOR2_X1 U576 ( .A(n512), .B(n450), .ZN(n451) );
  NAND2_X1 U577 ( .A1(G227), .A2(n761), .ZN(n452) );
  XNOR2_X1 U578 ( .A(n453), .B(n452), .ZN(n457) );
  XNOR2_X1 U579 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U580 ( .A(n457), .B(n456), .ZN(n458) );
  INV_X1 U581 ( .A(KEYINPUT72), .ZN(n459) );
  XNOR2_X1 U582 ( .A(n459), .B(G469), .ZN(n460) );
  XNOR2_X1 U583 ( .A(KEYINPUT1), .B(KEYINPUT66), .ZN(n461) );
  XOR2_X1 U584 ( .A(KEYINPUT97), .B(KEYINPUT73), .Z(n463) );
  XNOR2_X1 U585 ( .A(n463), .B(n359), .ZN(n464) );
  XNOR2_X1 U586 ( .A(n465), .B(n464), .ZN(n469) );
  NAND2_X1 U587 ( .A1(n761), .A2(G234), .ZN(n467) );
  XNOR2_X1 U588 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n466) );
  XNOR2_X1 U589 ( .A(n467), .B(n466), .ZN(n526) );
  NAND2_X1 U590 ( .A1(G221), .A2(n526), .ZN(n468) );
  XNOR2_X1 U591 ( .A(KEYINPUT10), .B(n360), .ZN(n756) );
  XNOR2_X1 U592 ( .A(G146), .B(n756), .ZN(n518) );
  XOR2_X1 U593 ( .A(KEYINPUT25), .B(KEYINPUT79), .Z(n471) );
  NAND2_X1 U594 ( .A1(G234), .A2(n629), .ZN(n470) );
  XOR2_X1 U595 ( .A(KEYINPUT99), .B(KEYINPUT21), .Z(n473) );
  INV_X1 U596 ( .A(n532), .ZN(n474) );
  NAND2_X1 U597 ( .A1(n510), .A2(G210), .ZN(n476) );
  XNOR2_X1 U598 ( .A(n476), .B(n475), .ZN(n478) );
  XNOR2_X1 U599 ( .A(KEYINPUT101), .B(KEYINPUT5), .ZN(n477) );
  XNOR2_X1 U600 ( .A(n478), .B(n477), .ZN(n480) );
  XNOR2_X1 U601 ( .A(n479), .B(G101), .ZN(n497) );
  XNOR2_X1 U602 ( .A(n480), .B(n497), .ZN(n481) );
  XNOR2_X1 U603 ( .A(n755), .B(n481), .ZN(n635) );
  INV_X1 U604 ( .A(n594), .ZN(n483) );
  NOR2_X1 U605 ( .A1(G898), .A2(n761), .ZN(n745) );
  XNOR2_X1 U606 ( .A(KEYINPUT14), .B(n485), .ZN(n487) );
  NAND2_X1 U607 ( .A1(G902), .A2(n487), .ZN(n568) );
  INV_X1 U608 ( .A(n568), .ZN(n486) );
  NAND2_X1 U609 ( .A1(n745), .A2(n486), .ZN(n489) );
  NAND2_X1 U610 ( .A1(G952), .A2(n487), .ZN(n713) );
  NOR2_X1 U611 ( .A1(G953), .A2(n713), .ZN(n488) );
  XOR2_X1 U612 ( .A(KEYINPUT96), .B(n488), .Z(n571) );
  NAND2_X1 U613 ( .A1(n489), .A2(n571), .ZN(n507) );
  NAND2_X1 U614 ( .A1(G224), .A2(n761), .ZN(n490) );
  XNOR2_X1 U615 ( .A(n491), .B(n490), .ZN(n494) );
  XNOR2_X1 U616 ( .A(n496), .B(n495), .ZN(n501) );
  XNOR2_X1 U617 ( .A(n498), .B(n497), .ZN(n499) );
  NAND2_X1 U618 ( .A1(n653), .A2(n629), .ZN(n502) );
  NAND2_X1 U619 ( .A1(G214), .A2(n503), .ZN(n505) );
  INV_X1 U620 ( .A(KEYINPUT95), .ZN(n504) );
  XNOR2_X1 U621 ( .A(n505), .B(n504), .ZN(n596) );
  XNOR2_X1 U622 ( .A(n506), .B(KEYINPUT19), .ZN(n599) );
  NAND2_X1 U623 ( .A1(n507), .A2(n599), .ZN(n508) );
  XOR2_X1 U624 ( .A(KEYINPUT34), .B(KEYINPUT82), .Z(n509) );
  NAND2_X1 U625 ( .A1(n510), .A2(G214), .ZN(n511) );
  XNOR2_X1 U626 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U627 ( .A(n514), .B(n513), .ZN(n517) );
  XOR2_X1 U628 ( .A(KEYINPUT13), .B(G475), .Z(n520) );
  XNOR2_X1 U629 ( .A(G134), .B(G122), .ZN(n522) );
  INV_X1 U630 ( .A(n606), .ZN(n528) );
  XNOR2_X2 U631 ( .A(n529), .B(KEYINPUT35), .ZN(n769) );
  NAND2_X1 U632 ( .A1(n769), .A2(KEYINPUT44), .ZN(n531) );
  INV_X1 U633 ( .A(KEYINPUT92), .ZN(n530) );
  NAND2_X1 U634 ( .A1(n531), .A2(n530), .ZN(n550) );
  NAND2_X1 U635 ( .A1(n685), .A2(n532), .ZN(n533) );
  XNOR2_X1 U636 ( .A(n535), .B(KEYINPUT22), .ZN(n556) );
  NAND2_X1 U637 ( .A1(n556), .A2(n594), .ZN(n552) );
  NAND2_X1 U638 ( .A1(n584), .A2(n417), .ZN(n537) );
  NOR2_X1 U639 ( .A1(n552), .A2(n537), .ZN(n659) );
  NAND2_X1 U640 ( .A1(n672), .A2(n667), .ZN(n687) );
  INV_X1 U641 ( .A(n687), .ZN(n610) );
  XOR2_X1 U642 ( .A(KEYINPUT103), .B(KEYINPUT31), .Z(n543) );
  INV_X1 U643 ( .A(n574), .ZN(n540) );
  INV_X1 U644 ( .A(n540), .ZN(n700) );
  NAND2_X1 U645 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U646 ( .A1(n546), .A2(n700), .ZN(n663) );
  NOR2_X1 U647 ( .A1(n677), .A2(n663), .ZN(n547) );
  NOR2_X1 U648 ( .A1(n610), .A2(n547), .ZN(n548) );
  NOR2_X1 U649 ( .A1(n659), .A2(n548), .ZN(n549) );
  NOR2_X1 U650 ( .A1(n769), .A2(KEYINPUT44), .ZN(n559) );
  INV_X1 U651 ( .A(n693), .ZN(n620) );
  XOR2_X1 U652 ( .A(KEYINPUT94), .B(n620), .Z(n597) );
  OR2_X1 U653 ( .A1(n584), .A2(n597), .ZN(n551) );
  NOR2_X1 U654 ( .A1(n584), .A2(n620), .ZN(n557) );
  NAND2_X1 U655 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U656 ( .A1(n558), .A2(n700), .ZN(n644) );
  NAND2_X1 U657 ( .A1(n559), .A2(n562), .ZN(n560) );
  NAND2_X1 U658 ( .A1(n561), .A2(n560), .ZN(n566) );
  NAND2_X1 U659 ( .A1(n769), .A2(KEYINPUT92), .ZN(n563) );
  NAND2_X1 U660 ( .A1(n563), .A2(n562), .ZN(n564) );
  AND2_X1 U661 ( .A1(n564), .A2(KEYINPUT44), .ZN(n565) );
  NOR2_X1 U662 ( .A1(G900), .A2(n568), .ZN(n569) );
  NAND2_X1 U663 ( .A1(n569), .A2(G953), .ZN(n570) );
  AND2_X1 U664 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U665 ( .A(n572), .B(KEYINPUT85), .ZN(n586) );
  INV_X1 U666 ( .A(n586), .ZN(n573) );
  NAND2_X1 U667 ( .A1(n574), .A2(n596), .ZN(n575) );
  XNOR2_X1 U668 ( .A(n575), .B(KEYINPUT30), .ZN(n576) );
  NOR2_X2 U669 ( .A1(n577), .A2(n576), .ZN(n609) );
  NAND2_X1 U670 ( .A1(n609), .A2(n583), .ZN(n580) );
  INV_X1 U671 ( .A(KEYINPUT74), .ZN(n578) );
  XNOR2_X1 U672 ( .A(n578), .B(KEYINPUT39), .ZN(n579) );
  OR2_X1 U673 ( .A1(n592), .A2(n667), .ZN(n581) );
  XNOR2_X1 U674 ( .A(n581), .B(KEYINPUT112), .ZN(n765) );
  NAND2_X1 U675 ( .A1(KEYINPUT2), .A2(n765), .ZN(n582) );
  XOR2_X1 U676 ( .A(KEYINPUT86), .B(n582), .Z(n721) );
  INV_X1 U677 ( .A(n596), .ZN(n683) );
  INV_X1 U678 ( .A(n695), .ZN(n585) );
  NAND2_X1 U679 ( .A1(n595), .A2(n700), .ZN(n590) );
  XNOR2_X1 U680 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n589) );
  XNOR2_X1 U681 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U682 ( .A(n593), .B(KEYINPUT46), .ZN(n617) );
  NAND2_X1 U683 ( .A1(n599), .A2(n598), .ZN(n671) );
  NOR2_X1 U684 ( .A1(KEYINPUT89), .A2(n687), .ZN(n600) );
  NOR2_X1 U685 ( .A1(n671), .A2(n600), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n601), .A2(KEYINPUT76), .ZN(n602) );
  XOR2_X1 U687 ( .A(KEYINPUT76), .B(n610), .Z(n604) );
  INV_X1 U688 ( .A(KEYINPUT47), .ZN(n603) );
  NAND2_X1 U689 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U690 ( .A1(n671), .A2(n605), .ZN(n614) );
  NOR2_X1 U691 ( .A1(n607), .A2(n606), .ZN(n608) );
  NAND2_X1 U692 ( .A1(n609), .A2(n608), .ZN(n642) );
  NAND2_X1 U693 ( .A1(KEYINPUT47), .A2(n610), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n611), .A2(KEYINPUT89), .ZN(n612) );
  NAND2_X1 U695 ( .A1(n642), .A2(n612), .ZN(n613) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n619) );
  XNOR2_X1 U697 ( .A(KEYINPUT91), .B(KEYINPUT48), .ZN(n618) );
  XNOR2_X1 U698 ( .A(n619), .B(n618), .ZN(n626) );
  XNOR2_X1 U699 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n621) );
  XNOR2_X1 U700 ( .A(n622), .B(n621), .ZN(n624) );
  NOR2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n679) );
  INV_X1 U702 ( .A(n679), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n720), .B(n630), .ZN(n632) );
  INV_X1 U704 ( .A(n750), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n736), .A2(G472), .ZN(n637) );
  XOR2_X1 U706 ( .A(KEYINPUT93), .B(KEYINPUT62), .Z(n634) );
  XNOR2_X1 U707 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n637), .B(n636), .ZN(n639) );
  INV_X1 U709 ( .A(G952), .ZN(n638) );
  NOR2_X2 U710 ( .A1(n639), .A2(n743), .ZN(n641) );
  INV_X1 U711 ( .A(KEYINPUT63), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n641), .B(n640), .ZN(G57) );
  XNOR2_X1 U713 ( .A(n642), .B(G143), .ZN(G45) );
  XOR2_X1 U714 ( .A(n355), .B(G131), .Z(G33) );
  XOR2_X1 U715 ( .A(G110), .B(n644), .Z(G12) );
  NAND2_X1 U716 ( .A1(n736), .A2(G475), .ZN(n648) );
  XOR2_X1 U717 ( .A(KEYINPUT67), .B(KEYINPUT59), .Z(n645) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(n649) );
  NOR2_X2 U719 ( .A1(n649), .A2(n743), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n650), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U721 ( .A1(n736), .A2(G210), .ZN(n655) );
  XNOR2_X1 U722 ( .A(KEYINPUT87), .B(KEYINPUT54), .ZN(n651) );
  XOR2_X1 U723 ( .A(n651), .B(KEYINPUT55), .Z(n652) );
  XNOR2_X1 U724 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X2 U725 ( .A1(n656), .A2(n743), .ZN(n658) );
  XNOR2_X1 U726 ( .A(KEYINPUT124), .B(KEYINPUT56), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n658), .B(n657), .ZN(G51) );
  XOR2_X1 U728 ( .A(G101), .B(n659), .Z(G3) );
  XOR2_X1 U729 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n661) );
  NAND2_X1 U730 ( .A1(n663), .A2(n674), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U732 ( .A(G104), .B(n662), .ZN(G6) );
  XOR2_X1 U733 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n665) );
  INV_X1 U734 ( .A(n667), .ZN(n676) );
  NAND2_X1 U735 ( .A1(n663), .A2(n676), .ZN(n664) );
  XNOR2_X1 U736 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U737 ( .A(G107), .B(n666), .ZN(G9) );
  NOR2_X1 U738 ( .A1(n667), .A2(n671), .ZN(n669) );
  XNOR2_X1 U739 ( .A(KEYINPUT115), .B(KEYINPUT29), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n669), .B(n668), .ZN(n670) );
  XOR2_X1 U741 ( .A(G128), .B(n670), .Z(G30) );
  NOR2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U743 ( .A(G146), .B(n673), .Z(G48) );
  NAND2_X1 U744 ( .A1(n677), .A2(n674), .ZN(n675) );
  XNOR2_X1 U745 ( .A(n675), .B(G113), .ZN(G15) );
  NAND2_X1 U746 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n678), .B(G116), .ZN(G18) );
  XNOR2_X1 U748 ( .A(G140), .B(n679), .ZN(n680) );
  XNOR2_X1 U749 ( .A(n680), .B(KEYINPUT117), .ZN(G42) );
  XOR2_X1 U750 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n681) );
  NOR2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n727) );
  NAND2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n686) );
  NAND2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n690) );
  NAND2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n692) );
  NAND2_X1 U756 ( .A1(n692), .A2(n714), .ZN(n709) );
  XNOR2_X1 U757 ( .A(KEYINPUT50), .B(n694), .ZN(n699) );
  XOR2_X1 U758 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n697) );
  NAND2_X1 U759 ( .A1(n695), .A2(n588), .ZN(n696) );
  XNOR2_X1 U760 ( .A(n697), .B(n696), .ZN(n698) );
  NAND2_X1 U761 ( .A1(n699), .A2(n698), .ZN(n701) );
  NOR2_X1 U762 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U763 ( .A(KEYINPUT119), .B(n702), .Z(n703) );
  NOR2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U765 ( .A(KEYINPUT120), .B(n705), .ZN(n706) );
  XNOR2_X1 U766 ( .A(n706), .B(KEYINPUT51), .ZN(n707) );
  NAND2_X1 U767 ( .A1(n707), .A2(n715), .ZN(n708) );
  NAND2_X1 U768 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U769 ( .A(n710), .B(KEYINPUT121), .ZN(n711) );
  XNOR2_X1 U770 ( .A(n711), .B(KEYINPUT52), .ZN(n712) );
  NOR2_X1 U771 ( .A1(n713), .A2(n712), .ZN(n719) );
  NAND2_X1 U772 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U773 ( .A(n716), .B(KEYINPUT122), .ZN(n717) );
  NAND2_X1 U774 ( .A1(n717), .A2(n761), .ZN(n718) );
  NOR2_X1 U775 ( .A1(n719), .A2(n718), .ZN(n725) );
  INV_X1 U776 ( .A(n760), .ZN(n723) );
  NOR2_X1 U777 ( .A1(n750), .A2(n721), .ZN(n722) );
  NAND2_X1 U778 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U779 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U780 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U781 ( .A(KEYINPUT123), .B(n728), .Z(n729) );
  XNOR2_X1 U782 ( .A(KEYINPUT53), .B(n729), .ZN(G75) );
  XOR2_X1 U783 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n732) );
  XNOR2_X1 U784 ( .A(n730), .B(KEYINPUT125), .ZN(n731) );
  XNOR2_X1 U785 ( .A(n732), .B(n731), .ZN(n734) );
  NAND2_X1 U786 ( .A1(n736), .A2(G469), .ZN(n733) );
  XOR2_X1 U787 ( .A(n734), .B(n733), .Z(n735) );
  NOR2_X1 U788 ( .A1(n743), .A2(n735), .ZN(G54) );
  NAND2_X1 U789 ( .A1(n736), .A2(G478), .ZN(n738) );
  XNOR2_X1 U790 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U791 ( .A1(n743), .A2(n739), .ZN(G63) );
  NAND2_X1 U792 ( .A1(n736), .A2(G217), .ZN(n741) );
  XNOR2_X1 U793 ( .A(n740), .B(n741), .ZN(n742) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(G66) );
  NOR2_X1 U795 ( .A1(n745), .A2(n744), .ZN(n747) );
  XNOR2_X1 U796 ( .A(KEYINPUT127), .B(KEYINPUT126), .ZN(n746) );
  XNOR2_X1 U797 ( .A(n747), .B(n746), .ZN(n754) );
  NAND2_X1 U798 ( .A1(G953), .A2(G224), .ZN(n748) );
  XNOR2_X1 U799 ( .A(KEYINPUT61), .B(n748), .ZN(n749) );
  NAND2_X1 U800 ( .A1(n749), .A2(G898), .ZN(n752) );
  OR2_X1 U801 ( .A1(n750), .A2(G953), .ZN(n751) );
  NAND2_X1 U802 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U803 ( .A(n754), .B(n753), .Z(G69) );
  XOR2_X1 U804 ( .A(n755), .B(n756), .Z(n759) );
  XNOR2_X1 U805 ( .A(n759), .B(G227), .ZN(n757) );
  NAND2_X1 U806 ( .A1(G900), .A2(n757), .ZN(n758) );
  NAND2_X1 U807 ( .A1(n758), .A2(G953), .ZN(n764) );
  XNOR2_X1 U808 ( .A(n760), .B(n759), .ZN(n762) );
  NAND2_X1 U809 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U810 ( .A1(n764), .A2(n763), .ZN(G72) );
  XNOR2_X1 U811 ( .A(G134), .B(n765), .ZN(n766) );
  XNOR2_X1 U812 ( .A(n766), .B(KEYINPUT116), .ZN(G36) );
  XOR2_X1 U813 ( .A(G125), .B(KEYINPUT37), .Z(n768) );
  XNOR2_X1 U814 ( .A(n767), .B(n768), .ZN(G27) );
  XOR2_X1 U815 ( .A(n769), .B(G122), .Z(G24) );
  XOR2_X1 U816 ( .A(n770), .B(G137), .Z(G39) );
  XOR2_X1 U817 ( .A(n771), .B(G119), .Z(G21) );
endmodule

