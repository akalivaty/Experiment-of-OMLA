//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1308, new_n1309;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n210));
  INV_X1    g0010(.A(G50), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G116), .ZN(new_n213));
  INV_X1    g0013(.A(G270), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(G58), .A2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(KEYINPUT65), .B1(G58), .B2(G68), .ZN(new_n227));
  AND3_X1   g0027(.A1(new_n226), .A2(G50), .A3(new_n227), .ZN(new_n228));
  AND2_X1   g0028(.A1(KEYINPUT64), .A2(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(KEYINPUT64), .A2(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n209), .A2(new_n223), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  AND2_X1   g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  OAI21_X1  g0054(.A(G274), .B1(new_n254), .B2(new_n232), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT68), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n256), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  OAI211_X1 g0060(.A(G1), .B(G13), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n258), .A2(new_n261), .A3(new_n262), .A4(G274), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n254), .A2(new_n232), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n258), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G226), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT69), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OR2_X1    g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1698), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G222), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n272), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G223), .A3(G1698), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n274), .B(new_n276), .C1(new_n217), .C2(new_n275), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n265), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n270), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT70), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n268), .A2(new_n269), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G169), .ZN(new_n285));
  OAI21_X1  g0085(.A(KEYINPUT70), .B1(new_n279), .B2(new_n282), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(G179), .B1(new_n284), .B2(new_n286), .ZN(new_n288));
  INV_X1    g0088(.A(G13), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(G1), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G20), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n232), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n204), .A2(G1), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  MUX2_X1   g0096(.A(new_n292), .B(new_n296), .S(G50), .Z(new_n297));
  INV_X1    g0097(.A(KEYINPUT72), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n294), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT71), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(G33), .A3(new_n231), .ZN(new_n303));
  INV_X1    g0103(.A(G58), .ZN(new_n304));
  INV_X1    g0104(.A(G68), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n211), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(G20), .A2(G33), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n306), .A2(G20), .B1(G150), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n300), .B1(new_n303), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n299), .A2(new_n309), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n287), .A2(new_n288), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT74), .B1(new_n299), .B2(new_n309), .ZN(new_n312));
  INV_X1    g0112(.A(new_n309), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n297), .B(KEYINPUT72), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT74), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n312), .A2(new_n316), .A3(KEYINPUT9), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT9), .B1(new_n312), .B2(new_n316), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n284), .A2(G200), .A3(new_n286), .ZN(new_n320));
  INV_X1    g0120(.A(G190), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n284), .B2(new_n286), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n319), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT10), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n322), .A2(new_n317), .A3(new_n318), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT10), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(new_n320), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n311), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n212), .A2(G1698), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(G223), .B2(G1698), .ZN(new_n331));
  AND2_X1   g0131(.A1(KEYINPUT76), .A2(G33), .ZN(new_n332));
  NOR2_X1   g0132(.A1(KEYINPUT76), .A2(G33), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT3), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n331), .B1(new_n271), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G87), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n259), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n265), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n257), .A2(new_n263), .B1(new_n266), .B2(G232), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT78), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT78), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n338), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G179), .ZN(new_n345));
  INV_X1    g0145(.A(new_n340), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n344), .A2(new_n285), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n302), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n291), .ZN(new_n349));
  INV_X1    g0149(.A(new_n296), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n302), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n304), .A2(new_n305), .ZN(new_n353));
  OAI21_X1  g0153(.A(G20), .B1(new_n353), .B2(new_n224), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n307), .A2(G159), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT3), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT64), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n204), .ZN(new_n359));
  NAND2_X1  g0159(.A1(KEYINPUT64), .A2(G20), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n359), .A2(KEYINPUT7), .A3(new_n360), .A4(new_n272), .ZN(new_n361));
  AND2_X1   g0161(.A1(KEYINPUT3), .A2(G33), .ZN(new_n362));
  NOR2_X1   g0162(.A1(KEYINPUT3), .A2(G33), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n362), .A2(new_n363), .A3(G20), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n357), .A2(new_n361), .B1(new_n364), .B2(KEYINPUT7), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n356), .B1(new_n365), .B2(G68), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n294), .B1(new_n366), .B2(KEYINPUT16), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT76), .B(G33), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n363), .B1(new_n369), .B2(KEYINPUT3), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n359), .A2(new_n360), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(KEYINPUT7), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n305), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n334), .A2(new_n204), .A3(new_n271), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT7), .ZN(new_n375));
  AOI211_X1 g0175(.A(new_n368), .B(new_n356), .C1(new_n373), .C2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n352), .B1(new_n367), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT77), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT77), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n379), .B(new_n352), .C1(new_n367), .C2(new_n376), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n347), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT18), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT18), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n347), .A2(new_n378), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  INV_X1    g0185(.A(new_n343), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n342), .B1(new_n338), .B2(new_n339), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n346), .A2(new_n321), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n377), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT17), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n377), .B1(new_n388), .B2(new_n389), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT17), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n382), .A2(new_n384), .A3(new_n394), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n266), .A2(G238), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n264), .A2(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n273), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n275), .A2(G232), .A3(G1698), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n265), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(new_n403), .A3(KEYINPUT13), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT13), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n264), .A2(new_n398), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n261), .B1(new_n400), .B2(new_n401), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT14), .B1(new_n409), .B2(new_n285), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n399), .A2(new_n403), .A3(KEYINPUT75), .A4(KEYINPUT13), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT75), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n406), .A2(new_n407), .B1(new_n412), .B2(new_n405), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G179), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT14), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n404), .A2(new_n408), .A3(new_n416), .A4(G169), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n410), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n307), .A2(G50), .B1(G20), .B2(new_n305), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n231), .A2(G33), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n419), .B1(new_n420), .B2(new_n217), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n421), .A2(KEYINPUT11), .A3(new_n294), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT11), .B1(new_n421), .B2(new_n294), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT12), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n292), .B2(new_n305), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n291), .A2(KEYINPUT12), .A3(G68), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n425), .A2(new_n426), .B1(new_n305), .B2(new_n350), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n422), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n418), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n428), .B1(new_n409), .B2(new_n385), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n321), .B1(new_n411), .B2(new_n413), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n292), .A2(new_n217), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n296), .A2(G77), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  XOR2_X1   g0238(.A(KEYINPUT8), .B(G58), .Z(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n307), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n371), .A2(G77), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT15), .B(G87), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n440), .B(new_n441), .C1(new_n420), .C2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n438), .B1(new_n443), .B2(new_n294), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n257), .A2(new_n263), .B1(new_n266), .B2(G244), .ZN(new_n445));
  INV_X1    g0245(.A(G1698), .ZN(new_n446));
  OAI211_X1 g0246(.A(G232), .B(new_n446), .C1(new_n362), .C2(new_n363), .ZN(new_n447));
  OAI211_X1 g0247(.A(G238), .B(G1698), .C1(new_n362), .C2(new_n363), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n447), .B(new_n448), .C1(new_n219), .C2(new_n275), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n265), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G179), .ZN(new_n452));
  AOI211_X1 g0252(.A(new_n444), .B(new_n452), .C1(new_n285), .C2(new_n451), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n385), .B1(new_n445), .B2(new_n450), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n420), .A2(new_n442), .ZN(new_n455));
  INV_X1    g0255(.A(new_n307), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n231), .A2(new_n217), .B1(new_n301), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n294), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(new_n436), .A3(new_n437), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n445), .A2(new_n450), .A3(G190), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT73), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n445), .A2(new_n450), .A3(KEYINPUT73), .A4(G190), .ZN(new_n463));
  AOI211_X1 g0263(.A(new_n454), .B(new_n459), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NOR4_X1   g0264(.A1(new_n397), .A2(new_n435), .A3(new_n453), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n329), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n300), .B(new_n291), .C1(G1), .C2(new_n259), .ZN(new_n467));
  OR2_X1    g0267(.A1(new_n467), .A2(new_n213), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n292), .A2(new_n213), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  INV_X1    g0270(.A(G97), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n231), .B(new_n470), .C1(G33), .C2(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n293), .A2(new_n232), .B1(G20), .B2(new_n213), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(KEYINPUT20), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT20), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n468), .B(new_n469), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n220), .A2(G1698), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(G257), .B2(G1698), .ZN(new_n479));
  INV_X1    g0279(.A(G303), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n370), .A2(new_n479), .B1(new_n480), .B2(new_n275), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n265), .ZN(new_n482));
  XNOR2_X1  g0282(.A(KEYINPUT5), .B(G41), .ZN(new_n483));
  INV_X1    g0283(.A(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(new_n255), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n265), .B1(new_n485), .B2(new_n483), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n487), .B1(G270), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n477), .A2(new_n490), .A3(KEYINPUT21), .A4(G169), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT82), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n472), .A2(new_n473), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT20), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n474), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n291), .A2(G116), .ZN(new_n497));
  INV_X1    g0297(.A(new_n467), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(G116), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n285), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT82), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT21), .A4(new_n490), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n492), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n500), .A2(new_n490), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT21), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n490), .A2(new_n345), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(new_n477), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n477), .B1(new_n490), .B2(G200), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n486), .A2(new_n261), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n509), .A2(new_n214), .B1(new_n255), .B2(new_n486), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n265), .B2(new_n481), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G190), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n503), .A2(new_n507), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n369), .A2(G294), .ZN(new_n515));
  INV_X1    g0315(.A(G257), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G1698), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(G250), .B2(G1698), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n515), .B1(new_n370), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(new_n265), .B1(new_n488), .B2(G264), .ZN(new_n520));
  INV_X1    g0320(.A(new_n487), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n385), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n321), .A3(new_n521), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(KEYINPUT84), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT22), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n359), .A2(G87), .A3(new_n360), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n362), .A2(new_n363), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n369), .A2(new_n204), .A3(G116), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT23), .B1(new_n204), .B2(G107), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT23), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n371), .A2(new_n532), .A3(new_n219), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n529), .A2(new_n530), .A3(new_n531), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(KEYINPUT22), .A2(G87), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n370), .A2(new_n371), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT83), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n533), .A2(new_n530), .A3(new_n531), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT83), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n334), .A2(new_n271), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n540), .A2(KEYINPUT22), .A3(G87), .A4(new_n231), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n538), .A2(new_n539), .A3(new_n541), .A4(new_n529), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n537), .A2(KEYINPUT24), .A3(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n543), .B(new_n294), .C1(KEYINPUT24), .C2(new_n537), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT25), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n291), .B2(G107), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n292), .A2(KEYINPUT25), .A3(new_n219), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n498), .A2(G107), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT84), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n522), .A2(new_n549), .A3(new_n385), .ZN(new_n550));
  AND4_X1   g0350(.A1(new_n525), .A2(new_n544), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n543), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n294), .B1(new_n537), .B2(KEYINPUT24), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n548), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n522), .A2(G179), .ZN(new_n555));
  AOI21_X1  g0355(.A(G169), .B1(new_n520), .B2(new_n521), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT6), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n559), .A2(new_n471), .A3(G107), .ZN(new_n560));
  XNOR2_X1  g0360(.A(G97), .B(G107), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n560), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n562), .A2(new_n231), .B1(new_n217), .B2(new_n456), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n365), .A2(G107), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n563), .B1(new_n564), .B2(KEYINPUT79), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT79), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n365), .A2(new_n566), .A3(G107), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n300), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n292), .A2(KEYINPUT80), .A3(new_n471), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT80), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n291), .B2(G97), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n571), .C1(new_n467), .C2(new_n471), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(KEYINPUT81), .B1(new_n509), .B2(new_n516), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT81), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n488), .A2(new_n575), .A3(G257), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n487), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n273), .A2(KEYINPUT4), .A3(G244), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n275), .A2(G250), .A3(G1698), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n470), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n446), .A2(G244), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT4), .B1(new_n540), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n265), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G190), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(G200), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n573), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n442), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n291), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n231), .A2(G33), .A3(G97), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT19), .ZN(new_n593));
  NAND3_X1  g0393(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n231), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n336), .A2(new_n471), .A3(new_n219), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n592), .A2(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n540), .A2(G68), .A3(new_n231), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n591), .B1(new_n599), .B2(new_n294), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n498), .A2(new_n590), .ZN(new_n601));
  INV_X1    g0401(.A(new_n255), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n485), .ZN(new_n603));
  INV_X1    g0403(.A(G250), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n485), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n261), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n369), .A2(G116), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n218), .A2(G1698), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(G238), .B2(G1698), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n608), .B1(new_n370), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n607), .B1(new_n265), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n600), .A2(new_n601), .B1(new_n345), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n265), .ZN(new_n614));
  INV_X1    g0414(.A(new_n607), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n285), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n614), .A2(new_n615), .A3(G190), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n385), .B1(new_n614), .B2(new_n615), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n467), .A2(new_n336), .ZN(new_n621));
  AOI211_X1 g0421(.A(new_n591), .B(new_n621), .C1(new_n599), .C2(new_n294), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n613), .A2(new_n617), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n585), .A2(new_n285), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n577), .A2(new_n584), .A3(new_n345), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n624), .B(new_n625), .C1(new_n568), .C2(new_n572), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n558), .A2(new_n589), .A3(new_n623), .A4(new_n626), .ZN(new_n627));
  NOR4_X1   g0427(.A1(new_n466), .A2(new_n514), .A3(new_n551), .A4(new_n627), .ZN(G372));
  NAND2_X1  g0428(.A1(new_n325), .A2(new_n328), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n347), .A2(new_n377), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT18), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n347), .A2(new_n383), .A3(new_n377), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n434), .A2(new_n453), .B1(new_n418), .B2(new_n429), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n394), .A2(new_n396), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n311), .B1(new_n629), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  INV_X1    g0438(.A(new_n626), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT85), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n617), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n613), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n620), .A2(new_n622), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(KEYINPUT86), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT86), .B1(new_n642), .B2(new_n643), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n638), .B(new_n639), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n639), .A2(new_n623), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(KEYINPUT26), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n645), .A2(new_n646), .ZN(new_n651));
  INV_X1    g0451(.A(new_n551), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n589), .A2(new_n626), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n558), .A2(new_n503), .A3(new_n507), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n642), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n637), .B1(new_n657), .B2(new_n466), .ZN(G369));
  NAND2_X1  g0458(.A1(new_n503), .A2(new_n507), .ZN(new_n659));
  INV_X1    g0459(.A(new_n514), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT27), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n290), .A2(new_n359), .A3(new_n661), .A4(new_n360), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT87), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n231), .A2(KEYINPUT87), .A3(new_n661), .A4(new_n290), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G213), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n231), .A2(new_n290), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n667), .B1(new_n668), .B2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT88), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n666), .A2(new_n669), .A3(new_n673), .A4(G343), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n477), .ZN(new_n676));
  MUX2_X1   g0476(.A(new_n659), .B(new_n660), .S(new_n676), .Z(new_n677));
  AND2_X1   g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n558), .A2(new_n675), .ZN(new_n679));
  INV_X1    g0479(.A(new_n554), .ZN(new_n680));
  INV_X1    g0480(.A(new_n675), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n652), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n679), .B1(new_n682), .B2(new_n558), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n675), .B1(new_n503), .B2(new_n507), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n558), .B2(new_n675), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT89), .ZN(G399));
  INV_X1    g0490(.A(new_n207), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n596), .A2(G116), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G1), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n228), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(new_n693), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(G330), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n511), .A2(G179), .A3(new_n612), .A4(new_n520), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n585), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n511), .A2(new_n612), .A3(G179), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(new_n522), .A3(new_n585), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT90), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n612), .A2(new_n520), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n586), .A2(new_n707), .A3(new_n506), .A4(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n705), .A2(KEYINPUT90), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n681), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n702), .A2(new_n704), .A3(new_n708), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n675), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n710), .A2(new_n712), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  NOR4_X1   g0515(.A1(new_n627), .A2(new_n514), .A3(new_n551), .A4(new_n675), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n699), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT26), .B1(new_n651), .B2(new_n626), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(KEYINPUT26), .B2(new_n648), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT29), .B(new_n681), .C1(new_n720), .C2(new_n656), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n681), .B1(new_n650), .B2(new_n656), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT91), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT29), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n722), .A2(new_n724), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT91), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n718), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n698), .B1(new_n729), .B2(G1), .ZN(G364));
  NOR2_X1   g0530(.A1(new_n371), .A2(new_n289), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n203), .B1(new_n731), .B2(G45), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n692), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n678), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(G330), .B2(new_n677), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n691), .A2(new_n528), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G355), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(G116), .B2(new_n207), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n249), .A2(new_n484), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n691), .A2(new_n540), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n484), .B2(new_n228), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n739), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  OR3_X1    g0544(.A1(KEYINPUT92), .A2(G13), .A3(G33), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT92), .B1(G13), .B2(G33), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n232), .B1(G20), .B2(new_n285), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n734), .B1(new_n744), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT93), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n231), .A2(new_n345), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G190), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n321), .A2(new_n385), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G311), .A2(new_n759), .B1(new_n762), .B2(G326), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n385), .A2(G190), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n371), .A2(new_n345), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n321), .A2(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n371), .B1(new_n768), .B2(G179), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n766), .A2(G283), .B1(G294), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n756), .A2(new_n764), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT33), .B(G317), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n371), .A2(new_n345), .A3(new_n757), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n772), .A2(new_n773), .B1(G329), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n760), .A2(G20), .A3(new_n345), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n528), .B1(new_n777), .B2(new_n480), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n756), .A2(new_n767), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n778), .B1(new_n780), .B2(G322), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n763), .A2(new_n770), .A3(new_n776), .A4(new_n781), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n211), .A2(new_n761), .B1(new_n758), .B2(new_n217), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G107), .B2(new_n766), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n769), .B(KEYINPUT96), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n779), .B(KEYINPUT94), .Z(new_n786));
  OAI221_X1 g0586(.A(new_n784), .B1(new_n471), .B2(new_n785), .C1(new_n304), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n772), .A2(G68), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT95), .B(G159), .ZN(new_n789));
  OR3_X1    g0589(.A1(new_n774), .A2(KEYINPUT32), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(KEYINPUT32), .B1(new_n774), .B2(new_n789), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n777), .A2(new_n336), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n528), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n788), .A2(new_n790), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n782), .B1(new_n787), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n755), .B1(new_n750), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n749), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n796), .B1(new_n754), .B2(new_n753), .C1(new_n677), .C2(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n736), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  INV_X1    g0600(.A(new_n734), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n747), .A2(new_n750), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT97), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n801), .B1(new_n804), .B2(new_n217), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n453), .A2(new_n681), .ZN(new_n806));
  AOI21_X1  g0606(.A(KEYINPUT100), .B1(new_n675), .B2(new_n459), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT100), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n808), .B(new_n444), .C1(new_n672), .C2(new_n674), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n464), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n806), .B1(new_n810), .B2(new_n453), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n775), .A2(G311), .ZN(new_n813));
  INV_X1    g0613(.A(G294), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n779), .B2(new_n814), .C1(new_n213), .C2(new_n758), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n762), .A2(G303), .B1(new_n772), .B2(G283), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n766), .A2(G87), .ZN(new_n817));
  INV_X1    g0617(.A(new_n777), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n275), .B1(new_n818), .B2(G107), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n785), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n815), .B(new_n820), .C1(G97), .C2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n789), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G137), .A2(new_n762), .B1(new_n759), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G150), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n825), .B2(new_n771), .ZN(new_n826));
  INV_X1    g0626(.A(new_n786), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(G143), .B2(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT34), .Z(new_n829));
  OAI22_X1  g0629(.A1(new_n765), .A2(new_n305), .B1(new_n211), .B2(new_n777), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n830), .A2(KEYINPUT98), .B1(G58), .B2(new_n769), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n830), .A2(KEYINPUT98), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n540), .B1(new_n774), .B2(new_n833), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n834), .A2(KEYINPUT99), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(KEYINPUT99), .ZN(new_n836));
  AND4_X1   g0636(.A1(new_n831), .A2(new_n832), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n822), .B1(new_n829), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n750), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n805), .B1(new_n812), .B2(new_n748), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n722), .A2(new_n811), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n681), .B(new_n812), .C1(new_n650), .C2(new_n656), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n718), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(KEYINPUT101), .A3(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n845), .B(new_n801), .C1(new_n844), .C2(new_n843), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT101), .B1(new_n843), .B2(new_n844), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n840), .B1(new_n846), .B2(new_n847), .ZN(G384));
  INV_X1    g0648(.A(new_n562), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n849), .A2(KEYINPUT35), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(KEYINPUT35), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n850), .A2(G116), .A3(new_n233), .A4(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(KEYINPUT102), .B(KEYINPUT36), .Z(new_n853));
  XNOR2_X1  g0653(.A(new_n852), .B(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n228), .B(G77), .C1(new_n304), .C2(new_n305), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n211), .A2(G68), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n203), .B(G13), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n430), .A2(new_n675), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT105), .ZN(new_n860));
  INV_X1    g0660(.A(new_n352), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n356), .B1(new_n373), .B2(new_n375), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n294), .B1(new_n862), .B2(KEYINPUT16), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n376), .B1(new_n863), .B2(KEYINPUT103), .ZN(new_n864));
  INV_X1    g0664(.A(new_n356), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT7), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n370), .B2(new_n204), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n231), .A2(new_n866), .ZN(new_n868));
  OAI21_X1  g0668(.A(G68), .B1(new_n540), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n865), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n300), .B1(new_n870), .B2(new_n368), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT103), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n861), .B1(new_n864), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT104), .B1(new_n874), .B2(new_n670), .ZN(new_n875));
  INV_X1    g0675(.A(new_n376), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n871), .B2(new_n872), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n863), .A2(KEYINPUT103), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n352), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT104), .ZN(new_n880));
  INV_X1    g0680(.A(new_n670), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n397), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT37), .B1(new_n390), .B2(new_n391), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n378), .A2(new_n380), .A3(new_n881), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n885), .A2(new_n381), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n395), .B1(new_n879), .B2(new_n347), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(new_n875), .A3(new_n882), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n887), .B1(new_n889), .B2(KEYINPUT37), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n884), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n885), .A2(new_n381), .A3(new_n886), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n397), .A2(new_n883), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT38), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n860), .B(KEYINPUT39), .C1(new_n892), .C2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n631), .A2(new_n394), .A3(new_n396), .A4(new_n632), .ZN(new_n899));
  INV_X1    g0699(.A(new_n886), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n886), .A2(new_n630), .A3(new_n392), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n894), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n893), .A2(new_n894), .B1(new_n397), .B2(new_n883), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n905), .B1(new_n906), .B2(KEYINPUT38), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n898), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n895), .A2(KEYINPUT38), .A3(new_n896), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n891), .B1(new_n884), .B2(new_n890), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n908), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n913), .A2(new_n860), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n910), .A2(new_n914), .A3(KEYINPUT106), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT106), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n913), .A2(new_n860), .B1(new_n908), .B2(new_n907), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n911), .A2(new_n912), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT39), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT105), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n916), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n859), .B1(new_n915), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n842), .A2(new_n806), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n429), .A2(new_n675), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n430), .A2(new_n434), .A3(new_n924), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n429), .B(new_n675), .C1(new_n418), .C2(new_n433), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n918), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n928), .A2(new_n929), .B1(new_n633), .B2(new_n881), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n922), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n466), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n728), .A2(new_n721), .A3(new_n933), .A4(new_n725), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n637), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n932), .B(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n811), .B1(new_n925), .B2(new_n926), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n714), .A2(new_n711), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n937), .B1(new_n716), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT107), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n892), .B2(new_n905), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT40), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n911), .A2(new_n912), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n941), .B1(new_n942), .B2(KEYINPUT40), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n944), .A2(KEYINPUT40), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n940), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n466), .B1(new_n717), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n699), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n951), .B2(new_n949), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n936), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n203), .B2(new_n731), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n936), .A2(new_n953), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n858), .B1(new_n955), .B2(new_n956), .ZN(G367));
  OAI22_X1  g0757(.A1(new_n645), .A2(new_n646), .B1(new_n622), .B2(new_n681), .ZN(new_n958));
  OR3_X1    g0758(.A1(new_n642), .A2(new_n622), .A3(new_n681), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT43), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n653), .B1(new_n573), .B2(new_n681), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n639), .A2(new_n675), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n683), .A2(new_n686), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(KEYINPUT42), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT108), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n964), .A2(new_n558), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n675), .B1(new_n970), .B2(new_n626), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n967), .B2(KEYINPUT42), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n963), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n973), .A2(KEYINPUT43), .A3(new_n960), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n973), .B1(KEYINPUT43), .B2(new_n960), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n966), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n684), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n977), .B(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n692), .B(KEYINPUT41), .Z(new_n981));
  NAND2_X1  g0781(.A1(new_n687), .A2(KEYINPUT110), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(new_n678), .Z(new_n983));
  NOR2_X1   g0783(.A1(new_n683), .A2(new_n686), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n729), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n688), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n988), .A2(KEYINPUT109), .A3(new_n966), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT44), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT109), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n688), .B2(new_n978), .ZN(new_n992));
  OR3_X1    g0792(.A1(new_n989), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n990), .B1(new_n989), .B2(new_n992), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n988), .A2(new_n966), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT45), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n993), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n685), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n993), .A2(new_n684), .A3(new_n997), .A4(new_n994), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n987), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n981), .B1(new_n1001), .B2(new_n729), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n980), .B1(new_n1002), .B2(new_n733), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n751), .B1(new_n207), .B2(new_n442), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n742), .A2(new_n243), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n734), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n275), .B1(new_n777), .B2(new_n304), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n779), .A2(new_n825), .B1(new_n217), .B2(new_n765), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(G143), .C2(new_n762), .ZN(new_n1009));
  INV_X1    g0809(.A(G137), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n758), .A2(new_n211), .B1(new_n1010), .B2(new_n774), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(new_n772), .B2(new_n823), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1009), .B(new_n1012), .C1(new_n305), .C2(new_n785), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT112), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n818), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT46), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n777), .B2(new_n213), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1015), .B(new_n1017), .C1(new_n814), .C2(new_n771), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n827), .A2(G303), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1020));
  XOR2_X1   g0820(.A(KEYINPUT111), .B(G311), .Z(new_n1021));
  AOI22_X1  g0821(.A1(G283), .A2(new_n759), .B1(new_n762), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n540), .B1(new_n775), .B2(G317), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n769), .A2(G107), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n766), .A2(G97), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1013), .B1(new_n1020), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT47), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1006), .B1(new_n1028), .B2(new_n750), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n960), .B2(new_n797), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1003), .A2(new_n1030), .ZN(G387));
  NAND2_X1  g0831(.A1(new_n985), .A2(new_n733), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n683), .A2(new_n797), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n694), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n737), .A2(new_n1034), .B1(new_n219), .B2(new_n691), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n240), .A2(new_n484), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n439), .A2(new_n211), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT50), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n694), .B(new_n484), .C1(new_n305), .C2(new_n217), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n741), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1035), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n801), .B1(new_n1041), .B2(new_n751), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n762), .A2(G322), .B1(new_n772), .B2(new_n1021), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n480), .B2(new_n758), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G317), .B2(new_n827), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT48), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(KEYINPUT48), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n769), .A2(G283), .B1(new_n818), .B2(G294), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT49), .Z(new_n1050));
  OR2_X1    g0850(.A1(new_n1050), .A2(KEYINPUT113), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n540), .B1(new_n775), .B2(G326), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n213), .B2(new_n765), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n1050), .B2(KEYINPUT113), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n821), .A2(new_n590), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n348), .A2(new_n771), .B1(new_n758), .B2(new_n305), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n762), .A2(G159), .B1(new_n780), .B2(G50), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n370), .B1(G77), .B2(new_n818), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n1025), .A3(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1056), .B(new_n1059), .C1(G150), .C2(new_n775), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1051), .A2(new_n1054), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1042), .B1(new_n1061), .B2(new_n839), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n692), .B(KEYINPUT114), .Z(new_n1063));
  NAND2_X1  g0863(.A1(new_n986), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n985), .A2(new_n729), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1032), .B1(new_n1033), .B2(new_n1062), .C1(new_n1064), .C2(new_n1065), .ZN(G393));
  INV_X1    g0866(.A(KEYINPUT115), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n999), .A2(new_n1067), .A3(new_n1000), .ZN(new_n1068));
  OR3_X1    g0868(.A1(new_n998), .A2(new_n1067), .A3(new_n685), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1001), .B(new_n1063), .C1(new_n1070), .C2(new_n987), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n751), .B1(new_n471), .B2(new_n207), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n742), .A2(new_n252), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n734), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n966), .A2(new_n797), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n759), .A2(new_n439), .B1(G143), .B2(new_n775), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n211), .B2(new_n771), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n817), .B(new_n540), .C1(new_n305), .C2(new_n777), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(G159), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n825), .A2(new_n761), .B1(new_n779), .B2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT51), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n821), .A2(G77), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1079), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(G283), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n528), .B1(new_n777), .B2(new_n1085), .C1(new_n765), .C2(new_n219), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G322), .B2(new_n775), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT117), .Z(new_n1088));
  AOI22_X1  g0888(.A1(new_n762), .A2(G317), .B1(new_n780), .B2(G311), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n1090));
  OR2_X1    g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n759), .A2(G294), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n772), .A2(G303), .B1(G116), .B2(new_n769), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1084), .B1(new_n1088), .B2(new_n1095), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1074), .B(new_n1075), .C1(new_n750), .C2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n1070), .B2(new_n733), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1071), .A2(new_n1098), .ZN(G390));
  OR2_X1    g0899(.A1(new_n810), .A2(new_n453), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n681), .B(new_n1100), .C1(new_n720), .C2(new_n656), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n718), .A2(new_n812), .A3(new_n927), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n1101), .A2(new_n806), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n699), .B1(new_n717), .B2(new_n950), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n927), .B1(new_n1104), .B2(new_n812), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n927), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n844), .B2(new_n811), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1104), .A2(new_n937), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1103), .A2(new_n1106), .B1(new_n1110), .B2(new_n923), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n933), .A2(new_n1104), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n934), .A2(new_n637), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT106), .B1(new_n910), .B2(new_n914), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n917), .A2(new_n920), .A3(new_n916), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n859), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n928), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1117), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n905), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n911), .A2(new_n1122), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1101), .A2(new_n806), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1119), .B(new_n1123), .C1(new_n1124), .C2(new_n1107), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1121), .A2(new_n1125), .A3(new_n1102), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1109), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1127));
  OAI211_X1 g0927(.A(KEYINPUT118), .B(new_n1116), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1109), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1121), .A2(new_n1125), .A3(new_n1102), .ZN(new_n1132));
  OAI21_X1  g0932(.A(KEYINPUT118), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1128), .A2(new_n1063), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1117), .A2(new_n747), .A3(new_n1118), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n734), .B1(new_n803), .B2(new_n302), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n771), .A2(new_n219), .B1(new_n814), .B2(new_n774), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n765), .A2(new_n305), .ZN(new_n1140));
  NOR4_X1   g0940(.A1(new_n1139), .A2(new_n275), .A3(new_n792), .A4(new_n1140), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n213), .A2(new_n779), .B1(new_n761), .B2(new_n1085), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G97), .B2(new_n759), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1141), .A2(new_n1143), .A3(new_n1083), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n775), .A2(G125), .ZN(new_n1145));
  INV_X1    g0945(.A(G128), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1146), .A2(new_n761), .B1(new_n771), .B2(new_n1010), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT54), .B(G143), .Z(new_n1148));
  AOI211_X1 g0948(.A(new_n1145), .B(new_n1147), .C1(new_n759), .C2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n818), .A2(G150), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT53), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G132), .B2(new_n780), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1149), .B(new_n1152), .C1(new_n1080), .C2(new_n785), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n275), .B1(new_n765), .B2(new_n211), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT119), .Z(new_n1155));
  OAI21_X1  g0955(.A(new_n1144), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1138), .B1(new_n1156), .B2(new_n750), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1136), .A2(new_n733), .B1(new_n1137), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1135), .A2(new_n1158), .ZN(G378));
  INV_X1    g0959(.A(KEYINPUT121), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n311), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n629), .A2(new_n1161), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n312), .A2(new_n316), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1163), .A2(new_n670), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1164), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n329), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1168), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n329), .A2(new_n1166), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n311), .B(new_n1164), .C1(new_n325), .C2(new_n328), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1169), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n948), .B2(new_n699), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1169), .A2(new_n1173), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n946), .A2(new_n947), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n945), .B1(new_n1123), .B2(new_n943), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1176), .B(G330), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n922), .A2(new_n931), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1119), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1175), .A2(new_n1179), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1181), .A2(new_n1182), .A3(new_n930), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1160), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n922), .A2(new_n931), .A3(new_n1175), .A4(new_n1179), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1182), .B1(new_n1181), .B2(new_n930), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1185), .A2(new_n1186), .A3(KEYINPUT121), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1174), .A2(new_n747), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n747), .A2(G50), .A3(new_n750), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n370), .A2(new_n260), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G77), .B2(new_n818), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n821), .A2(G68), .B1(new_n1192), .B2(KEYINPUT120), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(KEYINPUT120), .B2(new_n1192), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n772), .A2(G97), .B1(new_n766), .B2(G58), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n219), .B2(new_n779), .C1(new_n442), .C2(new_n758), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n761), .A2(new_n213), .B1(new_n1085), .B2(new_n774), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(new_n1194), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(G50), .B1(new_n259), .B2(new_n260), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1198), .A2(KEYINPUT58), .B1(new_n1191), .B2(new_n1199), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G125), .A2(new_n762), .B1(new_n759), .B2(G137), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n772), .A2(G132), .B1(new_n818), .B2(new_n1148), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n1146), .C2(new_n779), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G150), .B2(new_n821), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n259), .B(new_n260), .C1(new_n765), .C2(new_n789), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G124), .B2(new_n775), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT59), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1208), .B1(new_n1204), .B2(new_n1209), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1200), .B1(KEYINPUT58), .B2(new_n1198), .C1(new_n1206), .C2(new_n1210), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n801), .B(new_n1190), .C1(new_n1211), .C2(new_n750), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1188), .A2(new_n733), .B1(new_n1189), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1131), .A2(new_n1132), .A3(new_n1112), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1184), .A2(new_n1187), .B1(new_n1215), .B2(new_n1115), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1063), .B1(new_n1216), .B2(KEYINPUT57), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1215), .A2(new_n1115), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n932), .A2(KEYINPUT122), .A3(new_n1182), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT122), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1185), .A2(new_n1186), .A3(new_n1221), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1219), .A2(KEYINPUT57), .A3(new_n1220), .A4(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1214), .B1(new_n1218), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(G375));
  INV_X1    g1025(.A(new_n981), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1116), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1107), .A2(new_n747), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n734), .B1(new_n803), .B2(G68), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n827), .A2(G137), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n540), .B1(new_n777), .B2(new_n1080), .C1(new_n765), .C2(new_n304), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n758), .A2(new_n825), .B1(new_n1146), .B2(new_n774), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(new_n772), .C2(new_n1148), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n821), .A2(G50), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n762), .A2(G132), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT124), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1231), .A2(new_n1234), .A3(new_n1235), .A4(new_n1237), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n774), .A2(new_n480), .B1(new_n471), .B2(new_n777), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT123), .Z(new_n1240));
  OAI22_X1  g1040(.A1(new_n219), .A2(new_n758), .B1(new_n771), .B2(new_n213), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1085), .A2(new_n779), .B1(new_n761), .B2(new_n814), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n275), .B1(new_n766), .B2(G77), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1055), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1238), .B1(new_n1240), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1230), .B1(new_n1246), .B2(new_n750), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1112), .A2(new_n733), .B1(new_n1229), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1228), .A2(new_n1248), .ZN(G381));
  OR2_X1    g1049(.A1(G393), .A2(G396), .ZN(new_n1250));
  OR4_X1    g1050(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT125), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G378), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1135), .A2(new_n1158), .A3(KEYINPUT125), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OR4_X1    g1055(.A1(G387), .A2(new_n1251), .A3(G375), .A4(new_n1255), .ZN(G407));
  NOR2_X1   g1056(.A1(new_n667), .A2(G343), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1224), .A2(new_n1253), .A3(new_n1254), .A4(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(G407), .A2(new_n1258), .A3(G213), .ZN(G409));
  NAND3_X1  g1059(.A1(G387), .A2(new_n1071), .A3(new_n1098), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(G390), .A2(new_n1003), .A3(new_n1030), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(G393), .B(new_n799), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1260), .A2(new_n1263), .A3(new_n1261), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1265), .A2(KEYINPUT127), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT127), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1223), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G378), .B(new_n1213), .C1(new_n1217), .C2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1222), .A2(new_n733), .A3(new_n1220), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1189), .A2(new_n1212), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1188), .A2(new_n1226), .A3(new_n1219), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1257), .B1(new_n1271), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT60), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1227), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(new_n1116), .A3(new_n1063), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1227), .A2(new_n1279), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1248), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(G384), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT62), .B1(new_n1278), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1271), .A2(new_n1277), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1257), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT126), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT126), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n1289), .B(new_n1257), .C1(new_n1271), .C2(new_n1277), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1284), .A2(KEYINPUT62), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1285), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1257), .A2(G2897), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1284), .B(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1269), .B1(new_n1293), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1265), .A2(new_n1298), .A3(new_n1266), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT63), .B1(new_n1278), .B2(new_n1284), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1278), .A2(new_n1295), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1291), .A2(KEYINPUT63), .A3(new_n1284), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1300), .A2(new_n1306), .ZN(G405));
  OAI21_X1  g1107(.A(new_n1271), .B1(new_n1224), .B2(new_n1255), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1308), .B(new_n1284), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1269), .B(new_n1309), .ZN(G402));
endmodule


