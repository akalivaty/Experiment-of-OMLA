//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT65), .Z(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G50), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G116), .B2(G270), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT67), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT68), .Z(new_n218));
  NAND2_X1  g0018(.A1(G87), .A2(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n218), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n210), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT1), .Z(new_n224));
  OR3_X1    g0024(.A1(new_n210), .A2(KEYINPUT66), .A3(G13), .ZN(new_n225));
  OAI21_X1  g0025(.A(KEYINPUT66), .B1(new_n210), .B2(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n206), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n229), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n224), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT69), .ZN(G361));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT70), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n212), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n201), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT71), .B(G107), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n249), .B(new_n253), .ZN(G351));
  OAI21_X1  g0054(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G150), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n231), .A2(G33), .ZN(new_n258));
  XOR2_X1   g0058(.A(KEYINPUT8), .B(G58), .Z(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n255), .B(new_n257), .C1(new_n258), .C2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n230), .ZN(new_n263));
  INV_X1    g0063(.A(G13), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n264), .A2(new_n231), .A3(G1), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n261), .A2(new_n263), .B1(new_n212), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n263), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n266), .B1(new_n212), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G222), .ZN(new_n278));
  INV_X1    g0078(.A(G223), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n276), .B(new_n278), .C1(new_n279), .C2(new_n277), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G1), .A3(G13), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n280), .B(new_n283), .C1(G77), .C2(new_n276), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n285), .A2(KEYINPUT72), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(KEYINPUT72), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n286), .A2(G274), .A3(new_n287), .A4(new_n282), .ZN(new_n288));
  AND3_X1   g0088(.A1(new_n282), .A2(KEYINPUT73), .A3(new_n285), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT73), .B1(new_n282), .B2(new_n285), .ZN(new_n290));
  OAI21_X1  g0090(.A(G226), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n284), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G169), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n292), .A2(G179), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n271), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(G200), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n297), .B(new_n299), .C1(new_n271), .C2(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n271), .A2(new_n300), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT10), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n296), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(G238), .B1(new_n289), .B2(new_n290), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n213), .A2(new_n277), .ZN(new_n309));
  INV_X1    g0109(.A(G232), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G1698), .ZN(new_n311));
  AND2_X1   g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NOR2_X1   g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n309), .B(new_n311), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G33), .A2(G97), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n283), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n308), .A2(new_n317), .A3(new_n288), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT13), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT13), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n308), .A2(new_n317), .A3(new_n320), .A4(new_n288), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT77), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT14), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n322), .A2(G169), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n324), .ZN(new_n326));
  AOI211_X1 g0126(.A(new_n293), .B(new_n326), .C1(new_n319), .C2(new_n321), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n319), .A2(G179), .A3(new_n321), .ZN(new_n328));
  NAND2_X1  g0128(.A1(KEYINPUT77), .A2(KEYINPUT14), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n325), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n267), .A2(G68), .A3(new_n269), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT75), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n267), .A2(KEYINPUT75), .A3(G68), .A4(new_n269), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n264), .A2(G1), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(G20), .A3(new_n202), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT12), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT11), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n256), .A2(G50), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n202), .A2(G20), .ZN(new_n342));
  INV_X1    g0142(.A(G77), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n341), .B(new_n342), .C1(new_n343), .C2(new_n258), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n340), .B1(new_n344), .B2(new_n263), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n340), .A3(new_n263), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n336), .B(new_n339), .C1(new_n345), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT76), .ZN(new_n349));
  INV_X1    g0149(.A(new_n345), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n346), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT76), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n351), .A2(new_n352), .A3(new_n339), .A4(new_n336), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n331), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n270), .A2(new_n343), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n259), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT15), .B(G87), .Z(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n357), .B1(new_n258), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n356), .B1(new_n360), .B2(new_n263), .ZN(new_n361));
  INV_X1    g0161(.A(new_n265), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(G77), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n277), .A2(G232), .ZN(new_n366));
  INV_X1    g0166(.A(G238), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n276), .B(new_n366), .C1(new_n367), .C2(new_n277), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(new_n283), .C1(G107), .C2(new_n276), .ZN(new_n369));
  OAI21_X1  g0169(.A(G244), .B1(new_n289), .B2(new_n290), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(new_n288), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n293), .ZN(new_n372));
  INV_X1    g0172(.A(G179), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n369), .A2(new_n373), .A3(new_n288), .A4(new_n370), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n365), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n371), .A2(G200), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n369), .A2(G190), .A3(new_n288), .A4(new_n370), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n375), .B1(new_n365), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT74), .B1(new_n322), .B2(new_n298), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n322), .A2(G200), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT74), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n319), .A2(new_n383), .A3(G190), .A4(new_n321), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n381), .A2(new_n354), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n355), .A2(new_n380), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n260), .A2(new_n265), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n270), .B2(new_n260), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n274), .A2(new_n231), .A3(new_n275), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n231), .A4(new_n275), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT79), .B1(new_n395), .B2(G68), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT79), .ZN(new_n397));
  AOI211_X1 g0197(.A(new_n397), .B(new_n202), .C1(new_n393), .C2(new_n394), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n400), .A2(G20), .B1(G159), .B2(new_n256), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT16), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT78), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n393), .A2(new_n403), .A3(new_n394), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n391), .A2(KEYINPUT78), .A3(new_n392), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(G68), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(KEYINPUT16), .A3(new_n401), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n263), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n390), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G87), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT80), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n279), .A2(new_n277), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n213), .A2(G1698), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(new_n413), .C1(new_n312), .C2(new_n313), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n283), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n282), .A2(G232), .A3(new_n285), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(new_n288), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT81), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n417), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n415), .B2(new_n283), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(KEYINPUT81), .A3(new_n288), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G200), .ZN(new_n425));
  INV_X1    g0225(.A(new_n418), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n424), .A2(new_n425), .B1(new_n298), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n387), .B1(new_n409), .B2(new_n427), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n407), .A2(new_n263), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n395), .A2(G68), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n397), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n395), .A2(KEYINPUT79), .A3(G68), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n401), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT16), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n389), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n422), .A2(KEYINPUT81), .A3(new_n288), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT81), .B1(new_n422), .B2(new_n288), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n425), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n426), .A2(new_n298), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n436), .A2(KEYINPUT17), .A3(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n428), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n437), .A2(new_n438), .ZN(new_n445));
  OAI22_X1  g0245(.A1(new_n445), .A2(G169), .B1(G179), .B2(new_n418), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n444), .B1(new_n436), .B2(new_n446), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n424), .A2(new_n293), .B1(new_n373), .B2(new_n426), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n409), .A2(KEYINPUT18), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n307), .A2(new_n386), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n231), .A2(G33), .A3(G116), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n231), .A2(G107), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n454), .B(KEYINPUT23), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT22), .ZN(new_n456));
  AOI21_X1  g0256(.A(G20), .B1(new_n274), .B2(new_n275), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(G87), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n231), .B(G87), .C1(new_n312), .C2(new_n313), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(KEYINPUT22), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n453), .B(new_n455), .C1(new_n458), .C2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT24), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n457), .A2(new_n456), .A3(G87), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(KEYINPUT22), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n466), .A2(KEYINPUT24), .A3(new_n453), .A4(new_n455), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(new_n263), .A3(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n362), .B(new_n267), .C1(G1), .C2(new_n273), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G107), .ZN(new_n471));
  INV_X1    g0271(.A(G107), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n265), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g0273(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n474));
  XNOR2_X1  g0274(.A(new_n473), .B(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n276), .B1(G257), .B2(new_n277), .ZN(new_n476));
  NOR2_X1   g0276(.A1(G250), .A2(G1698), .ZN(new_n477));
  INV_X1    g0277(.A(G294), .ZN(new_n478));
  OAI22_X1  g0278(.A1(new_n476), .A2(new_n477), .B1(new_n273), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n283), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n268), .A2(G45), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n481), .A2(new_n483), .A3(G274), .A4(new_n282), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n283), .B1(new_n483), .B2(new_n481), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G264), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n480), .A2(G190), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n468), .A2(new_n471), .A3(new_n475), .A4(new_n487), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n479), .A2(new_n283), .B1(G264), .B2(new_n485), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n425), .B1(new_n489), .B2(new_n484), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n468), .A2(new_n471), .A3(new_n475), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT90), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n468), .A2(KEYINPUT90), .A3(new_n471), .A4(new_n475), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n489), .A2(new_n484), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G169), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n373), .B2(new_n497), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n491), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT88), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G264), .A2(G1698), .ZN(new_n502));
  OAI221_X1 g0302(.A(new_n502), .B1(new_n221), .B2(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n503), .B(new_n283), .C1(G303), .C2(new_n276), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n481), .A2(new_n483), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G270), .A3(new_n282), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n506), .A3(new_n484), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G169), .ZN(new_n508));
  INV_X1    g0308(.A(G116), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n469), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G283), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n220), .A2(KEYINPUT83), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT83), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G97), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n231), .B(new_n511), .C1(new_n515), .C2(G33), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n262), .A2(new_n230), .B1(G20), .B2(new_n509), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT20), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n516), .A2(KEYINPUT20), .A3(new_n517), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n510), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n265), .A2(new_n509), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n508), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n501), .B1(new_n524), .B2(KEYINPUT21), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n504), .A2(new_n506), .A3(G179), .A4(new_n484), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT21), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n508), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n470), .A2(G116), .ZN(new_n529));
  INV_X1    g0329(.A(new_n521), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT20), .B1(new_n516), .B2(new_n517), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n529), .B(new_n523), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n507), .A2(G169), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(KEYINPUT88), .A3(new_n527), .ZN(new_n536));
  OR2_X1    g0336(.A1(new_n507), .A2(new_n298), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n507), .A2(G200), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n537), .A2(new_n523), .A3(new_n522), .A4(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n525), .A2(new_n533), .A3(new_n536), .A4(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT19), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n515), .B2(new_n258), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n457), .A2(G68), .ZN(new_n543));
  XNOR2_X1  g0343(.A(KEYINPUT83), .B(G97), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n544), .A2(G87), .A3(G107), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n315), .A2(new_n541), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n546), .A2(G20), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n542), .B(new_n543), .C1(new_n545), .C2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(new_n263), .B1(new_n265), .B2(new_n359), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n470), .A2(new_n358), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n367), .A2(new_n277), .ZN(new_n552));
  INV_X1    g0352(.A(G244), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G1698), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n552), .B(new_n554), .C1(new_n312), .C2(new_n313), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G116), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n283), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n268), .A2(G45), .A3(G274), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n559), .B(KEYINPUT87), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n282), .A2(G250), .A3(new_n482), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n558), .A2(new_n561), .A3(new_n373), .A4(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n558), .A2(new_n561), .A3(new_n562), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n293), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n551), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(G200), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n282), .B1(new_n555), .B2(new_n556), .ZN(new_n568));
  INV_X1    g0368(.A(new_n562), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n568), .A2(new_n560), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G190), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n470), .A2(G87), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n549), .A2(new_n567), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n540), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT85), .ZN(new_n576));
  OAI21_X1  g0376(.A(G244), .B1(new_n312), .B2(new_n313), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT4), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(G1698), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n580), .B(G244), .C1(new_n313), .C2(new_n312), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n511), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(G250), .B1(new_n312), .B2(new_n313), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n277), .B1(new_n583), .B2(KEYINPUT4), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n576), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(KEYINPUT4), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G1698), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n577), .A2(new_n578), .B1(G33), .B2(G283), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(KEYINPUT85), .A4(new_n581), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n283), .ZN(new_n591));
  INV_X1    g0391(.A(new_n484), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT86), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n485), .B2(G257), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n485), .A2(new_n593), .A3(G257), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n591), .A2(G190), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n312), .A2(new_n313), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT7), .B1(new_n599), .B2(new_n231), .ZN(new_n600));
  INV_X1    g0400(.A(new_n394), .ZN(new_n601));
  OAI21_X1  g0401(.A(G107), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT6), .A4(new_n472), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT6), .ZN(new_n604));
  AND2_X1   g0404(.A1(G97), .A2(G107), .ZN(new_n605));
  NOR2_X1   g0405(.A1(G97), .A2(G107), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(G20), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n256), .A2(G77), .ZN(new_n610));
  XOR2_X1   g0410(.A(new_n610), .B(KEYINPUT82), .Z(new_n611));
  NAND3_X1  g0411(.A1(new_n602), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n263), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT84), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT84), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n615), .A3(new_n263), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n282), .B1(new_n585), .B2(new_n589), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n485), .A2(new_n593), .A3(G257), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n484), .B1(new_n619), .B2(new_n594), .ZN(new_n620));
  OAI21_X1  g0420(.A(G200), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n362), .A2(G97), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n470), .B2(G97), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n598), .A2(new_n617), .A3(new_n621), .A4(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n612), .A2(new_n615), .A3(new_n263), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n615), .B1(new_n612), .B2(new_n263), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n293), .B1(new_n618), .B2(new_n620), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n591), .A2(new_n373), .A3(new_n597), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n452), .A2(new_n500), .A3(new_n575), .A4(new_n631), .ZN(G372));
  AND3_X1   g0432(.A1(new_n409), .A2(KEYINPUT18), .A3(new_n448), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT18), .B1(new_n409), .B2(new_n448), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT93), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n375), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n365), .A2(KEYINPUT93), .A3(new_n372), .A4(new_n374), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n385), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n355), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n635), .B1(new_n641), .B2(new_n443), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n305), .A2(new_n306), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n296), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n452), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT92), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  NOR4_X1   g0448(.A1(new_n630), .A2(new_n574), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n569), .B1(new_n557), .B2(new_n283), .ZN(new_n650));
  AOI21_X1  g0450(.A(G169), .B1(new_n650), .B2(new_n561), .ZN(new_n651));
  NOR4_X1   g0451(.A1(new_n568), .A2(new_n560), .A3(new_n569), .A4(G179), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT91), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT91), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n565), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(new_n551), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n573), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n648), .B1(new_n630), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT92), .ZN(new_n659));
  INV_X1    g0459(.A(new_n630), .ZN(new_n660));
  INV_X1    g0460(.A(new_n574), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(KEYINPUT26), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n649), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n525), .A2(new_n533), .A3(new_n536), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n499), .A2(new_n492), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n488), .A2(new_n490), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n563), .B1(new_n570), .B2(G169), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n668), .A2(KEYINPUT91), .B1(new_n549), .B2(new_n550), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n549), .A2(new_n571), .A3(new_n572), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n669), .A2(new_n655), .B1(new_n670), .B2(new_n567), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n667), .A2(new_n630), .A3(new_n624), .A4(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n656), .B1(new_n666), .B2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n663), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n645), .B1(new_n646), .B2(new_n675), .ZN(G369));
  NAND2_X1  g0476(.A1(new_n337), .A2(new_n231), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n679), .A3(G213), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n500), .A2(new_n664), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n665), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(new_n682), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n496), .A2(new_n682), .ZN(new_n688));
  AND4_X1   g0488(.A1(G179), .A2(new_n480), .A3(new_n484), .A4(new_n486), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(G169), .B2(new_n497), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n494), .B2(new_n495), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n500), .A2(new_n688), .B1(new_n691), .B2(new_n682), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n664), .A2(new_n532), .A3(new_n682), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n683), .B1(new_n522), .B2(new_n523), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n540), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n687), .B1(new_n692), .B2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n227), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n545), .A2(new_n509), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n699), .A2(new_n268), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n234), .B2(new_n699), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT28), .Z(new_n703));
  NOR2_X1   g0503(.A1(new_n691), .A2(new_n664), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n672), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n627), .A2(new_n628), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(new_n661), .A3(new_n648), .A4(new_n629), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT26), .B1(new_n630), .B2(new_n657), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n656), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n683), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT94), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT94), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n712), .B(new_n683), .C1(new_n705), .C2(new_n709), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(KEYINPUT29), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n674), .A2(new_n715), .A3(new_n683), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G330), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n526), .A2(new_n564), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n591), .A2(new_n597), .A3(new_n489), .A4(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n618), .A2(new_n620), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(KEYINPUT30), .A3(new_n489), .A4(new_n719), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n507), .A2(new_n564), .A3(new_n373), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n725), .B(new_n497), .C1(new_n618), .C2(new_n620), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n722), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT31), .B1(new_n727), .B2(new_n682), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n575), .A2(new_n500), .A3(new_n631), .A4(new_n683), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n718), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n717), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n703), .B1(new_n733), .B2(G1), .ZN(G364));
  NAND3_X1  g0534(.A1(G355), .A2(new_n227), .A3(new_n276), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n249), .A2(G45), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n698), .A2(new_n276), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(G45), .B2(new_n233), .ZN(new_n738));
  OAI221_X1 g0538(.A(new_n735), .B1(G116), .B2(new_n227), .C1(new_n736), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n230), .B1(G20), .B2(new_n293), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n231), .A2(new_n373), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n298), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n298), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n373), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n748), .A2(G326), .B1(new_n751), .B2(G294), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n231), .A2(G179), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G190), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G329), .ZN(new_n757));
  INV_X1    g0557(.A(G283), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n753), .A2(new_n298), .A3(G200), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n752), .B(new_n757), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT95), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n746), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(KEYINPUT95), .B1(new_n231), .B2(new_n373), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n762), .A2(new_n763), .A3(new_n749), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n276), .B(new_n760), .C1(G322), .C2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n747), .A2(G190), .ZN(new_n767));
  INV_X1    g0567(.A(G317), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(KEYINPUT33), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n768), .A2(KEYINPUT33), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n767), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n753), .A2(G190), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G303), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n762), .A2(new_n763), .A3(new_n754), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G311), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n766), .A2(new_n771), .A3(new_n774), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G87), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n772), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n767), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n781), .A2(new_n202), .B1(new_n343), .B2(new_n775), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n780), .B(new_n782), .C1(G50), .C2(new_n748), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n276), .B1(new_n759), .B2(new_n472), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(G97), .B2(new_n751), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n783), .B(new_n785), .C1(new_n201), .C2(new_n764), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n756), .A2(G159), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT32), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n778), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT96), .Z(new_n790));
  AOI21_X1  g0590(.A(new_n745), .B1(new_n790), .B2(new_n743), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n264), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n268), .B1(new_n792), .B2(G45), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n699), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n742), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n791), .B(new_n795), .C1(new_n695), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n695), .A2(G330), .ZN(new_n798));
  INV_X1    g0598(.A(new_n795), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n696), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n797), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT97), .ZN(G396));
  NAND4_X1  g0602(.A1(new_n637), .A2(new_n365), .A3(new_n638), .A4(new_n682), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n365), .A2(new_n682), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n379), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT101), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n675), .B2(new_n682), .ZN(new_n809));
  INV_X1    g0609(.A(new_n806), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n683), .B(new_n810), .C1(new_n663), .C2(new_n673), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n729), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n731), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G330), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n812), .B(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n795), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n776), .A2(G116), .B1(G303), .B2(new_n748), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n758), .B2(new_n781), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT99), .Z(new_n821));
  AOI211_X1 g0621(.A(new_n276), .B(new_n821), .C1(G311), .C2(new_n756), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n773), .A2(G107), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n759), .A2(new_n779), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n765), .A2(G294), .B1(G97), .B2(new_n751), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT100), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n822), .A2(new_n823), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n756), .A2(G132), .ZN(new_n829));
  INV_X1    g0629(.A(new_n751), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n276), .B(new_n829), .C1(new_n830), .C2(new_n201), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n765), .A2(G143), .B1(G150), .B2(new_n767), .ZN(new_n832));
  INV_X1    g0632(.A(G137), .ZN(new_n833));
  INV_X1    g0633(.A(new_n748), .ZN(new_n834));
  INV_X1    g0634(.A(G159), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n832), .B1(new_n833), .B2(new_n834), .C1(new_n835), .C2(new_n775), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT34), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n759), .A2(new_n202), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n837), .B(new_n838), .C1(new_n212), .C2(new_n772), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n828), .B1(new_n831), .B2(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n840), .A2(new_n743), .B1(new_n740), .B2(new_n806), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n743), .A2(new_n740), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n795), .B1(G77), .B2(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT98), .Z(new_n845));
  AND2_X1   g0645(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n818), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G384));
  NOR2_X1   g0648(.A1(new_n375), .A2(new_n682), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n811), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT38), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n429), .A2(new_n435), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(new_n441), .A3(new_n390), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT16), .B1(new_n406), .B2(new_n401), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n390), .B1(new_n408), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n680), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n448), .A2(new_n856), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n854), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n409), .A2(new_n448), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n409), .A2(new_n857), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n854), .A2(new_n862), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n858), .B1(new_n443), .B2(new_n450), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n852), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n858), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n428), .A2(new_n442), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n869), .B1(new_n635), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n861), .A2(new_n865), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(KEYINPUT38), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n349), .A2(KEYINPUT102), .A3(new_n353), .A4(new_n682), .ZN(new_n875));
  NOR4_X1   g0675(.A1(new_n325), .A2(new_n875), .A3(new_n327), .A4(new_n330), .ZN(new_n876));
  OAI211_X1 g0676(.A(KEYINPUT102), .B(new_n385), .C1(new_n331), .C2(new_n354), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n349), .A2(new_n353), .A3(new_n682), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n851), .A2(new_n874), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n450), .A2(new_n857), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT103), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n854), .A2(new_n862), .A3(new_n863), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT37), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n886), .A2(new_n865), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n863), .B1(new_n443), .B2(new_n450), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n852), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT39), .B1(new_n889), .B2(new_n873), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n355), .A2(new_n682), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n868), .A2(KEYINPUT39), .A3(new_n873), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT103), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n880), .A2(new_n895), .A3(new_n882), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n884), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n646), .B1(new_n714), .B2(new_n716), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n898), .A2(new_n644), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n897), .B(new_n899), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n876), .B(new_n806), .C1(new_n877), .C2(new_n878), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n815), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n874), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n863), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n451), .A2(new_n906), .B1(new_n865), .B2(new_n886), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n873), .B1(new_n907), .B2(KEYINPUT38), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n902), .A2(new_n908), .A3(KEYINPUT40), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n452), .A2(new_n815), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(G330), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n900), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n268), .B2(new_n792), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n509), .B1(new_n608), .B2(KEYINPUT35), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n916), .B(new_n232), .C1(KEYINPUT35), .C2(new_n608), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT36), .ZN(new_n918));
  OAI21_X1  g0718(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n233), .A2(new_n919), .B1(G50), .B2(new_n202), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(G1), .A3(new_n264), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n915), .A2(new_n918), .A3(new_n921), .ZN(G367));
  INV_X1    g0722(.A(G143), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n276), .B1(new_n834), .B2(new_n923), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n767), .A2(G159), .B1(new_n751), .B2(G68), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n925), .B1(new_n343), .B2(new_n759), .C1(new_n833), .C2(new_n755), .ZN(new_n926));
  AOI211_X1 g0726(.A(new_n924), .B(new_n926), .C1(G150), .C2(new_n765), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n927), .B1(new_n212), .B2(new_n775), .C1(new_n201), .C2(new_n772), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n775), .A2(new_n758), .ZN(new_n929));
  OAI221_X1 g0729(.A(new_n599), .B1(new_n755), .B2(new_n768), .C1(new_n515), .C2(new_n759), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT108), .Z(new_n931));
  NAND2_X1  g0731(.A1(new_n773), .A2(G116), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT46), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n767), .A2(G294), .B1(new_n751), .B2(G107), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n765), .A2(G303), .B1(G311), .B2(new_n748), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n931), .A2(new_n933), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n928), .B1(new_n929), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT47), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n743), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n683), .B1(new_n549), .B2(new_n572), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n657), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n669), .A2(new_n655), .A3(new_n940), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n742), .ZN(new_n945));
  INV_X1    g0745(.A(new_n737), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n744), .B1(new_n227), .B2(new_n359), .C1(new_n245), .C2(new_n946), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n939), .A2(new_n945), .A3(new_n795), .A4(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT106), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n627), .A2(new_n682), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n631), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT104), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n660), .A2(new_n682), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n954), .A2(KEYINPUT42), .A3(new_n684), .ZN(new_n955));
  INV_X1    g0755(.A(new_n691), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n630), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n683), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT42), .B1(new_n954), .B2(new_n684), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n955), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT105), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT105), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n955), .A2(new_n962), .A3(new_n958), .A4(new_n959), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(new_n965), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n961), .A2(new_n968), .A3(new_n963), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n952), .A2(new_n953), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n696), .A2(new_n692), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n949), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n973), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n966), .A2(KEYINPUT106), .A3(new_n975), .A4(new_n969), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n970), .A2(new_n973), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n699), .B(KEYINPUT41), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n971), .A2(new_n687), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT44), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n954), .B2(new_n686), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n971), .A2(KEYINPUT44), .A3(new_n687), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n988), .A2(KEYINPUT107), .A3(new_n972), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n972), .A2(KEYINPUT107), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n983), .A2(new_n990), .A3(new_n987), .ZN(new_n991));
  INV_X1    g0791(.A(new_n733), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n664), .A2(new_n683), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n696), .A2(new_n692), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n994), .B2(new_n972), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n684), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n989), .A2(new_n991), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n980), .B1(new_n998), .B2(new_n733), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n978), .B1(new_n999), .B2(new_n794), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n948), .B1(new_n977), .B2(new_n1000), .ZN(G387));
  NAND3_X1  g0801(.A1(new_n700), .A2(new_n227), .A3(new_n276), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(G107), .B2(new_n227), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT109), .Z(new_n1004));
  INV_X1    g0804(.A(G45), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n737), .B1(new_n241), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(G68), .A2(G77), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n259), .A2(new_n212), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n545), .B(new_n509), .C1(new_n1008), .C2(KEYINPUT50), .ZN(new_n1009));
  AOI211_X1 g0809(.A(G45), .B(new_n1009), .C1(KEYINPUT50), .C2(new_n1008), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1006), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n744), .B1(new_n1004), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n795), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n743), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n756), .A2(G326), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n765), .A2(G317), .B1(G311), .B2(new_n767), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n748), .A2(G322), .ZN(new_n1017));
  INV_X1    g0817(.A(G303), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1016), .B(new_n1017), .C1(new_n1018), .C2(new_n775), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT48), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n758), .B2(new_n830), .C1(new_n478), .C2(new_n772), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n276), .B(new_n1015), .C1(new_n1022), .C2(KEYINPUT49), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(KEYINPUT49), .B2(new_n1022), .C1(new_n509), .C2(new_n759), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n767), .A2(new_n259), .B1(new_n751), .B2(new_n358), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n220), .B2(new_n759), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n748), .A2(G159), .B1(new_n773), .B2(G77), .ZN(new_n1027));
  INV_X1    g0827(.A(G150), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1027), .B1(new_n1028), .B2(new_n755), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n276), .B1(new_n764), .B2(new_n212), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n202), .B2(new_n775), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT110), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1014), .B1(new_n1024), .B2(new_n1033), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1013), .B(new_n1034), .C1(new_n692), .C2(new_n742), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n996), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1035), .B1(new_n1036), .B2(new_n794), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n699), .B1(new_n733), .B2(new_n1036), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1037), .B1(new_n1038), .B2(new_n997), .ZN(G393));
  INV_X1    g0839(.A(KEYINPUT111), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n972), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT111), .B1(new_n696), .B2(new_n692), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n988), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n983), .A2(new_n987), .A3(new_n1040), .A4(new_n972), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(new_n992), .C2(new_n996), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1045), .A2(new_n699), .A3(new_n998), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n793), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n253), .A2(new_n737), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n744), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n227), .A2(new_n515), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n795), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n765), .A2(G311), .B1(G317), .B2(new_n748), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n1055));
  AOI22_X1  g0855(.A1(new_n1054), .A2(new_n1055), .B1(G116), .B2(new_n751), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n599), .B1(new_n775), .B2(new_n478), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n472), .A2(new_n759), .B1(new_n772), .B2(new_n758), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1055), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1057), .B(new_n1058), .C1(new_n1053), .C2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n767), .A2(G303), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n756), .A2(G322), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1056), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n765), .A2(G159), .B1(G150), .B2(new_n748), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT51), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n830), .A2(new_n343), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n259), .B2(new_n776), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n212), .B2(new_n781), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT112), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1065), .B(new_n1069), .C1(G68), .C2(new_n773), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n276), .C1(new_n923), .C2(new_n755), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1063), .B1(new_n1071), .B2(new_n824), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1052), .B1(new_n1072), .B2(new_n743), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT114), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n971), .A2(new_n796), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OR3_X1    g0876(.A1(new_n1048), .A2(KEYINPUT115), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(KEYINPUT115), .B1(new_n1048), .B2(new_n1076), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1047), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(G390));
  NAND2_X1  g0880(.A1(new_n717), .A2(new_n452), .ZN(new_n1081));
  AND3_X1   g0881(.A1(new_n452), .A2(G330), .A3(new_n815), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n645), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n711), .A2(new_n713), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n849), .B1(new_n1085), .B2(new_n810), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n732), .A2(new_n807), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n879), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1087), .A2(new_n1088), .B1(new_n732), .B2(new_n901), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n732), .A2(new_n901), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n718), .B(new_n806), .C1(new_n730), .C2(new_n731), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1090), .B1(new_n1091), .B2(new_n879), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1086), .A2(new_n1089), .B1(new_n1092), .B2(new_n851), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1084), .A2(new_n1093), .A3(KEYINPUT116), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT116), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n898), .A2(new_n644), .A3(new_n1082), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n708), .A2(new_n656), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1097), .B(new_n707), .C1(new_n672), .C2(new_n704), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n712), .B1(new_n1098), .B2(new_n683), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n713), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n810), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1101), .A2(new_n1102), .A3(new_n850), .A4(new_n1090), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1092), .A2(new_n851), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1095), .B1(new_n1096), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1094), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n892), .B1(new_n889), .B2(new_n873), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n893), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1088), .B1(new_n811), .B2(new_n850), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n1110), .A2(new_n890), .B1(new_n1111), .B2(new_n892), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1090), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1088), .B1(new_n1101), .B2(new_n850), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1108), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1112), .B(new_n1090), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1107), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1114), .B(new_n1117), .C1(new_n1094), .C2(new_n1106), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1119), .A2(new_n699), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n741), .B1(new_n891), .B2(new_n893), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n838), .B1(new_n478), .B2(new_n755), .C1(new_n781), .C2(new_n472), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1066), .B(new_n1123), .C1(new_n544), .C2(new_n776), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n509), .B2(new_n764), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n599), .B1(new_n834), .B2(new_n758), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1125), .A2(new_n780), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n759), .A2(new_n212), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n756), .A2(G125), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n599), .B(new_n1129), .C1(G128), .C2(new_n748), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n772), .A2(new_n1028), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n765), .A2(G132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n767), .A2(G137), .B1(new_n751), .B2(G159), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT54), .B(G143), .Z(new_n1136));
  AOI211_X1 g0936(.A(new_n1128), .B(new_n1135), .C1(new_n776), .C2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n743), .B1(new_n1127), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1138), .B(new_n795), .C1(new_n259), .C2(new_n843), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1118), .A2(new_n793), .B1(new_n1122), .B2(new_n1139), .ZN(new_n1140));
  OR2_X1    g0940(.A1(new_n1121), .A2(new_n1140), .ZN(G378));
  OAI22_X1  g0941(.A1(new_n830), .A2(new_n202), .B1(new_n764), .B2(new_n472), .ZN(new_n1142));
  AOI211_X1 g0942(.A(G41), .B(new_n276), .C1(new_n756), .C2(G283), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n201), .B2(new_n759), .C1(new_n343), .C2(new_n772), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT118), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1142), .B(new_n1145), .C1(G116), .C2(new_n748), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n220), .B2(new_n781), .C1(new_n359), .C2(new_n775), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT58), .Z(new_n1148));
  INV_X1    g0948(.A(G124), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n273), .B1(new_n755), .B2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n765), .A2(G128), .B1(G125), .B2(new_n748), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n776), .A2(G137), .B1(G150), .B2(new_n751), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n767), .A2(G132), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n773), .A2(new_n1136), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  XOR2_X1   g0955(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1156));
  AOI211_X1 g0956(.A(G41), .B(new_n1150), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n835), .B2(new_n759), .C1(new_n1156), .C2(new_n1155), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n212), .B1(new_n312), .B2(G41), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT117), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n743), .B1(new_n1148), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n799), .B1(new_n212), .B2(new_n842), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1164));
  NOR2_X1   g0964(.A1(new_n307), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n307), .A2(new_n1164), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1166), .A2(new_n271), .A3(new_n857), .A4(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n271), .A2(new_n857), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1167), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1169), .B1(new_n1170), .B2(new_n1165), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1162), .B(new_n1163), .C1(new_n1173), .C2(new_n741), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT120), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n815), .A2(new_n901), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n868), .B2(new_n873), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n909), .B(G330), .C1(new_n1178), .C2(KEYINPUT40), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n1173), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n905), .A2(new_n1172), .A3(G330), .A4(new_n909), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1182), .A2(new_n897), .ZN(new_n1183));
  AOI211_X1 g0983(.A(KEYINPUT103), .B(new_n881), .C1(new_n1111), .C2(new_n874), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n895), .B1(new_n880), .B2(new_n882), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1186), .A2(new_n894), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1176), .B1(new_n1183), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1182), .A2(new_n897), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1186), .A2(new_n894), .A3(new_n1181), .A4(new_n1180), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n1190), .A3(KEYINPUT120), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1175), .B1(new_n1192), .B2(new_n794), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1120), .A2(new_n1096), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT57), .B1(new_n1120), .B2(new_n1096), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1197), .A2(KEYINPUT57), .B1(new_n1198), .B2(new_n1192), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n699), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1193), .B1(new_n1199), .B2(new_n1200), .ZN(G375));
  NAND2_X1  g1001(.A1(new_n1084), .A2(new_n1093), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1107), .A2(new_n979), .A3(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n772), .A2(new_n835), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n276), .B1(new_n759), .B2(new_n201), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT121), .Z(new_n1206));
  AOI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(G128), .C2(new_n756), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n212), .B2(new_n830), .C1(new_n1028), .C2(new_n775), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT122), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n765), .A2(G137), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n767), .A2(new_n1136), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n748), .A2(G132), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n599), .B1(new_n781), .B2(new_n509), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n748), .A2(G294), .B1(new_n751), .B2(new_n358), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n343), .B2(new_n759), .C1(new_n1018), .C2(new_n755), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1214), .B(new_n1216), .C1(G107), .C2(new_n776), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n220), .B2(new_n772), .C1(new_n758), .C2(new_n764), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1213), .A2(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n795), .B1(G68), .B2(new_n843), .C1(new_n1219), .C2(new_n1014), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n740), .B2(new_n1088), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n794), .B2(new_n1105), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1203), .A2(new_n1222), .ZN(G381));
  NOR2_X1   g1023(.A1(new_n1121), .A2(new_n1140), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1224), .B(new_n1193), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1225), .A2(G396), .A3(G393), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1079), .B(new_n948), .C1(new_n1000), .C2(new_n977), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1227), .A2(G384), .A3(G381), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(G407));
  OAI211_X1 g1029(.A(G407), .B(G213), .C1(G343), .C2(new_n1225), .ZN(G409));
  NAND2_X1  g1030(.A1(G387), .A2(G390), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1227), .ZN(new_n1232));
  XOR2_X1   g1032(.A(G393), .B(G396), .Z(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1231), .A2(new_n1227), .A3(new_n1233), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G213), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(G343), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G375), .B2(G378), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1192), .A2(new_n979), .A3(new_n1194), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT123), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1183), .A2(new_n1187), .A3(KEYINPUT124), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT124), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1175), .B1(new_n1247), .B2(new_n794), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT123), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1192), .A2(new_n1249), .A3(new_n979), .A4(new_n1194), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1243), .A2(new_n1224), .A3(new_n1248), .A4(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(KEYINPUT116), .B1(new_n1084), .B2(new_n1093), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1096), .A2(new_n1105), .A3(new_n1095), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(new_n1253), .A3(new_n1202), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(KEYINPUT60), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1202), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1255), .B(new_n699), .C1(KEYINPUT60), .C2(new_n1256), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1257), .A2(G384), .A3(new_n1222), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G384), .B1(new_n1257), .B2(new_n1222), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1241), .A2(new_n1251), .A3(new_n1260), .A4(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1198), .A2(new_n1192), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1117), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1266), .A2(new_n1113), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1084), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT57), .B1(new_n1268), .B2(new_n1195), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1200), .B1(new_n1264), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1193), .ZN(new_n1271));
  OAI21_X1  g1071(.A(G378), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1240), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1272), .A2(new_n1273), .A3(new_n1251), .A4(new_n1260), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1261), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1263), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1257), .A2(new_n1222), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n847), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1257), .A2(G384), .A3(new_n1222), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1240), .A2(G2897), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1272), .A2(new_n1273), .A3(new_n1251), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT61), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT125), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1238), .B1(new_n1277), .B2(new_n1288), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n1274), .A2(KEYINPUT63), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1274), .A2(KEYINPUT63), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1237), .A3(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT61), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT125), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1235), .A2(new_n1294), .A3(new_n1236), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1292), .A2(new_n1293), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1289), .A2(new_n1296), .ZN(G405));
  AND2_X1   g1097(.A1(new_n1272), .A2(new_n1225), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1260), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1302));
  OR3_X1    g1102(.A1(new_n1301), .A2(new_n1237), .A3(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1237), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(G402));
endmodule


