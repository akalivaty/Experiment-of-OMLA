//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1191, new_n1192, new_n1193, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(new_n201), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  INV_X1    g0015(.A(G1), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n212), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  AOI211_X1 g0022(.A(new_n215), .B(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n214), .B1(new_n223), .B2(KEYINPUT0), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT0), .B2(new_n223), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT64), .Z(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT66), .ZN(new_n229));
  AND2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n228), .A2(new_n229), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n227), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OR2_X1    g0032(.A1(new_n232), .A2(KEYINPUT67), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(KEYINPUT67), .ZN(new_n235));
  AOI22_X1  g0035(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  AOI22_X1  g0037(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n238));
  NAND3_X1  g0038(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g0039(.A(new_n218), .B1(new_n234), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g0040(.A(new_n226), .B1(KEYINPUT1), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g0041(.A(new_n241), .B1(KEYINPUT1), .B2(new_n240), .ZN(G361));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  INV_X1    g0043(.A(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT2), .B(G226), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G264), .B(G270), .Z(new_n248));
  XNOR2_X1  g0048(.A(G250), .B(G257), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G358));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n202), .A2(G68), .ZN(new_n255));
  INV_X1    g0055(.A(G68), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G50), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(G58), .B(G77), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n254), .B(new_n260), .ZN(G351));
  OAI21_X1  g0061(.A(new_n216), .B1(G41), .B2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n266), .A2(new_n262), .ZN(new_n267));
  XOR2_X1   g0067(.A(KEYINPUT68), .B(G226), .Z(new_n268));
  AND2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(G222), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(G223), .A3(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(G77), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n276), .B(new_n277), .C1(new_n278), .C2(new_n274), .ZN(new_n279));
  AOI211_X1 g0079(.A(new_n264), .B(new_n269), .C1(new_n265), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G190), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n212), .A2(new_n270), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AOI22_X1  g0083(.A1(G150), .A2(new_n283), .B1(new_n203), .B2(G20), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n212), .A2(G33), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n211), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n216), .A2(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G50), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT69), .ZN(new_n293));
  INV_X1    g0093(.A(new_n289), .ZN(new_n294));
  INV_X1    g0094(.A(G13), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n293), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n290), .B(new_n298), .C1(G50), .C2(new_n297), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n300), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n281), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G200), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n280), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n281), .A2(new_n301), .A3(KEYINPUT71), .A4(new_n302), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G20), .A2(G77), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n311), .B1(new_n285), .B2(new_n282), .C1(new_n286), .C2(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n313), .A2(new_n289), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n296), .A2(new_n278), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n289), .B1(new_n216), .B2(G20), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n315), .B1(new_n317), .B2(new_n278), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n264), .B1(new_n267), .B2(G244), .ZN(new_n321));
  NOR2_X1   g0121(.A1(G232), .A2(G1698), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n275), .A2(G238), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n274), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n324), .B(new_n265), .C1(G107), .C2(new_n274), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n320), .B1(G200), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(new_n326), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT70), .ZN(new_n330));
  INV_X1    g0130(.A(G169), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n330), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n326), .A2(G179), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n319), .B1(new_n333), .B2(KEYINPUT70), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n307), .B(new_n308), .C1(new_n303), .C2(new_n305), .ZN(new_n338));
  INV_X1    g0138(.A(G179), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n280), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n340), .B(new_n299), .C1(G169), .C2(new_n280), .ZN(new_n341));
  AND4_X1   g0141(.A1(new_n310), .A2(new_n337), .A3(new_n338), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n244), .A2(G1698), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n274), .B(new_n343), .C1(G226), .C2(G1698), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G97), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n266), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n266), .A2(new_n262), .ZN(new_n347));
  INV_X1    g0147(.A(G238), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n347), .A2(new_n348), .B1(new_n263), .B2(new_n262), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT13), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT13), .B1(new_n346), .B2(new_n349), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(G179), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT73), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT14), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n352), .A2(KEYINPUT72), .A3(new_n353), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT72), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n350), .A2(new_n359), .A3(new_n351), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(G169), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(KEYINPUT73), .A2(KEYINPUT14), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n362), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n358), .A2(G169), .A3(new_n364), .A4(new_n360), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n357), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n297), .A2(KEYINPUT12), .A3(G68), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT12), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n296), .B2(new_n256), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n367), .A2(new_n369), .B1(new_n317), .B2(new_n256), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n286), .A2(new_n278), .B1(new_n212), .B2(G68), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n282), .A2(new_n202), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n289), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT11), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n373), .A2(new_n374), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n370), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n366), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n358), .A2(G200), .A3(new_n360), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n352), .A2(G190), .A3(new_n353), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n342), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n285), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n296), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n317), .B2(new_n383), .ZN(new_n385));
  INV_X1    g0185(.A(G58), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(new_n256), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n387), .A2(new_n201), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(G20), .B1(G159), .B2(new_n283), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n272), .A2(KEYINPUT74), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT74), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT3), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n393), .A3(G33), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n271), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT75), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .A4(new_n212), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G68), .ZN(new_n399));
  AOI21_X1  g0199(.A(G20), .B1(new_n394), .B2(new_n271), .ZN(new_n400));
  NAND2_X1  g0200(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT76), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n403), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n394), .A2(new_n271), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n401), .B(new_n406), .C1(new_n407), .C2(G20), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT76), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(G68), .A4(new_n398), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n390), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n294), .B1(new_n411), .B2(KEYINPUT16), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n273), .B1(new_n414), .B2(G33), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n415), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n397), .B1(new_n274), .B2(G20), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n256), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n413), .B1(new_n418), .B2(new_n390), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n385), .B1(new_n412), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n264), .B1(new_n267), .B2(G232), .ZN(new_n421));
  MUX2_X1   g0221(.A(G223), .B(G226), .S(G1698), .Z(new_n422));
  AOI22_X1  g0222(.A1(new_n407), .A2(new_n422), .B1(G33), .B2(G87), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n421), .B1(new_n423), .B2(new_n266), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n328), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(G200), .B2(new_n424), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT17), .B1(new_n420), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n405), .A2(new_n410), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(KEYINPUT16), .A3(new_n389), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(new_n419), .A3(new_n289), .ZN(new_n430));
  INV_X1    g0230(.A(new_n385), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n431), .A3(new_n426), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT77), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT77), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n430), .A2(new_n434), .A3(new_n431), .A4(new_n426), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n427), .B1(new_n436), .B2(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n430), .A2(new_n431), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n424), .A2(G169), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n339), .B2(new_n424), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT18), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n441), .B(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n382), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n297), .B(new_n294), .C1(G1), .C2(new_n270), .ZN(new_n446));
  INV_X1    g0246(.A(G107), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n296), .A2(KEYINPUT25), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT25), .B1(new_n296), .B2(new_n447), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n446), .A2(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n407), .A2(KEYINPUT22), .A3(new_n212), .A4(G87), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT22), .ZN(new_n453));
  INV_X1    g0253(.A(new_n274), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n212), .A2(G87), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT23), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n212), .B2(G107), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n447), .A2(KEYINPUT23), .A3(G20), .ZN(new_n459));
  INV_X1    g0259(.A(G116), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n270), .A2(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n458), .A2(new_n459), .B1(new_n461), .B2(new_n212), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n452), .A2(new_n456), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n463), .B(KEYINPUT24), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n451), .B1(new_n464), .B2(new_n289), .ZN(new_n465));
  NOR2_X1   g0265(.A1(G250), .A2(G1698), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n221), .B2(G1698), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n407), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G294), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n266), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT85), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT85), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n407), .A2(new_n467), .B1(G33), .B2(G294), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n266), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT5), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT79), .B1(new_n475), .B2(G41), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT79), .ZN(new_n477));
  INV_X1    g0277(.A(G41), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT5), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n475), .A2(G41), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n476), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G45), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G1), .ZN(new_n483));
  AOI211_X1 g0283(.A(new_n222), .B(new_n265), .C1(new_n481), .C2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n481), .A2(G274), .A3(new_n266), .A4(new_n483), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n471), .A2(new_n474), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G169), .ZN(new_n489));
  OAI21_X1  g0289(.A(KEYINPUT86), .B1(new_n470), .B2(new_n484), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n265), .B1(new_n481), .B2(new_n483), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G264), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT86), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n492), .B(new_n493), .C1(new_n473), .C2(new_n266), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n486), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G179), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n465), .B1(new_n489), .B2(new_n496), .ZN(new_n497));
  OAI22_X1  g0297(.A1(new_n495), .A2(G200), .B1(G190), .B2(new_n488), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n465), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT87), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n498), .A2(new_n465), .A3(KEYINPUT87), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g0303(.A(KEYINPUT78), .B(G97), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(KEYINPUT6), .A3(new_n447), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT6), .ZN(new_n506));
  INV_X1    g0306(.A(G97), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(new_n447), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n508), .B2(new_n205), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G20), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n278), .B2(new_n282), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n447), .B1(new_n416), .B2(new_n417), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n289), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n297), .A2(G97), .ZN(new_n515));
  INV_X1    g0315(.A(new_n446), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(G97), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n486), .B1(new_n491), .B2(G257), .ZN(new_n519));
  INV_X1    g0319(.A(G244), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(G1698), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT4), .B1(new_n407), .B2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n275), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G283), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n274), .A2(G250), .A3(G1698), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n265), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n518), .B1(new_n528), .B2(G200), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n528), .A2(KEYINPUT80), .A3(new_n328), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT80), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n519), .A2(new_n527), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n532), .B2(G190), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n529), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n528), .A2(G169), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n519), .A2(new_n527), .A3(G179), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT81), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n514), .A2(new_n538), .A3(new_n517), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n538), .B1(new_n514), .B2(new_n517), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n407), .A2(new_n212), .A3(G68), .ZN(new_n543));
  INV_X1    g0343(.A(new_n504), .ZN(new_n544));
  INV_X1    g0344(.A(G87), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n545), .A3(new_n447), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT19), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n212), .B1(new_n345), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n547), .B1(new_n544), .B2(new_n270), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n543), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n551), .A2(new_n289), .B1(new_n296), .B2(new_n312), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n265), .A2(new_n215), .A3(new_n483), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(G274), .B2(new_n483), .ZN(new_n554));
  NOR2_X1   g0354(.A1(G238), .A2(G1698), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n520), .B2(G1698), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n461), .B1(new_n407), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n554), .B1(new_n557), .B2(new_n266), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G200), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n516), .A2(G87), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n552), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n554), .B(G190), .C1(new_n557), .C2(new_n266), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n562), .B(KEYINPUT82), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n558), .A2(new_n331), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n554), .B(new_n339), .C1(new_n557), .C2(new_n266), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OR2_X1    g0366(.A1(new_n446), .A2(new_n312), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n552), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n561), .A2(new_n563), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n534), .A2(new_n542), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT21), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n296), .A2(new_n460), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n516), .A2(G116), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n460), .A2(G20), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n289), .A2(KEYINPUT84), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT84), .B1(new_n289), .B2(new_n574), .ZN(new_n576));
  OR2_X1    g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n212), .B(new_n524), .C1(new_n544), .C2(G33), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(KEYINPUT20), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT20), .B1(new_n577), .B2(new_n578), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n572), .B(new_n573), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G169), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n491), .A2(G270), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT83), .B1(new_n584), .B2(new_n485), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(KEYINPUT83), .A3(new_n485), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n222), .A2(G1698), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(G257), .B2(G1698), .ZN(new_n589));
  INV_X1    g0389(.A(G303), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n395), .A2(new_n589), .B1(new_n590), .B2(new_n274), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n586), .A2(new_n587), .B1(new_n265), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n571), .B1(new_n583), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n582), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(new_n265), .ZN(new_n595));
  INV_X1    g0395(.A(new_n587), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n595), .B(G190), .C1(new_n596), .C2(new_n585), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n594), .B(new_n597), .C1(new_n592), .C2(new_n304), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n595), .B1(new_n596), .B2(new_n585), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n599), .A2(new_n582), .A3(KEYINPUT21), .A4(G169), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n592), .A2(G179), .A3(new_n582), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n593), .A2(new_n598), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n570), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n445), .A2(new_n503), .A3(new_n603), .ZN(G372));
  AND2_X1   g0404(.A1(new_n310), .A2(new_n338), .ZN(new_n605));
  INV_X1    g0405(.A(new_n427), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n434), .B1(new_n420), .B2(new_n426), .ZN(new_n607));
  INV_X1    g0407(.A(new_n435), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT17), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n336), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n381), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n611), .B1(new_n378), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n441), .B(KEYINPUT18), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n605), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n341), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT88), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n498), .A2(new_n465), .A3(KEYINPUT87), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT87), .B1(new_n498), .B2(new_n465), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n566), .A2(new_n568), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n552), .A2(new_n559), .A3(new_n560), .A4(new_n562), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n534), .A2(new_n625), .A3(new_n542), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n619), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n501), .A2(new_n502), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n534), .A2(new_n625), .A3(new_n542), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(KEYINPUT88), .ZN(new_n630));
  INV_X1    g0430(.A(new_n497), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n601), .A2(new_n600), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n593), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n627), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n623), .A2(new_n537), .A3(new_n518), .A4(new_n624), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(KEYINPUT89), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n541), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n638), .A2(new_n539), .B1(new_n535), .B2(new_n536), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(new_n569), .A3(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT89), .B1(new_n635), .B2(new_n636), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n623), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n634), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n445), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n618), .A2(new_n647), .ZN(G369));
  NAND2_X1  g0448(.A1(new_n632), .A2(new_n593), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n295), .A2(G20), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n216), .ZN(new_n651));
  XOR2_X1   g0451(.A(new_n651), .B(KEYINPUT90), .Z(new_n652));
  INV_X1    g0452(.A(KEYINPUT27), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n654), .A2(new_n655), .A3(G213), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT91), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(G343), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(G343), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(new_n594), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n649), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n602), .B2(new_n662), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G330), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n503), .B1(new_n465), .B2(new_n661), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n631), .B2(new_n661), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n649), .A2(new_n661), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n672), .A2(new_n503), .B1(new_n497), .B2(new_n661), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(G399));
  NOR2_X1   g0474(.A1(new_n220), .A2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n546), .A2(G116), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G1), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n209), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT31), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n603), .A2(new_n503), .A3(new_n661), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n592), .A2(G179), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n528), .A2(new_n558), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n490), .A2(new_n494), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT92), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT30), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  OAI211_X1 g0489(.A(KEYINPUT92), .B(new_n689), .C1(new_n683), .C2(new_n686), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n528), .A2(new_n339), .A3(new_n558), .ZN(new_n691));
  OR3_X1    g0491(.A1(new_n592), .A2(new_n691), .A3(new_n495), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n688), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n661), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n681), .B1(new_n682), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT31), .B1(new_n693), .B2(new_n694), .ZN(new_n697));
  OAI21_X1  g0497(.A(G330), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n646), .A2(new_n661), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n633), .A2(new_n628), .A3(new_n629), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n644), .B1(new_n635), .B2(KEYINPUT26), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n639), .A2(new_n569), .A3(new_n636), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT93), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n704), .A2(new_n705), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT93), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n703), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .A3(new_n661), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n699), .B1(new_n702), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n680), .B1(new_n712), .B2(G1), .ZN(G364));
  AOI21_X1  g0513(.A(new_n216), .B1(new_n650), .B2(G45), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n675), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(G13), .A2(G33), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G20), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n665), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n211), .B1(G20), .B2(new_n331), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n220), .A2(new_n407), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n482), .B2(new_n210), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n482), .B2(new_n260), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n219), .A2(new_n274), .ZN(new_n729));
  INV_X1    g0529(.A(G355), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n729), .A2(new_n730), .B1(G116), .B2(new_n219), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT94), .Z(new_n732));
  AOI21_X1  g0532(.A(new_n724), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n212), .A2(new_n328), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(G179), .A3(new_n304), .ZN(new_n735));
  INV_X1    g0535(.A(G322), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n212), .A2(G190), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(G179), .A3(new_n304), .ZN(new_n738));
  INV_X1    g0538(.A(G311), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n735), .A2(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n339), .A2(new_n304), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n737), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  XNOR2_X1  g0543(.A(KEYINPUT33), .B(G317), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n274), .B(new_n740), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n304), .A2(G179), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n734), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G179), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n737), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G303), .A2(new_n748), .B1(new_n751), .B2(G329), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n734), .A2(new_n741), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n737), .A2(new_n746), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G326), .A2(new_n754), .B1(new_n756), .B2(G283), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n212), .B1(new_n749), .B2(G190), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G294), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n745), .A2(new_n752), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n735), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n762), .A2(G58), .B1(new_n754), .B2(G50), .ZN(new_n763));
  INV_X1    g0563(.A(new_n738), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(KEYINPUT95), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n764), .A2(KEYINPUT95), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n763), .B1(new_n256), .B2(new_n742), .C1(new_n768), .C2(new_n278), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  OR3_X1    g0570(.A1(new_n750), .A2(KEYINPUT32), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(KEYINPUT32), .B1(new_n750), .B2(new_n770), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n771), .B(new_n772), .C1(new_n507), .C2(new_n758), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n274), .B1(new_n747), .B2(new_n545), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n775), .A2(KEYINPUT96), .B1(new_n447), .B2(new_n755), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(KEYINPUT96), .B2(new_n775), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT97), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n761), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n733), .B1(new_n779), .B2(new_n722), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n717), .B1(new_n721), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n664), .B(G330), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(new_n782), .B2(new_n717), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT98), .ZN(G396));
  NAND2_X1  g0584(.A1(new_n694), .A2(new_n320), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n612), .B1(new_n329), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n336), .A2(new_n694), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n700), .B(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n716), .B1(new_n790), .B2(new_n698), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n698), .B2(new_n790), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n722), .A2(new_n718), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n717), .B1(new_n278), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n722), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n762), .A2(G143), .B1(new_n754), .B2(G137), .ZN(new_n796));
  INV_X1    g0596(.A(G150), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n796), .B1(new_n797), .B2(new_n742), .C1(new_n768), .C2(new_n770), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(KEYINPUT34), .ZN(new_n800));
  INV_X1    g0600(.A(G132), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n747), .A2(new_n202), .B1(new_n750), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n407), .B1(new_n386), .B2(new_n758), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(G68), .C2(new_n756), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT34), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n798), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n800), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G283), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n768), .A2(new_n460), .B1(new_n808), .B2(new_n742), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(KEYINPUT99), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(KEYINPUT99), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n755), .A2(new_n545), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G311), .B2(new_n751), .ZN(new_n813));
  INV_X1    g0613(.A(G294), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n814), .B2(new_n735), .C1(new_n590), .C2(new_n753), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n454), .B1(new_n758), .B2(new_n507), .C1(new_n447), .C2(new_n747), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n811), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n807), .B1(new_n810), .B2(new_n817), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n794), .B1(new_n795), .B2(new_n818), .C1(new_n788), .C2(new_n719), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n792), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G384));
  OR2_X1    g0621(.A1(new_n661), .A2(new_n377), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n381), .B(new_n822), .C1(new_n366), .C2(new_n377), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n366), .A2(new_n822), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(KEYINPUT100), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT100), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n823), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n829), .B(new_n788), .C1(new_n696), .C2(new_n697), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n429), .A2(new_n289), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n411), .A2(KEYINPUT16), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n431), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT101), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(KEYINPUT101), .B(new_n431), .C1(new_n832), .C2(new_n833), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n836), .A2(new_n656), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n836), .A2(new_n440), .A3(new_n837), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n609), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(KEYINPUT37), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT37), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT102), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n656), .B(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n438), .B1(new_n844), .B2(new_n440), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n609), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n838), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n444), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n847), .A2(KEYINPUT38), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT103), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT38), .ZN(new_n852));
  AND4_X1   g0652(.A1(new_n842), .A2(new_n845), .A3(new_n433), .A4(new_n435), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n840), .B2(KEYINPUT37), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n838), .B1(new_n437), .B2(new_n443), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n850), .A2(new_n851), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n851), .B1(new_n850), .B2(new_n856), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n831), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT40), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n438), .A2(new_n844), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n615), .B1(new_n437), .B2(KEYINPUT105), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT105), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n611), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n861), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT104), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n846), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n853), .A2(KEYINPUT104), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n845), .A2(new_n432), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT37), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n852), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n850), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n830), .A2(new_n860), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n859), .A2(new_n860), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n445), .B1(new_n696), .B2(new_n697), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT107), .ZN(new_n878));
  OAI21_X1  g0678(.A(G330), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n878), .B2(new_n876), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT39), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n378), .A2(new_n694), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n850), .A2(KEYINPUT39), .A3(new_n856), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n829), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n694), .B1(new_n634), .B2(new_n645), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n788), .ZN(new_n888));
  INV_X1    g0688(.A(new_n787), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n857), .B2(new_n858), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n443), .A2(new_n844), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n885), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n702), .A2(KEYINPUT106), .A3(new_n445), .A4(new_n711), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n445), .B(new_n711), .C1(new_n887), .C2(KEYINPUT29), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT106), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n617), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n893), .B(new_n898), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n880), .A2(new_n899), .B1(new_n216), .B2(new_n650), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n899), .B2(new_n880), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n510), .A2(KEYINPUT35), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n510), .A2(KEYINPUT35), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n902), .A2(G116), .A3(new_n213), .A4(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT36), .Z(new_n905));
  OR3_X1    g0705(.A1(new_n209), .A2(new_n278), .A3(new_n387), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n216), .B(G13), .C1(new_n906), .C2(new_n255), .ZN(new_n907));
  OR3_X1    g0707(.A1(new_n901), .A2(new_n905), .A3(new_n907), .ZN(G367));
  NAND2_X1  g0708(.A1(new_n552), .A2(new_n560), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n694), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n625), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n623), .B2(new_n910), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT43), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT108), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n694), .A2(new_n518), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n534), .A2(new_n542), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n694), .A2(new_n537), .A3(new_n518), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n672), .A2(new_n503), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT42), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n631), .B1(new_n916), .B2(new_n917), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n661), .B1(new_n921), .B2(new_n639), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n919), .A2(KEYINPUT42), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n914), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n912), .A2(KEYINPUT43), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n925), .B(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n670), .B1(new_n916), .B2(new_n917), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n927), .B(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n675), .B(KEYINPUT41), .Z(new_n930));
  NAND2_X1  g0730(.A1(new_n673), .A2(new_n918), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT45), .Z(new_n932));
  NOR2_X1   g0732(.A1(new_n673), .A2(new_n918), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT44), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n670), .A2(KEYINPUT109), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n935), .B(new_n936), .Z(new_n937));
  NAND2_X1  g0737(.A1(new_n672), .A2(new_n503), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n669), .B2(new_n672), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(new_n667), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n712), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n930), .B1(new_n943), .B2(new_n712), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n929), .B1(new_n944), .B2(new_n715), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n723), .B1(new_n219), .B2(new_n312), .C1(new_n726), .C2(new_n250), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n946), .A2(new_n716), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n747), .A2(new_n460), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT46), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(G107), .B2(new_n759), .ZN(new_n950));
  INV_X1    g0750(.A(new_n768), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(G283), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n735), .A2(new_n590), .B1(new_n753), .B2(new_n739), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n504), .B2(new_n756), .ZN(new_n954));
  INV_X1    g0754(.A(G317), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n742), .A2(new_n814), .B1(new_n750), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n407), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n950), .A2(new_n952), .A3(new_n954), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n951), .A2(G50), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n759), .A2(G68), .ZN(new_n960));
  INV_X1    g0760(.A(G143), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n753), .A2(new_n961), .B1(new_n747), .B2(new_n386), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n454), .B(new_n962), .C1(G150), .C2(new_n762), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n755), .A2(new_n278), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n742), .A2(new_n770), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(G137), .C2(new_n751), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n959), .A2(new_n960), .A3(new_n963), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n958), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT47), .Z(new_n969));
  INV_X1    g0769(.A(new_n720), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n947), .B1(new_n969), .B2(new_n795), .C1(new_n912), .C2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n945), .A2(new_n971), .ZN(G387));
  OR2_X1    g0772(.A1(new_n669), .A2(new_n970), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n677), .A2(new_n729), .B1(G107), .B2(new_n219), .ZN(new_n974));
  INV_X1    g0774(.A(new_n247), .ZN(new_n975));
  AOI21_X1  g0775(.A(G45), .B1(G68), .B2(G77), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT50), .B1(new_n383), .B2(new_n202), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n383), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n677), .B(new_n976), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n725), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n975), .A2(G45), .B1(KEYINPUT110), .B2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n980), .A2(KEYINPUT110), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n974), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n716), .B1(new_n983), .B2(new_n724), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n753), .A2(new_n736), .B1(new_n742), .B2(new_n739), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT112), .Z(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n590), .B2(new_n768), .C1(new_n955), .C2(new_n735), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT48), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n747), .A2(new_n814), .B1(new_n758), .B2(new_n808), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT49), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G116), .A2(new_n756), .B1(new_n751), .B2(G326), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n993), .A2(new_n395), .A3(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n992), .A2(KEYINPUT49), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n758), .A2(new_n312), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G50), .B2(new_n762), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT111), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G159), .A2(new_n754), .B1(new_n743), .B2(new_n383), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G68), .A2(new_n764), .B1(new_n756), .B2(G97), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G77), .A2(new_n748), .B1(new_n751), .B2(G150), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .A4(new_n407), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n995), .A2(new_n996), .B1(new_n999), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n984), .B1(new_n1004), .B2(new_n722), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n940), .A2(new_n715), .B1(new_n973), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n941), .A2(new_n675), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n712), .A2(new_n940), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(G393));
  OAI221_X1 g0809(.A(new_n723), .B1(new_n219), .B2(new_n544), .C1(new_n726), .C2(new_n254), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n716), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n747), .A2(new_n256), .B1(new_n750), .B2(new_n961), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n812), .B(new_n1012), .C1(G50), .C2(new_n743), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n395), .B1(G77), .B2(new_n759), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(new_n285), .C2(new_n768), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n735), .A2(new_n770), .B1(new_n753), .B2(new_n797), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT51), .Z(new_n1017));
  OAI22_X1  g0817(.A1(new_n735), .A2(new_n739), .B1(new_n753), .B2(new_n955), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT52), .Z(new_n1019));
  OAI221_X1 g0819(.A(new_n454), .B1(new_n758), .B2(new_n460), .C1(new_n447), .C2(new_n755), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n738), .A2(new_n814), .B1(new_n742), .B2(new_n590), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n747), .A2(new_n808), .B1(new_n750), .B2(new_n736), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n1015), .A2(new_n1017), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1011), .B1(new_n1024), .B2(new_n722), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n918), .B2(new_n970), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n935), .ZN(new_n1027));
  AOI21_X1  g0827(.A(KEYINPUT113), .B1(new_n1027), .B2(new_n670), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n670), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n935), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1027), .A2(KEYINPUT113), .A3(new_n670), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n942), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n943), .A2(new_n675), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1026), .B1(new_n1032), .B2(new_n714), .C1(new_n1033), .C2(new_n1034), .ZN(G390));
  AOI21_X1  g0835(.A(KEYINPUT39), .B1(new_n872), .B2(new_n850), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n884), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1036), .A2(new_n1037), .B1(new_n883), .B2(new_n890), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n786), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n710), .A2(new_n661), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n889), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n883), .B1(new_n1041), .B2(new_n829), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n873), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1038), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(G330), .B(new_n788), .C1(new_n696), .C2(new_n697), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1045), .A2(new_n886), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1038), .B(new_n1043), .C1(new_n886), .C2(new_n1045), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n715), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n718), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n717), .B1(new_n285), .B2(new_n793), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G68), .A2(new_n756), .B1(new_n751), .B2(G294), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n447), .B2(new_n742), .C1(new_n808), .C2(new_n753), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n274), .B(new_n1053), .C1(G87), .C2(new_n748), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n735), .A2(new_n460), .B1(new_n758), .B2(new_n278), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT118), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1054), .B(new_n1056), .C1(new_n544), .C2(new_n768), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G128), .A2(new_n754), .B1(new_n743), .B2(G137), .ZN(new_n1058));
  INV_X1    g0858(.A(G125), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1058), .B1(new_n1059), .B2(new_n750), .C1(new_n801), .C2(new_n735), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(KEYINPUT54), .B(G143), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1060), .B1(new_n951), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n274), .B1(new_n755), .B2(new_n202), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT117), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n748), .A2(G150), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT53), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G159), .B2(new_n759), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1063), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1057), .A2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1050), .B(new_n1051), .C1(new_n795), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1049), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n894), .A2(new_n897), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n699), .A2(new_n445), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1074), .A2(new_n618), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT114), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n898), .A2(KEYINPUT114), .A3(new_n1075), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n889), .B(new_n1040), .C1(new_n1045), .C2(new_n886), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT115), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n698), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g0882(.A(KEYINPUT115), .B(G330), .C1(new_n696), .C2(new_n697), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1082), .A2(new_n788), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1080), .B1(new_n1084), .B2(new_n886), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(KEYINPUT116), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n888), .A2(new_n889), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1045), .A2(new_n886), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1088), .B1(new_n1089), .B2(new_n1046), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n1085), .B2(KEYINPUT116), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1078), .B(new_n1079), .C1(new_n1087), .C2(new_n1091), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1073), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n676), .B1(new_n1073), .B2(new_n1092), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1072), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(G378));
  NAND2_X1  g0896(.A1(new_n605), .A2(new_n341), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n656), .A2(new_n299), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1097), .B(new_n1098), .Z(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n875), .B2(G330), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n873), .A2(new_n874), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT38), .B1(new_n847), .B2(new_n849), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n854), .A2(new_n855), .A3(new_n852), .ZN(new_n1106));
  OAI21_X1  g0906(.A(KEYINPUT103), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n850), .A2(new_n851), .A3(new_n856), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n830), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(G330), .B(new_n1104), .C1(new_n1109), .C2(KEYINPUT40), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1110), .A2(new_n1101), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n893), .B1(new_n1103), .B2(new_n1111), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n885), .A2(new_n891), .A3(new_n892), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n875), .A2(G330), .A3(new_n1102), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1110), .A2(new_n1101), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1112), .A2(KEYINPUT120), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT120), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1118), .B(new_n893), .C1(new_n1103), .C2(new_n1111), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n898), .A2(KEYINPUT114), .A3(new_n1075), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT114), .B1(new_n898), .B2(new_n1075), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1122), .B1(new_n1073), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1117), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT57), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n676), .B1(new_n1128), .B2(new_n1124), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n793), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n756), .A2(G58), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1132), .B1(new_n278), .B2(new_n747), .C1(new_n808), .C2(new_n750), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n395), .A2(new_n478), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT119), .Z(new_n1136));
  OAI22_X1  g0936(.A1(new_n735), .A2(new_n447), .B1(new_n738), .B2(new_n312), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n753), .A2(new_n460), .B1(new_n742), .B2(new_n507), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1136), .A2(new_n960), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT58), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n753), .A2(new_n1059), .B1(new_n742), .B2(new_n801), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G150), .B2(new_n759), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G137), .A2(new_n764), .B1(new_n748), .B2(new_n1062), .ZN(new_n1145));
  INV_X1    g0945(.A(G128), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1144), .B(new_n1145), .C1(new_n1146), .C2(new_n735), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(G33), .A2(G41), .ZN(new_n1149));
  INV_X1    g0949(.A(G124), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1149), .B1(new_n750), .B2(new_n1150), .C1(new_n770), .C2(new_n755), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n1147), .B2(KEYINPUT59), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1149), .A2(G50), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1148), .A2(new_n1152), .B1(new_n1134), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1142), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n1141), .B2(new_n1140), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n716), .B1(G50), .B2(new_n1131), .C1(new_n1156), .C2(new_n795), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1101), .B2(new_n718), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n715), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1130), .A2(new_n1160), .ZN(G375));
  OAI21_X1  g0961(.A(new_n1123), .B1(new_n1121), .B2(new_n1120), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n930), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n1163), .A3(new_n1092), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n747), .A2(new_n770), .B1(new_n750), .B2(new_n1146), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT122), .Z(new_n1166));
  AOI22_X1  g0966(.A1(new_n762), .A2(G137), .B1(new_n754), .B2(G132), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1167), .B1(new_n797), .B2(new_n738), .C1(new_n742), .C2(new_n1061), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1166), .B(new_n1168), .C1(G50), .C2(new_n759), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1132), .A2(new_n407), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT121), .Z(new_n1171));
  OAI22_X1  g0971(.A1(new_n735), .A2(new_n808), .B1(new_n753), .B2(new_n814), .ZN(new_n1172));
  NOR4_X1   g0972(.A1(new_n1172), .A2(new_n274), .A3(new_n964), .A4(new_n997), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n743), .A2(G116), .B1(new_n751), .B2(G303), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n507), .B2(new_n747), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n951), .B2(G107), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1169), .A2(new_n1171), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n716), .B1(G68), .B2(new_n1131), .C1(new_n1177), .C2(new_n795), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n886), .B2(new_n718), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1085), .A2(KEYINPUT116), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(new_n1086), .A3(new_n1090), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1179), .B1(new_n1181), .B2(new_n715), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1164), .A2(new_n1182), .ZN(G381));
  NOR2_X1   g0983(.A1(G375), .A2(G378), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1026), .B1(new_n1032), .B2(new_n714), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n820), .ZN(new_n1188));
  NOR4_X1   g0988(.A1(new_n1188), .A2(G387), .A3(G396), .A4(G393), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1184), .A2(new_n1182), .A3(new_n1164), .A4(new_n1189), .ZN(G407));
  NAND3_X1  g0990(.A1(new_n658), .A2(new_n659), .A3(G213), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1184), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(G407), .A2(G213), .A3(new_n1193), .ZN(G409));
  AOI21_X1  g0994(.A(G390), .B1(new_n945), .B2(new_n971), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(G387), .A2(new_n1187), .ZN(new_n1196));
  XOR2_X1   g0996(.A(G393), .B(G396), .Z(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OR3_X1    g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1198), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1122), .A2(new_n1181), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n676), .B1(new_n1202), .B2(KEYINPUT60), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1092), .A2(KEYINPUT60), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1204), .A2(new_n1162), .A3(KEYINPUT125), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT125), .B1(new_n1204), .B2(new_n1162), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1182), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n820), .ZN(new_n1209));
  OAI211_X1 g1009(.A(G384), .B(new_n1182), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(KEYINPUT62), .A3(new_n1210), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1117), .A2(new_n1163), .A3(new_n1119), .A4(new_n1124), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1158), .B1(new_n1213), .B2(new_n715), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT123), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(new_n1216), .A3(new_n1095), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1216), .B1(new_n1215), .B2(new_n1095), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1130), .A2(new_n1160), .A3(G378), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1192), .B(new_n1211), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1215), .A2(new_n1095), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT123), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1221), .A2(new_n1224), .A3(new_n1217), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT124), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT124), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1221), .A2(new_n1224), .A3(new_n1228), .A4(new_n1217), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1226), .A2(new_n1191), .A3(new_n1227), .A4(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT62), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1222), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT61), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1192), .A2(G2897), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1227), .B(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1192), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1233), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1201), .B1(new_n1232), .B2(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1227), .A2(KEYINPUT63), .ZN(new_n1239));
  AOI211_X1 g1039(.A(KEYINPUT61), .B(new_n1201), .C1(new_n1236), .C2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT63), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1226), .A2(new_n1191), .A3(new_n1229), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1234), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1227), .B(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1241), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1230), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1240), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1238), .A2(new_n1247), .ZN(G405));
  INV_X1    g1048(.A(KEYINPUT126), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1201), .A2(new_n1249), .A3(new_n1227), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1227), .A2(new_n1249), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(G375), .B(G378), .ZN(new_n1254));
  XOR2_X1   g1054(.A(new_n1253), .B(new_n1254), .Z(G402));
endmodule


