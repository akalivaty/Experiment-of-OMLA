//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n540, new_n542, new_n543, new_n544,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n564, new_n565, new_n566, new_n567, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n599, new_n600, new_n601, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1205, new_n1206, new_n1207, new_n1208;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT64), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n464), .A2(new_n469), .ZN(G160));
  NOR2_X1   g045(.A1(new_n460), .A2(new_n461), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(new_n459), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n471), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G162));
  OAI21_X1  g054(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n482));
  INV_X1    g057(.A(G114), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n482), .A2(new_n483), .A3(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT65), .B1(new_n459), .B2(G114), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n490), .B(new_n492), .C1(new_n461), .C2(new_n460), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n490), .B1(new_n460), .B2(new_n461), .ZN(new_n494));
  INV_X1    g069(.A(new_n492), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n488), .B1(new_n493), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G50), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  OR2_X1    g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT5), .B(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G88), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n498), .A2(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n506), .A2(new_n509), .ZN(G303));
  INV_X1    g085(.A(G303), .ZN(G166));
  NAND3_X1  g086(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT7), .ZN(new_n513));
  INV_X1    g088(.A(G89), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n504), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT67), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT67), .ZN(new_n517));
  OAI211_X1 g092(.A(new_n517), .B(new_n513), .C1(new_n504), .C2(new_n514), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n499), .A2(new_n500), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(G63), .A2(G651), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n521), .A2(G51), .B1(new_n503), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n516), .A2(new_n518), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(G168));
  XOR2_X1   g100(.A(KEYINPUT69), .B(G90), .Z(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT68), .B(G52), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n504), .A2(new_n526), .B1(new_n502), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n508), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n528), .A2(new_n530), .ZN(G171));
  XOR2_X1   g106(.A(KEYINPUT5), .B(G543), .Z(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n519), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT70), .B(G81), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n533), .A2(new_n534), .B1(new_n521), .B2(G43), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n508), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  NAND4_X1  g114(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT71), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT72), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  INV_X1    g120(.A(G53), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT9), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n502), .A2(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g126(.A(new_n521), .B(G53), .C1(new_n547), .C2(new_n548), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n551), .A2(KEYINPUT74), .A3(new_n552), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n532), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G651), .B1(new_n533), .B2(G91), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  NAND2_X1  g138(.A1(new_n524), .A2(KEYINPUT75), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n516), .A2(new_n565), .A3(new_n518), .A4(new_n523), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G286));
  OR2_X1    g143(.A1(new_n503), .A2(G74), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(new_n521), .B2(G49), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n571));
  AND3_X1   g146(.A1(new_n533), .A2(new_n571), .A3(G87), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n571), .B1(new_n533), .B2(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(G288));
  AOI22_X1  g149(.A1(new_n503), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n508), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n533), .A2(G86), .B1(new_n521), .B2(G48), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G305));
  INV_X1    g154(.A(G47), .ZN(new_n580));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  OAI22_X1  g156(.A1(new_n580), .A2(new_n502), .B1(new_n504), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n508), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n533), .A2(G92), .ZN(new_n588));
  XOR2_X1   g163(.A(new_n588), .B(KEYINPUT10), .Z(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n532), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(new_n521), .B2(G54), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n587), .B1(new_n594), .B2(G868), .ZN(G284));
  OAI21_X1  g170(.A(new_n587), .B1(new_n594), .B2(G868), .ZN(G321));
  INV_X1    g171(.A(new_n561), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n555), .B2(new_n556), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT77), .B1(new_n598), .B2(G868), .ZN(new_n599));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n567), .A2(new_n600), .ZN(new_n601));
  MUX2_X1   g176(.A(new_n599), .B(KEYINPUT77), .S(new_n601), .Z(G297));
  MUX2_X1   g177(.A(new_n599), .B(KEYINPUT77), .S(new_n601), .Z(G280));
  XNOR2_X1  g178(.A(KEYINPUT78), .B(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n594), .B1(G860), .B2(new_n604), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT79), .Z(G148));
  NAND2_X1  g181(.A1(new_n537), .A2(new_n600), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n594), .A2(new_n604), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n609), .B2(new_n600), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n472), .A2(G123), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n474), .A2(G135), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n459), .A2(G111), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT80), .Z(new_n617));
  OR2_X1    g192(.A1(new_n617), .A2(G2096), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT3), .B(G2104), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n467), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n617), .A2(G2096), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n618), .A2(new_n623), .A3(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2443), .B(G2446), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n633), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT82), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n637), .A2(new_n639), .ZN(new_n642));
  AND2_X1   g217(.A1(new_n642), .A2(G14), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n641), .A2(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT83), .ZN(new_n646));
  NOR2_X1   g221(.A1(G2072), .A2(G2078), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n442), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT17), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT84), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n648), .ZN(new_n653));
  AOI211_X1 g228(.A(new_n646), .B(new_n652), .C1(new_n653), .C2(new_n651), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n646), .A2(new_n648), .A3(new_n650), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n649), .A2(new_n651), .A3(new_n646), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT85), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2096), .B(G2100), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT85), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n660), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n662), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n663), .A2(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n672), .B(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n677), .A2(KEYINPUT87), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n675), .B(new_n678), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n674), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT86), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n680), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(KEYINPUT20), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n679), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1991), .B(G1996), .Z(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n691), .B2(new_n692), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G19), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n538), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT92), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1341), .ZN(new_n703));
  NOR2_X1   g278(.A1(G4), .A2(G16), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT91), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n589), .A2(new_n593), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n699), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1348), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G26), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n472), .A2(G128), .ZN(new_n712));
  INV_X1    g287(.A(G140), .ZN(new_n713));
  INV_X1    g288(.A(new_n474), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G104), .ZN(new_n716));
  AND3_X1   g291(.A1(new_n716), .A2(new_n459), .A3(KEYINPUT93), .ZN(new_n717));
  AOI21_X1  g292(.A(KEYINPUT93), .B1(new_n716), .B2(new_n459), .ZN(new_n718));
  OAI221_X1 g293(.A(G2104), .B1(G116), .B2(new_n459), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n711), .B1(new_n721), .B2(new_n709), .ZN(new_n722));
  INV_X1    g297(.A(G2067), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n708), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n703), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT94), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n699), .A2(G20), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT23), .Z(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G299), .B2(G16), .ZN(new_n730));
  INV_X1    g305(.A(G1956), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n709), .A2(G35), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G162), .B2(new_n709), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT29), .Z(new_n735));
  INV_X1    g310(.A(G2090), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n699), .A2(G21), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G168), .B2(new_n699), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n737), .B1(G1966), .B2(new_n739), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n732), .B(new_n740), .C1(G1966), .C2(new_n739), .ZN(new_n741));
  NOR2_X1   g316(.A1(G171), .A2(new_n699), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G5), .B2(new_n699), .ZN(new_n743));
  INV_X1    g318(.A(G1961), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(KEYINPUT24), .A2(G34), .ZN(new_n746));
  NOR2_X1   g321(.A1(KEYINPUT24), .A2(G34), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n709), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT96), .Z(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G29), .B2(G160), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n745), .B1(G2084), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n709), .A2(G32), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT26), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G129), .B2(new_n472), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n474), .A2(G141), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n467), .A2(G105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT97), .ZN(new_n758));
  AND3_X1   g333(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(KEYINPUT98), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(KEYINPUT98), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n752), .B1(new_n762), .B2(new_n709), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT27), .B(G1996), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n751), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT99), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n709), .A2(G33), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n474), .A2(G139), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT95), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n619), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(new_n459), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n768), .B1(new_n776), .B2(new_n709), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2072), .ZN(new_n778));
  OAI22_X1  g353(.A1(new_n763), .A2(new_n765), .B1(new_n735), .B2(new_n736), .ZN(new_n779));
  INV_X1    g354(.A(new_n617), .ZN(new_n780));
  INV_X1    g355(.A(G2078), .ZN(new_n781));
  NOR2_X1   g356(.A1(G164), .A2(new_n709), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G27), .B2(new_n709), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n780), .A2(G29), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n743), .A2(new_n744), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT30), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n786), .A2(G28), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n709), .B1(new_n786), .B2(G28), .ZN(new_n788));
  AND2_X1   g363(.A1(KEYINPUT31), .A2(G11), .ZN(new_n789));
  NOR2_X1   g364(.A1(KEYINPUT31), .A2(G11), .ZN(new_n790));
  OAI22_X1  g365(.A1(new_n787), .A2(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n750), .B2(G2084), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n783), .A2(new_n781), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n784), .A2(new_n785), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n778), .A2(new_n779), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n741), .A2(new_n767), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n727), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(G6), .A2(G16), .ZN(new_n799));
  INV_X1    g374(.A(G305), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G16), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT32), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1981), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n699), .A2(G22), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G166), .B2(new_n699), .ZN(new_n805));
  INV_X1    g380(.A(G1971), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(G16), .A2(G23), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT88), .Z(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G288), .B2(new_n699), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT33), .B(G1976), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n807), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  OR3_X1    g389(.A1(new_n803), .A2(new_n814), .A3(KEYINPUT89), .ZN(new_n815));
  OAI21_X1  g390(.A(KEYINPUT89), .B1(new_n803), .B2(new_n814), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n815), .A2(new_n816), .A3(KEYINPUT34), .ZN(new_n820));
  NOR2_X1   g395(.A1(G16), .A2(G24), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n585), .B2(G16), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(G1986), .Z(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(KEYINPUT90), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n472), .A2(G119), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n474), .A2(G131), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n459), .A2(G107), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n826), .B(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  MUX2_X1   g405(.A(G25), .B(new_n830), .S(G29), .Z(new_n831));
  XOR2_X1   g406(.A(KEYINPUT35), .B(G1991), .Z(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n831), .B(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n825), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n819), .A2(new_n820), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n824), .A2(KEYINPUT90), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n838), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n798), .B1(new_n839), .B2(new_n840), .ZN(G311));
  AND2_X1   g416(.A1(new_n836), .A2(new_n838), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n836), .A2(new_n838), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n797), .B1(new_n842), .B2(new_n843), .ZN(G150));
  NAND2_X1  g419(.A1(new_n594), .A2(G559), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT100), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  INV_X1    g422(.A(G55), .ZN(new_n848));
  INV_X1    g423(.A(G93), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n848), .A2(new_n502), .B1(new_n504), .B2(new_n849), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n508), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n537), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n847), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n856));
  AOI21_X1  g431(.A(G860), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n856), .B2(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n853), .A2(G860), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT37), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(G145));
  AND2_X1   g436(.A1(new_n465), .A2(new_n468), .ZN(new_n862));
  INV_X1    g437(.A(G125), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT3), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n466), .ZN(new_n865));
  NAND2_X1  g440(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n863), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n463), .ZN(new_n868));
  OAI21_X1  g443(.A(G2105), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n617), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(G162), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n762), .A2(new_n721), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n760), .A2(new_n761), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n874), .A2(new_n720), .A3(new_n715), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n472), .A2(G130), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT102), .ZN(new_n878));
  OAI21_X1  g453(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n879));
  INV_X1    g454(.A(G118), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(new_n880), .B2(G2105), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(new_n474), .B2(G142), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n876), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n488), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n496), .A2(new_n493), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n486), .A2(KEYINPUT101), .A3(new_n487), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n776), .B(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n830), .B(new_n621), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n883), .B1(new_n873), .B2(new_n875), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n773), .A2(new_n775), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n896), .A2(new_n890), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n890), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n892), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AND4_X1   g474(.A1(new_n885), .A2(new_n894), .A3(new_n895), .A4(new_n899), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n885), .A2(new_n895), .B1(new_n899), .B2(new_n894), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n872), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI211_X1 g479(.A(KEYINPUT103), .B(new_n872), .C1(new_n900), .C2(new_n901), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n900), .A2(new_n901), .A3(new_n872), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n907), .A2(G37), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n906), .A2(new_n908), .A3(KEYINPUT40), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT40), .B1(new_n906), .B2(new_n908), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(G395));
  XNOR2_X1  g486(.A(G303), .B(new_n585), .ZN(new_n912));
  XNOR2_X1  g487(.A(G288), .B(G305), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n912), .B(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n594), .A2(new_n598), .ZN(new_n916));
  NAND2_X1  g491(.A1(G299), .A2(new_n706), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(KEYINPUT41), .A3(new_n917), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n850), .A2(new_n852), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(new_n537), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n854), .A2(KEYINPUT104), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n609), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n854), .A2(KEYINPUT104), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n924), .A2(new_n925), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n608), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n922), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n928), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n918), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n915), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(new_n934), .A3(new_n915), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n914), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n937), .ZN(new_n939));
  INV_X1    g514(.A(new_n914), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n939), .A2(new_n940), .A3(new_n935), .ZN(new_n941));
  OAI21_X1  g516(.A(G868), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n923), .A2(G868), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n936), .A2(new_n914), .A3(new_n937), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n940), .B1(new_n939), .B2(new_n935), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n600), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT105), .B1(new_n949), .B2(new_n944), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n946), .A2(new_n950), .ZN(G295));
  NAND2_X1  g526(.A1(new_n942), .A2(new_n945), .ZN(G331));
  AOI21_X1  g527(.A(G301), .B1(new_n564), .B2(new_n566), .ZN(new_n953));
  NOR2_X1   g528(.A1(G168), .A2(G171), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n953), .A2(new_n924), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n924), .B1(new_n953), .B2(new_n954), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n920), .A2(new_n956), .A3(new_n921), .A4(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n957), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n917), .B(new_n916), .C1(new_n959), .C2(new_n955), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(new_n960), .A3(new_n940), .ZN(new_n961));
  INV_X1    g536(.A(G37), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n958), .A2(new_n960), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n966), .A2(KEYINPUT107), .A3(new_n914), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT107), .B1(new_n966), .B2(new_n914), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n964), .B(new_n965), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n940), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n958), .A2(new_n960), .A3(KEYINPUT106), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n963), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n969), .B(KEYINPUT108), .C1(new_n973), .C2(new_n965), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n967), .A2(new_n968), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n976), .A2(new_n977), .A3(new_n965), .A4(new_n964), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n974), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n964), .B(KEYINPUT43), .C1(new_n967), .C2(new_n968), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(KEYINPUT43), .B2(new_n973), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT44), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n982), .ZN(G397));
  AOI21_X1  g558(.A(KEYINPUT109), .B1(G160), .B2(G40), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n985));
  INV_X1    g560(.A(G40), .ZN(new_n986));
  NOR4_X1   g561(.A1(new_n464), .A2(new_n469), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT45), .B1(new_n890), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1996), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n874), .B(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n721), .B(G2067), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n830), .A2(new_n833), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n830), .A2(new_n833), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  XOR2_X1   g573(.A(new_n585), .B(G1986), .Z(new_n999));
  OAI21_X1  g574(.A(new_n992), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n985), .B1(new_n870), .B2(new_n986), .ZN(new_n1002));
  NAND3_X1  g577(.A1(G160), .A2(KEYINPUT109), .A3(G40), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n888), .A2(new_n889), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT101), .B1(new_n486), .B2(new_n487), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n989), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n486), .A2(new_n487), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1384), .B1(new_n888), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1004), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(G1961), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT110), .B1(new_n1011), .B2(KEYINPUT45), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1016), .B(new_n1017), .C1(G164), .C2(G1384), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n890), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1019), .A2(new_n781), .A3(new_n988), .A4(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT123), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1014), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1021), .A2(KEYINPUT123), .A3(new_n1022), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1007), .A2(new_n1017), .ZN(new_n1027));
  NOR4_X1   g602(.A1(new_n870), .A2(new_n1022), .A3(new_n986), .A4(G2078), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1020), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1025), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1001), .B1(new_n1030), .B2(G171), .ZN(new_n1031));
  INV_X1    g606(.A(new_n493), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n492), .B1(new_n619), .B2(new_n490), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT45), .B(new_n989), .C1(new_n1034), .C2(new_n488), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1027), .A2(new_n988), .A3(new_n781), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT122), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1002), .A2(new_n1035), .A3(new_n1003), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT122), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1039), .A2(new_n1040), .A3(new_n781), .A4(new_n1027), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(new_n1041), .A3(KEYINPUT53), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1025), .A2(G301), .A3(new_n1026), .A4(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1043), .A2(KEYINPUT124), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(KEYINPUT124), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1031), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1014), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n1042), .A3(new_n1026), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G171), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(G171), .B2(new_n1030), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1001), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1004), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1971), .B1(new_n1053), .B2(new_n1020), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT50), .B1(new_n890), .B2(new_n989), .ZN(new_n1055));
  NOR3_X1   g630(.A1(G164), .A2(new_n1008), .A3(G1384), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n988), .B(new_n736), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT111), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1019), .A2(new_n988), .A3(new_n1020), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1060), .B(new_n1057), .C1(new_n1061), .C2(G1971), .ZN(new_n1062));
  NAND2_X1  g637(.A1(G303), .A2(G8), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT55), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1059), .A2(new_n1062), .A3(G8), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1011), .A2(new_n1008), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1008), .B1(new_n890), .B2(new_n989), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1068), .A2(G2090), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(G8), .B1(new_n1054), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n1064), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n1073));
  NOR2_X1   g648(.A1(G305), .A2(G1981), .ZN(new_n1074));
  INV_X1    g649(.A(G1981), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n577), .B2(new_n578), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1073), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT49), .ZN(new_n1078));
  INV_X1    g653(.A(G8), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1007), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1079), .B1(new_n988), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT49), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1073), .B(new_n1082), .C1(new_n1074), .C2(new_n1076), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1078), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G288), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(G1976), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1081), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT52), .ZN(new_n1088));
  INV_X1    g663(.A(G1976), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT52), .B1(G288), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1081), .A2(new_n1086), .A3(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1084), .A2(new_n1088), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1066), .A2(new_n1072), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n1095));
  INV_X1    g670(.A(G1966), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1038), .B2(new_n990), .ZN(new_n1097));
  INV_X1    g672(.A(G2084), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n988), .B(new_n1098), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1095), .B(G8), .C1(new_n1100), .C2(new_n524), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n524), .A2(G8), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g680(.A(KEYINPUT120), .B(new_n1102), .C1(new_n1097), .C2(new_n1099), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1101), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1100), .A2(G8), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(KEYINPUT51), .A3(new_n1102), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1094), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1103), .B(new_n1104), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1112), .A2(KEYINPUT121), .A3(new_n1109), .A4(new_n1101), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1093), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1046), .A2(new_n1052), .A3(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1061), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n731), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1118), .A2(KEYINPUT114), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT114), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1120), .B(new_n731), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1117), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n553), .A2(new_n1124), .A3(new_n561), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n598), .B2(new_n1124), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(KEYINPUT115), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1013), .A2(G1348), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n988), .A2(new_n1080), .A3(new_n723), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1128), .B1(new_n706), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1126), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1133), .B(new_n1117), .C1(new_n1119), .C2(new_n1122), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1118), .A2(KEYINPUT114), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1136), .A2(new_n1121), .B1(new_n1061), .B2(new_n1116), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT115), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1126), .B(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1134), .B(KEYINPUT61), .C1(new_n1137), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1128), .A2(KEYINPUT118), .A3(KEYINPUT61), .A4(new_n1134), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1129), .A2(KEYINPUT60), .A3(new_n1130), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1145), .A2(KEYINPUT119), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1145), .A2(KEYINPUT119), .A3(new_n706), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n706), .B1(new_n1145), .B2(KEYINPUT119), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1131), .A2(KEYINPUT60), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1134), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n1154));
  NAND2_X1  g729(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1053), .A2(new_n993), .A3(new_n1020), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT116), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT58), .B(G1341), .Z(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1157), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n538), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1153), .A2(new_n1154), .B1(new_n1155), .B2(new_n1162), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1162), .A2(new_n1155), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1144), .A2(new_n1151), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1115), .B1(new_n1135), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(KEYINPUT62), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1111), .A2(new_n1113), .A3(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1093), .A2(new_n1050), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  XOR2_X1   g747(.A(KEYINPUT113), .B(KEYINPUT63), .Z(new_n1173));
  NAND3_X1  g748(.A1(new_n1100), .A2(G8), .A3(new_n567), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1173), .B1(new_n1093), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1066), .A2(new_n1092), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1174), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1059), .A2(G8), .A3(new_n1062), .ZN(new_n1178));
  OAI211_X1 g753(.A(KEYINPUT63), .B(new_n1177), .C1(new_n1178), .C2(new_n1065), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1175), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1066), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1084), .A2(new_n1089), .A3(new_n1085), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(G1981), .B2(G305), .ZN(new_n1183));
  AOI22_X1  g758(.A1(new_n1181), .A2(new_n1092), .B1(new_n1183), .B2(new_n1081), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1172), .A2(new_n1180), .A3(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1000), .B1(new_n1166), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n991), .A2(G1996), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(KEYINPUT46), .ZN(new_n1188));
  XOR2_X1   g763(.A(new_n1188), .B(KEYINPUT125), .Z(new_n1189));
  AOI21_X1  g764(.A(new_n991), .B1(new_n762), .B2(new_n995), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT126), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1189), .B(new_n1191), .C1(KEYINPUT46), .C2(new_n1187), .ZN(new_n1192));
  XOR2_X1   g767(.A(new_n1192), .B(KEYINPUT47), .Z(new_n1193));
  NAND2_X1  g768(.A1(new_n998), .A2(new_n992), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT127), .ZN(new_n1195));
  NOR3_X1   g770(.A1(new_n991), .A2(G1986), .A3(G290), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT48), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n994), .A2(new_n995), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1198), .A2(new_n996), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1199), .B1(new_n723), .B2(new_n721), .ZN(new_n1200));
  OAI22_X1  g775(.A1(new_n1195), .A2(new_n1197), .B1(new_n991), .B2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1193), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1186), .A2(new_n1202), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g778(.A1(new_n663), .A2(new_n667), .A3(G319), .ZN(new_n1205));
  AOI21_X1  g779(.A(new_n1205), .B1(new_n641), .B2(new_n643), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n1206), .A2(new_n697), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n1207), .B1(new_n906), .B2(new_n908), .ZN(new_n1208));
  AND3_X1   g782(.A1(new_n1208), .A2(new_n974), .A3(new_n978), .ZN(G308));
  NAND3_X1  g783(.A1(new_n1208), .A2(new_n974), .A3(new_n978), .ZN(G225));
endmodule


