//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT73), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n202), .A2(KEYINPUT73), .ZN(new_n204));
  INV_X1    g003(.A(G183gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT27), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT27), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G183gat), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT28), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT27), .B(G183gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT28), .A3(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n218));
  INV_X1    g017(.A(G169gat), .ZN(new_n219));
  INV_X1    g018(.A(G176gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT26), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n217), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n215), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n228), .A3(KEYINPUT68), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G113gat), .B2(G120gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G127gat), .B(G134gat), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT70), .B(G113gat), .Z(new_n238));
  INV_X1    g037(.A(G120gat), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n236), .B(new_n237), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G113gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n239), .ZN(new_n242));
  NAND2_X1  g041(.A1(G113gat), .A2(G120gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n234), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n245));
  INV_X1    g044(.A(G134gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G127gat), .ZN(new_n247));
  INV_X1    g046(.A(G127gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(G134gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n244), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n245), .B1(new_n244), .B2(new_n250), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n240), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT71), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n243), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n235), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT69), .B1(new_n257), .B2(new_n237), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n244), .A2(new_n245), .A3(new_n250), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(KEYINPUT71), .A3(new_n240), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n216), .ZN(new_n263));
  NAND4_X1  g062(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n263), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n219), .A2(new_n220), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n226), .B1(new_n270), .B2(KEYINPUT23), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT23), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(KEYINPUT66), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n269), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g073(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n272), .A2(G169gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n268), .A2(new_n274), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT25), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n270), .A2(KEYINPUT23), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n272), .A2(KEYINPUT66), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(new_n226), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n281), .B1(new_n285), .B2(new_n269), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n221), .A2(KEYINPUT23), .A3(new_n223), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n263), .A2(new_n265), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n233), .A2(new_n255), .A3(new_n261), .A4(new_n290), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n215), .A2(KEYINPUT68), .A3(new_n228), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT68), .B1(new_n215), .B2(new_n228), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n285), .A2(new_n269), .B1(new_n277), .B2(new_n278), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT25), .B1(new_n294), .B2(new_n268), .ZN(new_n295));
  AND4_X1   g094(.A1(KEYINPUT25), .A2(new_n274), .A3(new_n287), .A4(new_n288), .ZN(new_n296));
  OAI22_X1  g095(.A1(new_n292), .A2(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n255), .A2(new_n261), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G227gat), .ZN(new_n300));
  INV_X1    g099(.A(G233gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n291), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n304), .B(KEYINPUT34), .Z(new_n305));
  XOR2_X1   g104(.A(G71gat), .B(G99gat), .Z(new_n306));
  XNOR2_X1  g105(.A(G15gat), .B(G43gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n303), .B1(new_n291), .B2(new_n299), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT33), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(KEYINPUT32), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n308), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n297), .A2(new_n298), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n233), .A2(new_n290), .B1(new_n255), .B2(new_n261), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n302), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n308), .A2(KEYINPUT33), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT32), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n315), .A2(KEYINPUT72), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n309), .B2(new_n317), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n305), .B1(new_n312), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT72), .B1(new_n315), .B2(new_n318), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n309), .A2(new_n320), .A3(new_n317), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n312), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n304), .B(KEYINPUT34), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n203), .B(new_n204), .C1(new_n323), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n326), .A2(new_n327), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n305), .A2(new_n322), .A3(new_n312), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT73), .A4(new_n202), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G228gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(new_n301), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336));
  XNOR2_X1  g135(.A(G197gat), .B(G204gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT22), .ZN(new_n338));
  INV_X1    g137(.A(G211gat), .ZN(new_n339));
  INV_X1    g138(.A(G218gat), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G211gat), .B(G218gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n336), .B1(new_n344), .B2(KEYINPUT29), .ZN(new_n345));
  AND2_X1   g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G141gat), .B(G148gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT2), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n350), .B1(G155gat), .B2(G162gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n348), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G141gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G148gat), .ZN(new_n354));
  INV_X1    g153(.A(G148gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G141gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G155gat), .B(G162gat), .ZN(new_n358));
  INV_X1    g157(.A(G155gat), .ZN(new_n359));
  INV_X1    g158(.A(G162gat), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT2), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n357), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n352), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n363), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n352), .A2(new_n362), .A3(new_n336), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n344), .B1(new_n365), .B2(KEYINPUT29), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n366), .A3(G22gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(G22gat), .B1(new_n364), .B2(new_n366), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n335), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n364), .A2(new_n366), .ZN(new_n371));
  INV_X1    g170(.A(G22gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n335), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n374), .A3(new_n367), .ZN(new_n375));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT31), .B(G50gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  AND2_X1   g177(.A1(new_n378), .A2(KEYINPUT79), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n370), .A2(new_n375), .A3(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n378), .A2(KEYINPUT79), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n383), .B1(new_n370), .B2(new_n375), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n282), .A2(new_n289), .B1(new_n215), .B2(new_n228), .ZN(new_n387));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n388), .B(KEYINPUT74), .Z(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT75), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT75), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n295), .A2(new_n296), .ZN(new_n393));
  INV_X1    g192(.A(new_n229), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n392), .B(new_n389), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT29), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n389), .B1(new_n297), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n344), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n297), .A2(new_n389), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n390), .B1(new_n387), .B2(KEYINPUT29), .ZN(new_n401));
  INV_X1    g200(.A(new_n344), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  AND3_X1   g205(.A1(new_n399), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(KEYINPUT76), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n408), .B1(new_n399), .B2(new_n403), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT30), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n399), .A2(new_n403), .A3(new_n406), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n298), .B2(new_n363), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT5), .ZN(new_n417));
  NAND2_X1  g216(.A1(G225gat), .A2(G233gat), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n336), .B1(new_n352), .B2(new_n362), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n365), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n419), .B1(new_n421), .B2(new_n253), .ZN(new_n422));
  INV_X1    g221(.A(new_n363), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(new_n260), .A3(new_n240), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n424), .A2(new_n415), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n416), .A2(new_n417), .A3(new_n422), .A4(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n255), .A2(KEYINPUT4), .A3(new_n423), .A4(new_n261), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n424), .A2(new_n415), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n422), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT77), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n253), .A2(new_n363), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n424), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n417), .B1(new_n432), .B2(new_n419), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n429), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n430), .B1(new_n429), .B2(new_n433), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n426), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(G1gat), .B(G29gat), .Z(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G57gat), .B(G85gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n436), .A2(KEYINPUT6), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT6), .B1(new_n436), .B2(new_n442), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n441), .B(new_n426), .C1(new_n434), .C2(new_n435), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n414), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n333), .B1(new_n386), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n444), .A2(KEYINPUT82), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n443), .B1(new_n446), .B2(new_n445), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(KEYINPUT82), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n399), .A2(new_n403), .ZN(new_n454));
  XOR2_X1   g253(.A(KEYINPUT81), .B(KEYINPUT37), .Z(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n406), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT37), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT38), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n408), .A2(KEYINPUT38), .ZN(new_n462));
  OR3_X1    g261(.A1(new_n396), .A2(new_n398), .A3(new_n344), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n400), .A2(new_n401), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n344), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n463), .A2(KEYINPUT80), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT37), .B1(new_n463), .B2(KEYINPUT80), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n456), .B(new_n462), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n461), .A2(new_n411), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n421), .A2(new_n253), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n416), .A2(new_n471), .A3(new_n425), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n419), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n473), .A2(KEYINPUT39), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n473), .B(KEYINPUT39), .C1(new_n419), .C2(new_n432), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n475), .A3(new_n441), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT40), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n436), .A2(new_n442), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n476), .A2(new_n477), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n414), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n385), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n450), .B1(new_n470), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n330), .A2(new_n385), .A3(new_n331), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT83), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT83), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n330), .A2(new_n331), .A3(new_n385), .A4(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n448), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT35), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT35), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n410), .A2(new_n491), .A3(new_n413), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n453), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n484), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g295(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n498));
  AOI21_X1  g297(.A(G36gat), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G29gat), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n500), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(KEYINPUT85), .ZN(new_n503));
  AND2_X1   g302(.A1(G43gat), .A2(G50gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(G43gat), .A2(G50gat), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT15), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n503), .B(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT86), .B(G43gat), .ZN(new_n508));
  INV_X1    g307(.A(G50gat), .ZN(new_n509));
  AOI211_X1 g308(.A(KEYINPUT15), .B(new_n504), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(new_n499), .B2(new_n501), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT87), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n512), .A2(new_n513), .ZN(new_n516));
  XNOR2_X1  g315(.A(G15gat), .B(G22gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(KEYINPUT88), .ZN(new_n518));
  INV_X1    g317(.A(G1gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n519), .A2(KEYINPUT16), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G8gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n515), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G229gat), .A2(G233gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n523), .B(KEYINPUT89), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n512), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT18), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n525), .A2(KEYINPUT18), .A3(new_n526), .A4(new_n528), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n526), .B(KEYINPUT13), .Z(new_n533));
  INV_X1    g332(.A(new_n528), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n527), .A2(new_n512), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n531), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(G169gat), .B(G197gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n542), .B(KEYINPUT12), .Z(new_n543));
  NAND2_X1  g342(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n543), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n531), .A2(new_n532), .A3(new_n536), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n496), .A2(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n549), .B(KEYINPUT90), .Z(new_n550));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n551), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(G71gat), .B2(G78gat), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n554));
  AND2_X1   g353(.A1(G57gat), .A2(G64gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(G57gat), .A2(G64gat), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n553), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT21), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n527), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT94), .ZN(new_n562));
  XOR2_X1   g361(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT93), .ZN(new_n564));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT92), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n564), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n562), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n558), .A2(new_n559), .ZN(new_n569));
  XOR2_X1   g368(.A(G127gat), .B(G155gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G183gat), .B(G211gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n568), .A2(new_n573), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT7), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT97), .B1(new_n577), .B2(KEYINPUT96), .ZN(new_n578));
  INV_X1    g377(.A(G85gat), .ZN(new_n579));
  INV_X1    g378(.A(G92gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n578), .B(new_n581), .C1(KEYINPUT97), .C2(new_n577), .ZN(new_n582));
  OAI221_X1 g381(.A(KEYINPUT97), .B1(new_n577), .B2(KEYINPUT96), .C1(new_n579), .C2(new_n580), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(KEYINPUT8), .A2(new_n584), .B1(new_n579), .B2(new_n580), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G99gat), .B(G106gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n516), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n515), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n512), .A2(new_n588), .B1(KEYINPUT41), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(G190gat), .B(G218gat), .Z(new_n594));
  OR2_X1    g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT95), .ZN(new_n599));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n595), .A2(new_n601), .A3(new_n596), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G120gat), .B(G148gat), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT99), .ZN(new_n608));
  XNOR2_X1  g407(.A(G176gat), .B(G204gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT101), .ZN(new_n611));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n558), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n588), .B(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n615), .A2(KEYINPUT10), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n588), .A2(new_n614), .A3(KEYINPUT10), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n615), .A2(new_n613), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n611), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n618), .ZN(new_n621));
  INV_X1    g420(.A(new_n610), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n622), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n621), .B(new_n624), .C1(new_n623), .C2(new_n619), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n625), .A2(KEYINPUT100), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(KEYINPUT100), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n620), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n576), .A2(new_n606), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n550), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n452), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT102), .B(G1gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(G1324gat));
  XOR2_X1   g434(.A(KEYINPUT16), .B(G8gat), .Z(new_n636));
  AND3_X1   g435(.A1(new_n632), .A2(new_n414), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(G8gat), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n638), .B1(new_n632), .B2(new_n414), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT42), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(KEYINPUT42), .B2(new_n637), .ZN(G1325gat));
  INV_X1    g440(.A(G15gat), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n323), .A2(new_n328), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n632), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n632), .A2(new_n333), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n644), .B1(new_n645), .B2(new_n642), .ZN(G1326gat));
  NAND2_X1  g445(.A1(new_n632), .A2(new_n386), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT43), .B(G22gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(G1327gat));
  NOR3_X1   g448(.A1(new_n576), .A2(new_n606), .A3(new_n628), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT103), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n550), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n444), .A2(new_n447), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n652), .A2(G29gat), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT45), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  AOI221_X4 g455(.A(KEYINPUT104), .B1(new_n453), .B2(new_n493), .C1(new_n489), .C2(KEYINPUT35), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n658), .B1(new_n490), .B2(new_n494), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n484), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT105), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n662), .B(new_n484), .C1(new_n657), .C2(new_n659), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n606), .A2(KEYINPUT44), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT44), .B1(new_n496), .B2(new_n606), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n576), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(new_n547), .A3(new_n629), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(G29gat), .B1(new_n671), .B2(new_n653), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n672), .ZN(G1328gat));
  NOR3_X1   g472(.A1(new_n652), .A2(G36gat), .A3(new_n482), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT46), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G36gat), .B1(new_n671), .B2(new_n482), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(G1329gat));
  INV_X1    g478(.A(new_n643), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n508), .B1(new_n652), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n333), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(new_n508), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n681), .B1(new_n671), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT47), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT47), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n681), .B(new_n686), .C1(new_n671), .C2(new_n683), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(G1330gat));
  NAND2_X1  g487(.A1(new_n386), .A2(new_n509), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT107), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n550), .A2(new_n651), .A3(new_n690), .ZN(new_n691));
  AOI211_X1 g490(.A(new_n385), .B(new_n669), .C1(new_n665), .C2(new_n666), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n691), .B(KEYINPUT48), .C1(new_n509), .C2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT106), .B1(new_n692), .B2(new_n509), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n667), .A2(new_n386), .A3(new_n670), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n696), .A3(G50gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n694), .A2(new_n697), .A3(new_n691), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT48), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n699), .B1(new_n698), .B2(new_n700), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n693), .B1(new_n701), .B2(new_n702), .ZN(G1331gat));
  NOR2_X1   g502(.A1(new_n668), .A2(new_n605), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n547), .A2(new_n629), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n661), .A2(new_n704), .A3(new_n663), .A4(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n653), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT109), .B(G57gat), .Z(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1332gat));
  NOR2_X1   g508(.A1(new_n706), .A2(new_n482), .ZN(new_n710));
  NOR2_X1   g509(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n711));
  AND2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n710), .B2(new_n711), .ZN(G1333gat));
  OAI21_X1  g513(.A(G71gat), .B1(new_n706), .B2(new_n682), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n680), .A2(G71gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(new_n706), .B2(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g517(.A1(new_n706), .A2(new_n385), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(G78gat), .Z(G1335gat));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(KEYINPUT51), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n576), .A2(new_n606), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n548), .A3(new_n660), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n721), .A2(KEYINPUT51), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n629), .B1(new_n724), .B2(new_n725), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(new_n579), .A3(new_n452), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n667), .A2(new_n668), .A3(new_n705), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n730), .A2(new_n452), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n731), .B2(new_n579), .ZN(G1336gat));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n414), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n482), .A2(G92gat), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n733), .A2(G92gat), .B1(new_n728), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1337gat));
  INV_X1    g536(.A(G99gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n728), .A2(new_n738), .A3(new_n643), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n730), .A2(new_n333), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n740), .A2(KEYINPUT111), .ZN(new_n741));
  OAI21_X1  g540(.A(G99gat), .B1(new_n740), .B2(KEYINPUT111), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(G1338gat));
  NOR2_X1   g542(.A1(new_n385), .A2(G106gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(KEYINPUT113), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(KEYINPUT53), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n386), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G106gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n745), .A2(KEYINPUT113), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n745), .A2(KEYINPUT112), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n728), .A2(new_n753), .A3(new_n744), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n749), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT53), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n751), .A2(new_n756), .ZN(G1339gat));
  NOR2_X1   g556(.A1(new_n630), .A2(new_n547), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n534), .A2(new_n535), .A3(new_n533), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n526), .B1(new_n525), .B2(new_n528), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n542), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n761), .A2(KEYINPUT116), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(KEYINPUT116), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n762), .A2(new_n546), .A3(new_n628), .A4(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n610), .B1(new_n618), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n618), .A2(new_n765), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n616), .A2(new_n613), .A3(new_n617), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n767), .A2(KEYINPUT114), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT114), .B1(new_n767), .B2(new_n768), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n766), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n547), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT115), .B1(new_n772), .B2(new_n773), .ZN(new_n776));
  INV_X1    g575(.A(new_n766), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n767), .A2(new_n768), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n777), .B1(new_n780), .B2(new_n769), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n782), .A3(KEYINPUT55), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n626), .A2(new_n627), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n776), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n764), .B1(new_n775), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n606), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n605), .A2(new_n774), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n762), .A2(new_n546), .A3(new_n763), .ZN(new_n790));
  OR3_X1    g589(.A1(new_n789), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n758), .B1(new_n792), .B2(new_n668), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n386), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n794), .A2(new_n452), .A3(new_n482), .A4(new_n643), .ZN(new_n795));
  OAI21_X1  g594(.A(G113gat), .B1(new_n795), .B2(new_n548), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n486), .A2(new_n488), .ZN(new_n797));
  NOR4_X1   g596(.A1(new_n793), .A2(new_n653), .A3(new_n414), .A4(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n238), .A3(new_n547), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(new_n799), .ZN(G1340gat));
  NOR3_X1   g599(.A1(new_n795), .A2(new_n239), .A3(new_n629), .ZN(new_n801));
  AOI21_X1  g600(.A(G120gat), .B1(new_n798), .B2(new_n628), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(G1341gat));
  NOR3_X1   g602(.A1(new_n795), .A2(new_n248), .A3(new_n668), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n798), .A2(new_n576), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n805), .A2(KEYINPUT117), .ZN(new_n806));
  AOI21_X1  g605(.A(G127gat), .B1(new_n805), .B2(KEYINPUT117), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(G1342gat));
  NAND3_X1  g607(.A1(new_n798), .A2(new_n246), .A3(new_n605), .ZN(new_n809));
  XNOR2_X1  g608(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  OAI21_X1  g611(.A(G134gat), .B1(new_n795), .B2(new_n606), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(G1343gat));
  NAND2_X1  g613(.A1(new_n452), .A2(new_n482), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n333), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n385), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n789), .A2(new_n786), .A3(new_n790), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n788), .B2(new_n821), .ZN(new_n822));
  AOI211_X1 g621(.A(new_n773), .B(new_n777), .C1(new_n780), .C2(new_n769), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n784), .B1(new_n823), .B2(new_n782), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n824), .A2(new_n547), .A3(new_n776), .A4(new_n774), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n605), .B1(new_n825), .B2(new_n764), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT119), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n576), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n819), .B1(new_n828), .B2(new_n758), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n818), .B1(new_n793), .B2(new_n385), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n817), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n353), .B1(new_n831), .B2(new_n547), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n793), .A2(new_n653), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n333), .A2(new_n385), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n482), .B1(new_n835), .B2(KEYINPUT120), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(KEYINPUT120), .B2(new_n835), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(G141gat), .A3(new_n548), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT58), .B1(new_n832), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n819), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n791), .B1(new_n826), .B2(KEYINPUT119), .ZN(new_n842));
  AOI211_X1 g641(.A(new_n821), .B(new_n605), .C1(new_n825), .C2(new_n764), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n668), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n631), .A2(new_n548), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n841), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n668), .B1(new_n826), .B2(new_n820), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n845), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(new_n848), .B2(new_n386), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n547), .B(new_n816), .C1(new_n846), .C2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n829), .A2(new_n830), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n853), .A2(KEYINPUT121), .A3(new_n547), .A4(new_n816), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n852), .A2(new_n854), .A3(G141gat), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n839), .A2(KEYINPUT58), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n840), .B1(new_n855), .B2(new_n856), .ZN(G1344gat));
  INV_X1    g656(.A(new_n838), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n355), .A3(new_n628), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n793), .A2(new_n818), .A3(new_n385), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(new_n849), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n628), .A3(new_n816), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n860), .B1(new_n863), .B2(G148gat), .ZN(new_n864));
  AOI211_X1 g663(.A(KEYINPUT59), .B(new_n355), .C1(new_n831), .C2(new_n628), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n859), .B1(new_n864), .B2(new_n865), .ZN(G1345gat));
  NAND3_X1  g665(.A1(new_n858), .A2(new_n359), .A3(new_n576), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n831), .A2(new_n576), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n868), .B2(new_n359), .ZN(G1346gat));
  AOI21_X1  g668(.A(G162gat), .B1(new_n858), .B2(new_n605), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n606), .A2(new_n360), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n831), .B2(new_n871), .ZN(G1347gat));
  NAND3_X1  g671(.A1(new_n643), .A2(new_n653), .A3(new_n414), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT123), .Z(new_n874));
  NAND2_X1  g673(.A1(new_n794), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n219), .A3(new_n548), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n793), .B2(new_n452), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n848), .A2(KEYINPUT122), .A3(new_n653), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n797), .A2(new_n482), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n547), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n876), .B1(new_n883), .B2(new_n219), .ZN(G1348gat));
  NOR3_X1   g683(.A1(new_n875), .A2(new_n277), .A3(new_n629), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n882), .A2(new_n628), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n220), .ZN(G1349gat));
  NAND4_X1  g686(.A1(new_n880), .A2(new_n213), .A3(new_n576), .A4(new_n881), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n794), .A2(new_n576), .A3(new_n874), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(G183gat), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n892), .B(new_n893), .ZN(G1350gat));
  NAND3_X1  g693(.A1(new_n882), .A2(new_n209), .A3(new_n605), .ZN(new_n895));
  OAI21_X1  g694(.A(G190gat), .B1(new_n875), .B2(new_n606), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n896), .A2(KEYINPUT61), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(KEYINPUT61), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(G1351gat));
  NOR3_X1   g698(.A1(new_n333), .A2(new_n452), .A3(new_n482), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n862), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G197gat), .B1(new_n901), .B2(new_n548), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n835), .A2(new_n482), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n904), .B1(new_n878), .B2(new_n879), .ZN(new_n905));
  INV_X1    g704(.A(G197gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n906), .A3(new_n547), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n902), .B1(new_n909), .B2(new_n910), .ZN(G1352gat));
  NOR2_X1   g710(.A1(new_n629), .A2(G204gat), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n793), .A2(new_n877), .A3(new_n452), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT122), .B1(new_n848), .B2(new_n653), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n903), .B(new_n912), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT127), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n905), .A2(new_n917), .A3(new_n912), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(G204gat), .B1(new_n901), .B2(new_n629), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n916), .A2(new_n918), .A3(KEYINPUT62), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G1353gat));
  NAND3_X1  g723(.A1(new_n905), .A2(new_n339), .A3(new_n576), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n576), .B(new_n900), .C1(new_n861), .C2(new_n849), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n926), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT63), .B1(new_n926), .B2(G211gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(G1354gat));
  OAI21_X1  g728(.A(G218gat), .B1(new_n901), .B2(new_n606), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n905), .A2(new_n340), .A3(new_n605), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1355gat));
endmodule


