

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U323 ( .A(n435), .B(n434), .ZN(n439) );
  XNOR2_X1 U324 ( .A(n405), .B(n291), .ZN(n362) );
  XNOR2_X1 U325 ( .A(n412), .B(n411), .ZN(n497) );
  AND2_X1 U326 ( .A1(G227GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U327 ( .A(KEYINPUT45), .B(KEYINPUT111), .ZN(n457) );
  XNOR2_X1 U328 ( .A(n458), .B(n457), .ZN(n459) );
  INV_X1 U329 ( .A(KEYINPUT112), .ZN(n463) );
  XNOR2_X1 U330 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U331 ( .A(n463), .B(KEYINPUT48), .ZN(n464) );
  XNOR2_X1 U332 ( .A(n362), .B(n435), .ZN(n366) );
  XNOR2_X1 U333 ( .A(n465), .B(n464), .ZN(n528) );
  XNOR2_X1 U334 ( .A(KEYINPUT37), .B(KEYINPUT99), .ZN(n411) );
  XOR2_X1 U335 ( .A(n445), .B(n444), .Z(n484) );
  NOR2_X1 U336 ( .A1(n376), .A2(n474), .ZN(n562) );
  XOR2_X1 U337 ( .A(n429), .B(n428), .Z(n567) );
  XNOR2_X1 U338 ( .A(KEYINPUT28), .B(n472), .ZN(n535) );
  XNOR2_X1 U339 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n475) );
  XNOR2_X1 U340 ( .A(n447), .B(G106GAT), .ZN(n448) );
  XNOR2_X1 U341 ( .A(n476), .B(n475), .ZN(G1351GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT12), .B(KEYINPUT74), .Z(n293) );
  XNOR2_X1 U343 ( .A(KEYINPUT14), .B(KEYINPUT73), .ZN(n292) );
  XNOR2_X1 U344 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U345 ( .A(G22GAT), .B(G155GAT), .Z(n346) );
  XOR2_X1 U346 ( .A(n346), .B(G71GAT), .Z(n295) );
  XOR2_X1 U347 ( .A(G15GAT), .B(G127GAT), .Z(n368) );
  XNOR2_X1 U348 ( .A(G1GAT), .B(n368), .ZN(n294) );
  XNOR2_X1 U349 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U350 ( .A(n297), .B(n296), .Z(n299) );
  NAND2_X1 U351 ( .A1(G231GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U353 ( .A(KEYINPUT15), .B(G64GAT), .Z(n301) );
  XNOR2_X1 U354 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U356 ( .A(n303), .B(n302), .Z(n307) );
  XNOR2_X1 U357 ( .A(G78GAT), .B(G57GAT), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n304), .B(KEYINPUT13), .ZN(n441) );
  XNOR2_X1 U359 ( .A(G8GAT), .B(G183GAT), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n305), .B(G211GAT), .ZN(n340) );
  XNOR2_X1 U361 ( .A(n441), .B(n340), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n307), .B(n306), .ZN(n578) );
  XOR2_X1 U363 ( .A(G113GAT), .B(KEYINPUT0), .Z(n367) );
  XOR2_X1 U364 ( .A(G85GAT), .B(G162GAT), .Z(n309) );
  XNOR2_X1 U365 ( .A(G29GAT), .B(G134GAT), .ZN(n308) );
  XNOR2_X1 U366 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U367 ( .A(n367), .B(n310), .Z(n312) );
  NAND2_X1 U368 ( .A1(G225GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U370 ( .A(n313), .B(KEYINPUT6), .Z(n317) );
  XOR2_X1 U371 ( .A(KEYINPUT83), .B(KEYINPUT3), .Z(n315) );
  XNOR2_X1 U372 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n314) );
  XNOR2_X1 U373 ( .A(n315), .B(n314), .ZN(n352) );
  XNOR2_X1 U374 ( .A(n352), .B(KEYINPUT1), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U376 ( .A(G148GAT), .B(G155GAT), .Z(n319) );
  XNOR2_X1 U377 ( .A(G127GAT), .B(G120GAT), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U379 ( .A(n321), .B(n320), .Z(n329) );
  XOR2_X1 U380 ( .A(KEYINPUT85), .B(G57GAT), .Z(n323) );
  XNOR2_X1 U381 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U383 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n325) );
  XNOR2_X1 U384 ( .A(KEYINPUT88), .B(KEYINPUT4), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n529) );
  XOR2_X1 U388 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n331) );
  XNOR2_X1 U389 ( .A(KEYINPUT18), .B(G176GAT), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U391 ( .A(G169GAT), .B(n332), .Z(n371) );
  INV_X1 U392 ( .A(n371), .ZN(n344) );
  XOR2_X1 U393 ( .A(G36GAT), .B(G190GAT), .Z(n397) );
  XOR2_X1 U394 ( .A(KEYINPUT89), .B(n397), .Z(n334) );
  NAND2_X1 U395 ( .A1(G226GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U396 ( .A(n334), .B(n333), .ZN(n336) );
  XNOR2_X1 U397 ( .A(G204GAT), .B(G92GAT), .ZN(n335) );
  XNOR2_X1 U398 ( .A(n335), .B(G64GAT), .ZN(n440) );
  XOR2_X1 U399 ( .A(n336), .B(n440), .Z(n342) );
  XOR2_X1 U400 ( .A(KEYINPUT21), .B(G218GAT), .Z(n338) );
  XNOR2_X1 U401 ( .A(KEYINPUT82), .B(KEYINPUT81), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U403 ( .A(G197GAT), .B(n339), .Z(n360) );
  XNOR2_X1 U404 ( .A(n360), .B(n340), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U406 ( .A(n344), .B(n343), .Z(n377) );
  INV_X1 U407 ( .A(n377), .ZN(n522) );
  XOR2_X1 U408 ( .A(KEYINPUT27), .B(KEYINPUT90), .Z(n345) );
  XOR2_X1 U409 ( .A(n522), .B(n345), .Z(n385) );
  INV_X1 U410 ( .A(n385), .ZN(n530) );
  XOR2_X1 U411 ( .A(KEYINPUT84), .B(G78GAT), .Z(n348) );
  XOR2_X1 U412 ( .A(G106GAT), .B(G148GAT), .Z(n431) );
  XNOR2_X1 U413 ( .A(n346), .B(n431), .ZN(n347) );
  XNOR2_X1 U414 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U415 ( .A(G50GAT), .B(G162GAT), .Z(n393) );
  XOR2_X1 U416 ( .A(n349), .B(n393), .Z(n358) );
  XOR2_X1 U417 ( .A(G211GAT), .B(KEYINPUT23), .Z(n351) );
  XNOR2_X1 U418 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n350) );
  XNOR2_X1 U419 ( .A(n351), .B(n350), .ZN(n356) );
  XOR2_X1 U420 ( .A(n352), .B(G204GAT), .Z(n354) );
  NAND2_X1 U421 ( .A1(G228GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U423 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U424 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U425 ( .A(n360), .B(n359), .ZN(n472) );
  XOR2_X1 U426 ( .A(G43GAT), .B(G134GAT), .Z(n405) );
  XNOR2_X1 U427 ( .A(G99GAT), .B(G71GAT), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n361), .B(G120GAT), .ZN(n435) );
  XOR2_X1 U429 ( .A(G183GAT), .B(KEYINPUT79), .Z(n364) );
  XNOR2_X1 U430 ( .A(G190GAT), .B(KEYINPUT20), .ZN(n363) );
  XNOR2_X1 U431 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U432 ( .A(n366), .B(n365), .Z(n370) );
  XNOR2_X1 U433 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U434 ( .A(n370), .B(n369), .ZN(n372) );
  XOR2_X1 U435 ( .A(n372), .B(n371), .Z(n376) );
  NAND2_X1 U436 ( .A1(n472), .A2(n376), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n373), .B(KEYINPUT26), .ZN(n564) );
  NOR2_X1 U438 ( .A1(n530), .A2(n564), .ZN(n374) );
  XOR2_X1 U439 ( .A(KEYINPUT91), .B(n374), .Z(n375) );
  NOR2_X1 U440 ( .A1(n529), .A2(n375), .ZN(n382) );
  NOR2_X1 U441 ( .A1(n376), .A2(n377), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n378), .B(KEYINPUT92), .ZN(n379) );
  NOR2_X1 U443 ( .A1(n472), .A2(n379), .ZN(n380) );
  XNOR2_X1 U444 ( .A(KEYINPUT25), .B(n380), .ZN(n381) );
  NAND2_X1 U445 ( .A1(n382), .A2(n381), .ZN(n388) );
  INV_X1 U446 ( .A(n376), .ZN(n526) );
  XNOR2_X1 U447 ( .A(n526), .B(KEYINPUT80), .ZN(n383) );
  NOR2_X1 U448 ( .A1(n535), .A2(n383), .ZN(n384) );
  NAND2_X1 U449 ( .A1(n385), .A2(n384), .ZN(n386) );
  NAND2_X1 U450 ( .A1(n386), .A2(n529), .ZN(n387) );
  NAND2_X1 U451 ( .A1(n388), .A2(n387), .ZN(n389) );
  XOR2_X1 U452 ( .A(KEYINPUT93), .B(n389), .Z(n482) );
  NOR2_X1 U453 ( .A1(n578), .A2(n482), .ZN(n390) );
  XNOR2_X1 U454 ( .A(KEYINPUT98), .B(n390), .ZN(n410) );
  XOR2_X1 U455 ( .A(KEYINPUT70), .B(KEYINPUT10), .Z(n392) );
  XNOR2_X1 U456 ( .A(G99GAT), .B(KEYINPUT9), .ZN(n391) );
  XNOR2_X1 U457 ( .A(n392), .B(n391), .ZN(n409) );
  XOR2_X1 U458 ( .A(G85GAT), .B(KEYINPUT68), .Z(n430) );
  XOR2_X1 U459 ( .A(G92GAT), .B(n430), .Z(n395) );
  XNOR2_X1 U460 ( .A(G218GAT), .B(n393), .ZN(n394) );
  XNOR2_X1 U461 ( .A(n395), .B(n394), .ZN(n401) );
  XNOR2_X1 U462 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n396), .B(KEYINPUT8), .ZN(n421) );
  XNOR2_X1 U464 ( .A(n421), .B(n397), .ZN(n399) );
  AND2_X1 U465 ( .A1(G232GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U466 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U467 ( .A(n401), .B(n400), .Z(n407) );
  XOR2_X1 U468 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n403) );
  XNOR2_X1 U469 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U471 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n409), .B(n408), .ZN(n553) );
  INV_X1 U474 ( .A(n553), .ZN(n477) );
  XOR2_X1 U475 ( .A(KEYINPUT36), .B(n477), .Z(n582) );
  NAND2_X1 U476 ( .A1(n410), .A2(n582), .ZN(n412) );
  XOR2_X1 U477 ( .A(G15GAT), .B(G197GAT), .Z(n414) );
  XNOR2_X1 U478 ( .A(G169GAT), .B(G141GAT), .ZN(n413) );
  XNOR2_X1 U479 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U480 ( .A(KEYINPUT29), .B(G8GAT), .Z(n416) );
  XNOR2_X1 U481 ( .A(G113GAT), .B(G1GAT), .ZN(n415) );
  XNOR2_X1 U482 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U483 ( .A(n418), .B(n417), .ZN(n429) );
  XOR2_X1 U484 ( .A(G43GAT), .B(G36GAT), .Z(n420) );
  XNOR2_X1 U485 ( .A(G50GAT), .B(G22GAT), .ZN(n419) );
  XNOR2_X1 U486 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U487 ( .A(n422), .B(n421), .Z(n427) );
  XOR2_X1 U488 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n424) );
  NAND2_X1 U489 ( .A1(G229GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U490 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U491 ( .A(KEYINPUT30), .B(n425), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n427), .B(n426), .ZN(n428) );
  INV_X1 U493 ( .A(n567), .ZN(n485) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n445) );
  NAND2_X1 U495 ( .A1(G230GAT), .A2(G233GAT), .ZN(n433) );
  INV_X1 U496 ( .A(KEYINPUT67), .ZN(n432) );
  XOR2_X1 U497 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n437) );
  XNOR2_X1 U498 ( .A(G176GAT), .B(KEYINPUT32), .ZN(n436) );
  XOR2_X1 U499 ( .A(n437), .B(n436), .Z(n438) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U503 ( .A(n484), .B(KEYINPUT41), .ZN(n450) );
  NAND2_X1 U504 ( .A1(n485), .A2(n450), .ZN(n512) );
  NOR2_X1 U505 ( .A1(n497), .A2(n512), .ZN(n446) );
  XOR2_X1 U506 ( .A(KEYINPUT105), .B(n446), .Z(n525) );
  NAND2_X1 U507 ( .A1(n525), .A2(n535), .ZN(n449) );
  XOR2_X1 U508 ( .A(KEYINPUT107), .B(KEYINPUT44), .Z(n447) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(G1339GAT) );
  XOR2_X1 U510 ( .A(n522), .B(KEYINPUT117), .Z(n466) );
  XNOR2_X1 U511 ( .A(n578), .B(KEYINPUT108), .ZN(n561) );
  AND2_X1 U512 ( .A1(n567), .A2(n450), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n451), .B(KEYINPUT46), .ZN(n452) );
  NOR2_X1 U514 ( .A1(n561), .A2(n452), .ZN(n453) );
  NAND2_X1 U515 ( .A1(n453), .A2(n477), .ZN(n455) );
  XOR2_X1 U516 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n454) );
  XNOR2_X1 U517 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U518 ( .A(n456), .B(KEYINPUT47), .ZN(n462) );
  NAND2_X1 U519 ( .A1(n578), .A2(n582), .ZN(n458) );
  NAND2_X1 U520 ( .A1(n459), .A2(n484), .ZN(n460) );
  NOR2_X1 U521 ( .A1(n567), .A2(n460), .ZN(n461) );
  NOR2_X1 U522 ( .A1(n462), .A2(n461), .ZN(n465) );
  NAND2_X1 U523 ( .A1(n466), .A2(n528), .ZN(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT54), .B(KEYINPUT118), .Z(n467) );
  XNOR2_X1 U525 ( .A(KEYINPUT119), .B(n467), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n469), .B(n468), .ZN(n470) );
  NOR2_X1 U527 ( .A1(n470), .A2(n529), .ZN(n471) );
  XOR2_X1 U528 ( .A(KEYINPUT64), .B(n471), .Z(n565) );
  NOR2_X1 U529 ( .A1(n565), .A2(n472), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n473), .B(KEYINPUT55), .ZN(n474) );
  NAND2_X1 U531 ( .A1(n553), .A2(n562), .ZN(n476) );
  XOR2_X1 U532 ( .A(KEYINPUT16), .B(KEYINPUT78), .Z(n479) );
  NAND2_X1 U533 ( .A1(n578), .A2(n477), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U535 ( .A(n480), .B(KEYINPUT77), .ZN(n481) );
  NOR2_X1 U536 ( .A1(n482), .A2(n481), .ZN(n483) );
  XOR2_X1 U537 ( .A(KEYINPUT94), .B(n483), .Z(n513) );
  INV_X1 U538 ( .A(n484), .ZN(n574) );
  NOR2_X1 U539 ( .A1(n574), .A2(n485), .ZN(n486) );
  XNOR2_X1 U540 ( .A(n486), .B(KEYINPUT69), .ZN(n498) );
  NOR2_X1 U541 ( .A1(n513), .A2(n498), .ZN(n495) );
  NAND2_X1 U542 ( .A1(n495), .A2(n529), .ZN(n490) );
  XOR2_X1 U543 ( .A(KEYINPUT34), .B(KEYINPUT95), .Z(n488) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(KEYINPUT96), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U546 ( .A(n490), .B(n489), .ZN(G1324GAT) );
  XOR2_X1 U547 ( .A(G8GAT), .B(KEYINPUT97), .Z(n492) );
  NAND2_X1 U548 ( .A1(n495), .A2(n522), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n492), .B(n491), .ZN(G1325GAT) );
  XOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT35), .Z(n494) );
  NAND2_X1 U551 ( .A1(n495), .A2(n526), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U553 ( .A1(n495), .A2(n535), .ZN(n496) );
  XNOR2_X1 U554 ( .A(n496), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT39), .Z(n502) );
  NOR2_X1 U556 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U557 ( .A(n499), .B(KEYINPUT38), .ZN(n500) );
  XNOR2_X1 U558 ( .A(KEYINPUT100), .B(n500), .ZN(n508) );
  NAND2_X1 U559 ( .A1(n508), .A2(n529), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  XOR2_X1 U561 ( .A(G36GAT), .B(KEYINPUT101), .Z(n504) );
  NAND2_X1 U562 ( .A1(n508), .A2(n522), .ZN(n503) );
  XNOR2_X1 U563 ( .A(n504), .B(n503), .ZN(G1329GAT) );
  NAND2_X1 U564 ( .A1(n526), .A2(n508), .ZN(n507) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n505), .B(KEYINPUT102), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n507), .B(n506), .ZN(G1330GAT) );
  NAND2_X1 U568 ( .A1(n508), .A2(n535), .ZN(n509) );
  XNOR2_X1 U569 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n510), .B(KEYINPUT103), .ZN(n511) );
  XOR2_X1 U572 ( .A(KEYINPUT104), .B(n511), .Z(n515) );
  NOR2_X1 U573 ( .A1(n513), .A2(n512), .ZN(n518) );
  NAND2_X1 U574 ( .A1(n518), .A2(n529), .ZN(n514) );
  XNOR2_X1 U575 ( .A(n515), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U576 ( .A1(n518), .A2(n522), .ZN(n516) );
  XNOR2_X1 U577 ( .A(n516), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n526), .A2(n518), .ZN(n517) );
  XNOR2_X1 U579 ( .A(n517), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U581 ( .A1(n518), .A2(n535), .ZN(n519) );
  XNOR2_X1 U582 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NAND2_X1 U583 ( .A1(n529), .A2(n525), .ZN(n521) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n525), .A2(n522), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n523), .B(KEYINPUT106), .ZN(n524) );
  XNOR2_X1 U587 ( .A(G92GAT), .B(n524), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U589 ( .A(n527), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n531) );
  NOR2_X1 U591 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U592 ( .A(n532), .B(KEYINPUT113), .ZN(n545) );
  NOR2_X1 U593 ( .A1(n376), .A2(n545), .ZN(n533) );
  XOR2_X1 U594 ( .A(KEYINPUT114), .B(n533), .Z(n534) );
  NOR2_X1 U595 ( .A1(n535), .A2(n534), .ZN(n542) );
  NAND2_X1 U596 ( .A1(n567), .A2(n542), .ZN(n536) );
  XNOR2_X1 U597 ( .A(n536), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U599 ( .A1(n542), .A2(n450), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n540) );
  NAND2_X1 U602 ( .A1(n542), .A2(n561), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U606 ( .A1(n542), .A2(n553), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NOR2_X1 U608 ( .A1(n564), .A2(n545), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n552), .A2(n567), .ZN(n546) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  NAND2_X1 U612 ( .A1(n552), .A2(n450), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n552), .A2(n578), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(KEYINPUT116), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(n551), .ZN(G1346GAT) );
  NAND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n562), .A2(n567), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(n555), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n557) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(KEYINPUT120), .B(n558), .Z(n560) );
  NAND2_X1 U626 ( .A1(n562), .A2(n450), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n569) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n566), .A2(n567), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n569), .B(n568), .ZN(n571) );
  INV_X1 U634 ( .A(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(n573) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n576) );
  NAND2_X1 U639 ( .A1(n566), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(n577), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n580) );
  NAND2_X1 U643 ( .A1(n566), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U647 ( .A1(n566), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

