//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT24), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n203), .A2(G183gat), .A3(G190gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(G183gat), .B(G190gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(new_n203), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT65), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n208), .B(new_n204), .C1(new_n205), .C2(new_n203), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT23), .ZN(new_n212));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT64), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(KEYINPUT64), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217));
  INV_X1    g016(.A(new_n211), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n210), .A2(new_n215), .A3(new_n216), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n214), .B1(KEYINPUT23), .B2(new_n211), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n217), .B1(new_n222), .B2(new_n206), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT27), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT27), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G183gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT28), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n229), .A2(new_n230), .A3(G190gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(G190gat), .B1(new_n226), .B2(KEYINPUT66), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n231), .B1(new_n235), .B2(new_n230), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT26), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n237), .A3(new_n213), .ZN(new_n238));
  INV_X1    g037(.A(G190gat), .ZN(new_n239));
  OAI221_X1 g038(.A(new_n238), .B1(new_n237), .B2(new_n218), .C1(new_n225), .C2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT67), .B1(new_n236), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n236), .A2(KEYINPUT67), .A3(new_n240), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n224), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G134gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(KEYINPUT68), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n246), .B1(new_n247), .B2(KEYINPUT1), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n249));
  INV_X1    g048(.A(G113gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(G120gat), .ZN(new_n251));
  INV_X1    g050(.A(G120gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n252), .A2(G113gat), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n249), .B(new_n245), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G127gat), .ZN(new_n256));
  INV_X1    g055(.A(G127gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n248), .A2(new_n257), .A3(new_n254), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n256), .A2(KEYINPUT69), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT69), .B1(new_n256), .B2(new_n258), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n256), .A2(KEYINPUT69), .A3(new_n258), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n224), .B(new_n263), .C1(new_n242), .C2(new_n243), .ZN(new_n264));
  AOI211_X1 g063(.A(KEYINPUT70), .B(new_n202), .C1(new_n262), .C2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n235), .A2(new_n230), .ZN(new_n267));
  INV_X1    g066(.A(new_n231), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n240), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n271), .A2(new_n241), .B1(new_n223), .B2(new_n221), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n259), .A2(new_n260), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n264), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n202), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n266), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT32), .B1(new_n265), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT33), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n265), .B2(new_n276), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT34), .B1(new_n274), .B2(new_n275), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT34), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n262), .A2(new_n281), .A3(new_n202), .A4(new_n264), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(G15gat), .B(G43gat), .Z(new_n284));
  XNOR2_X1  g083(.A(G71gat), .B(G99gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n279), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n283), .B1(new_n279), .B2(new_n286), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n277), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n283), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT70), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n266), .A3(new_n275), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT33), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n286), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n290), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n277), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n283), .A3(new_n286), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT79), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n301));
  INV_X1    g100(.A(G141gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(G148gat), .ZN(new_n303));
  INV_X1    g102(.A(G148gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(G141gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n301), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G155gat), .ZN(new_n307));
  INV_X1    g106(.A(G162gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT78), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(new_n302), .B2(G148gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n304), .A2(KEYINPUT78), .A3(G141gat), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n314), .B(new_n315), .C1(G141gat), .C2(new_n304), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n310), .B1(new_n309), .B2(KEYINPUT2), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n300), .B1(new_n319), .B2(KEYINPUT3), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n306), .A2(new_n311), .B1(new_n316), .B2(new_n317), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(KEYINPUT79), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT22), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n327), .A2(KEYINPUT71), .B1(G211gat), .B2(G218gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(KEYINPUT71), .B2(new_n327), .ZN(new_n329));
  XNOR2_X1  g128(.A(G197gat), .B(G204gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(G211gat), .B(G218gat), .Z(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT72), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n331), .B(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n326), .A2(new_n334), .ZN(new_n335));
  AND2_X1   g134(.A1(G228gat), .A2(G233gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n334), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT3), .B1(new_n337), .B2(new_n325), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n335), .B(new_n336), .C1(new_n321), .C2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n332), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT29), .B1(new_n331), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(new_n340), .B2(new_n331), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n321), .B1(new_n342), .B2(new_n322), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n326), .B2(new_n334), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n339), .B1(new_n336), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G78gat), .B(G106gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT31), .B(G50gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G22gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(KEYINPUT84), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n350), .B1(new_n349), .B2(new_n348), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n345), .B(new_n351), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n289), .A2(new_n299), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT35), .ZN(new_n354));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT0), .ZN(new_n356));
  XNOR2_X1  g155(.A(G57gat), .B(G85gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n257), .B1(new_n248), .B2(new_n254), .ZN(new_n360));
  INV_X1    g159(.A(new_n258), .ZN(new_n361));
  AOI211_X1 g160(.A(new_n360), .B(new_n361), .C1(KEYINPUT3), .C2(new_n319), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n321), .B1(new_n361), .B2(new_n360), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT4), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n365), .B(new_n321), .C1(new_n361), .C2(new_n360), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n362), .A2(new_n324), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n368), .B(KEYINPUT80), .Z(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n256), .A2(new_n319), .A3(new_n258), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n363), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n369), .ZN(new_n376));
  INV_X1    g175(.A(new_n371), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(KEYINPUT83), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT83), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n370), .B1(new_n363), .B2(new_n374), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n379), .B1(new_n380), .B2(new_n371), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n369), .B1(new_n362), .B2(new_n324), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n319), .B1(new_n256), .B2(new_n258), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(KEYINPUT81), .A3(new_n365), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n366), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n386), .A3(new_n364), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n378), .A2(new_n381), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n359), .B1(new_n373), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n378), .A2(new_n381), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n382), .A2(new_n387), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n392), .A2(new_n372), .A3(new_n358), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT6), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n389), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  OAI211_X1 g194(.A(KEYINPUT6), .B(new_n359), .C1(new_n373), .C2(new_n388), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n398), .B(KEYINPUT73), .Z(new_n399));
  NAND2_X1  g198(.A1(new_n244), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n399), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n269), .B1(new_n221), .B2(new_n223), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(KEYINPUT29), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n400), .A2(new_n337), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n399), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n401), .A2(new_n325), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n405), .B(new_n334), .C1(new_n272), .C2(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(G8gat), .B(G36gat), .Z(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(KEYINPUT74), .ZN(new_n409));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n404), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT76), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n413), .B1(new_n412), .B2(new_n414), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT75), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n407), .ZN(new_n420));
  INV_X1    g219(.A(new_n411), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI211_X1 g221(.A(KEYINPUT75), .B(new_n411), .C1(new_n404), .C2(new_n407), .ZN(new_n423));
  OAI22_X1  g222(.A1(new_n422), .A2(new_n423), .B1(new_n414), .B2(new_n412), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n353), .A2(new_n354), .A3(new_n397), .A4(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n289), .A2(new_n425), .A3(new_n299), .A4(new_n352), .ZN(new_n427));
  INV_X1    g226(.A(new_n397), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT35), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OR3_X1    g228(.A1(new_n367), .A2(KEYINPUT39), .A3(new_n370), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n363), .A2(new_n374), .A3(new_n370), .ZN(new_n431));
  OAI211_X1 g230(.A(KEYINPUT39), .B(new_n431), .C1(new_n367), .C2(new_n370), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n358), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT40), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n430), .A2(new_n432), .A3(KEYINPUT40), .A4(new_n358), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n389), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n412), .A2(new_n414), .ZN(new_n438));
  INV_X1    g237(.A(new_n422), .ZN(new_n439));
  INV_X1    g238(.A(new_n423), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n417), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n415), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n437), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT37), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n404), .A2(new_n445), .A3(new_n407), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n446), .A2(new_n421), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT38), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(new_n420), .B2(KEYINPUT37), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n400), .A2(new_n334), .A3(new_n403), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n405), .B(new_n337), .C1(new_n272), .C2(new_n406), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(KEYINPUT37), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n446), .A2(new_n452), .A3(new_n421), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n447), .A2(new_n449), .B1(new_n453), .B2(new_n448), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n395), .A2(new_n396), .A3(new_n412), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n352), .B1(new_n444), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n352), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n425), .A2(new_n397), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT36), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n287), .A2(new_n288), .A3(new_n277), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n297), .B1(new_n296), .B2(new_n298), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n289), .A2(KEYINPUT36), .A3(new_n299), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n426), .A2(new_n429), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(G71gat), .A2(G78gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(G71gat), .ZN(new_n470));
  INV_X1    g269(.A(G78gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT9), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G64gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(G57gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(G57gat), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(KEYINPUT96), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT96), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n478), .A2(new_n474), .A3(G57gat), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n473), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G57gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(G64gat), .ZN(new_n482));
  OAI22_X1  g281(.A1(new_n476), .A2(new_n482), .B1(KEYINPUT9), .B2(new_n468), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT94), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT94), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(G71gat), .B2(G78gat), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n468), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n483), .B1(new_n487), .B2(KEYINPUT95), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT95), .ZN(new_n489));
  AOI211_X1 g288(.A(new_n489), .B(new_n468), .C1(new_n484), .C2(new_n486), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n480), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  XOR2_X1   g290(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(G231gat), .A2(G233gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(G127gat), .ZN(new_n496));
  INV_X1    g295(.A(G1gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT16), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n349), .A2(G15gat), .ZN(new_n499));
  INV_X1    g298(.A(G15gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(G22gat), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT90), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT90), .B1(new_n499), .B2(new_n501), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n501), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT90), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n497), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT91), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n512), .A3(G8gat), .ZN(new_n513));
  INV_X1    g312(.A(G8gat), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n504), .B(new_n509), .C1(new_n511), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT21), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(new_n491), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n496), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(new_n307), .ZN(new_n522));
  XOR2_X1   g321(.A(G183gat), .B(G211gat), .Z(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n520), .B(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(G232gat), .A2(G233gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(KEYINPUT41), .ZN(new_n527));
  XNOR2_X1  g326(.A(G134gat), .B(G162gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G85gat), .A2(G92gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g330(.A1(G99gat), .A2(G106gat), .ZN(new_n532));
  INV_X1    g331(.A(G85gat), .ZN(new_n533));
  INV_X1    g332(.A(G92gat), .ZN(new_n534));
  AOI22_X1  g333(.A1(KEYINPUT8), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G99gat), .B(G106gat), .Z(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n537), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(new_n531), .A3(new_n535), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT98), .ZN(new_n542));
  XNOR2_X1  g341(.A(G43gat), .B(G50gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT15), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G29gat), .A2(G36gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT14), .ZN(new_n547));
  INV_X1    g346(.A(G29gat), .ZN(new_n548));
  INV_X1    g347(.A(G36gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT87), .ZN(new_n551));
  NOR3_X1   g350(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT87), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT86), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g356(.A(KEYINPUT86), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n551), .A2(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n546), .B1(new_n559), .B2(KEYINPUT88), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n551), .A2(new_n554), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n558), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n561), .A2(KEYINPUT88), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n545), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n550), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n543), .A2(KEYINPUT15), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n546), .B(KEYINPUT89), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n544), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n542), .A2(new_n569), .B1(KEYINPUT41), .B2(new_n526), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n552), .A2(new_n553), .ZN(new_n572));
  NOR4_X1   g371(.A1(KEYINPUT87), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n562), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT88), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n574), .A2(new_n575), .B1(G29gat), .B2(G36gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n561), .A2(KEYINPUT88), .A3(new_n562), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n544), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n568), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n571), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT98), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n541), .B(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n564), .A2(KEYINPUT17), .A3(new_n568), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n570), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT99), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n570), .B(new_n590), .C1(new_n583), .C2(new_n585), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n529), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(new_n529), .A3(new_n591), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n525), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G113gat), .B(G141gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(G169gat), .B(G197gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT12), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT93), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n604), .B1(new_n569), .B2(new_n516), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n574), .A2(new_n575), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(new_n577), .A3(new_n546), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n579), .B1(new_n607), .B2(new_n545), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n608), .A2(KEYINPUT93), .A3(new_n515), .A4(new_n513), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n569), .A2(new_n516), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT13), .Z(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n580), .A2(new_n517), .A3(new_n584), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT18), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT92), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n615), .A2(new_n617), .A3(new_n612), .A4(new_n610), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n564), .A2(new_n568), .B1(new_n513), .B2(new_n515), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n516), .B1(new_n569), .B2(new_n571), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n620), .B1(new_n621), .B2(new_n584), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n617), .B1(new_n622), .B2(new_n612), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n603), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n615), .A2(new_n612), .A3(new_n610), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(KEYINPUT92), .A3(new_n616), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n626), .A2(new_n614), .A3(new_n618), .A4(new_n602), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n491), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g430(.A(KEYINPUT100), .B(new_n480), .C1(new_n488), .C2(new_n490), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n541), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n632), .A2(new_n541), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n633), .A2(KEYINPUT10), .A3(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n484), .A2(new_n486), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n489), .B1(new_n636), .B2(new_n468), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n487), .A2(KEYINPUT95), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(new_n638), .A3(new_n483), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(KEYINPUT10), .A3(new_n480), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n582), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n629), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT101), .ZN(new_n644));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n633), .A2(new_n634), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n642), .B(new_n647), .C1(new_n629), .C2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n629), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n632), .A2(new_n541), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT100), .B1(new_n639), .B2(new_n480), .ZN(new_n653));
  INV_X1    g452(.A(new_n632), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n651), .B(new_n652), .C1(new_n655), .C2(new_n541), .ZN(new_n656));
  INV_X1    g455(.A(new_n640), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n542), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n650), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n648), .A2(new_n629), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n646), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n649), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n596), .A2(new_n628), .A3(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n467), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n428), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  NOR3_X1   g466(.A1(new_n467), .A2(new_n425), .A3(new_n664), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  AND3_X1   g468(.A1(new_n668), .A2(KEYINPUT42), .A3(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n670), .A2(KEYINPUT102), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(KEYINPUT102), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT42), .B1(new_n668), .B2(new_n514), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n671), .B1(new_n672), .B2(new_n675), .ZN(G1325gat));
  NOR2_X1   g475(.A1(new_n462), .A2(new_n463), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n665), .A2(new_n500), .A3(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n467), .A2(new_n466), .A3(new_n664), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(new_n500), .ZN(G1326gat));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n458), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  INV_X1    g482(.A(new_n594), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n592), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n467), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n525), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n624), .A2(new_n627), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n687), .A2(new_n688), .A3(new_n662), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n397), .A2(G29gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT103), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n690), .A2(new_n694), .A3(new_n691), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n693), .A2(KEYINPUT45), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT45), .B1(new_n693), .B2(new_n695), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n426), .A2(new_n429), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n460), .A2(new_n466), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(KEYINPUT44), .A3(new_n595), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n467), .B2(new_n685), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n428), .A3(new_n689), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n548), .B1(new_n706), .B2(KEYINPUT104), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(KEYINPUT104), .B2(new_n706), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n698), .A2(new_n708), .ZN(G1328gat));
  INV_X1    g508(.A(new_n425), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711));
  AOI21_X1  g510(.A(G36gat), .B1(new_n711), .B2(KEYINPUT46), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n690), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n711), .A2(KEYINPUT46), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n705), .A2(new_n710), .A3(new_n689), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(new_n549), .B2(new_n716), .ZN(G1329gat));
  INV_X1    g516(.A(new_n466), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n702), .A2(new_n704), .A3(new_n718), .A4(new_n689), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G43gat), .ZN(new_n720));
  INV_X1    g519(.A(G43gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n690), .A2(new_n721), .A3(new_n677), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n720), .A2(new_n722), .A3(KEYINPUT47), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(KEYINPUT107), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n719), .A2(new_n725), .A3(G43gat), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n724), .A2(new_n726), .A3(new_n722), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n728));
  OAI21_X1  g527(.A(new_n723), .B1(new_n727), .B2(new_n728), .ZN(G1330gat));
  NAND3_X1  g528(.A1(new_n705), .A2(new_n458), .A3(new_n689), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G50gat), .ZN(new_n731));
  NAND2_X1  g530(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n352), .A2(G50gat), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n690), .B2(new_n734), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n731), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n732), .B1(new_n731), .B2(new_n735), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(G1331gat));
  AND4_X1   g537(.A1(new_n701), .A2(new_n688), .A3(new_n596), .A4(new_n662), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n428), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n710), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT49), .B(G64gat), .Z(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(G1333gat));
  AOI21_X1  g544(.A(new_n470), .B1(new_n739), .B2(new_n718), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n462), .A2(new_n463), .A3(G71gat), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n739), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n739), .A2(new_n458), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT109), .B(G78gat), .Z(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1335gat));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n701), .A2(new_n753), .A3(new_n595), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT112), .B1(new_n467), .B2(new_n685), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n687), .A2(new_n628), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT51), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n754), .A2(new_n755), .A3(new_n759), .A4(new_n756), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n758), .A2(new_n662), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(new_n533), .A3(new_n428), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n687), .A2(new_n628), .A3(new_n663), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n702), .A2(new_n704), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT110), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n702), .A2(new_n704), .A3(new_n766), .A4(new_n763), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n428), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT111), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G85gat), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n768), .A2(KEYINPUT111), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n762), .B1(new_n770), .B2(new_n771), .ZN(G1336gat));
  NOR2_X1   g571(.A1(new_n425), .A2(G92gat), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n662), .A3(new_n760), .A4(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  OAI21_X1  g574(.A(G92gat), .B1(new_n764), .B2(new_n425), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n765), .A2(new_n710), .A3(new_n767), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n761), .A2(new_n773), .B1(new_n778), .B2(G92gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n779), .B2(new_n775), .ZN(G1337gat));
  NAND2_X1  g579(.A1(new_n761), .A2(new_n677), .ZN(new_n781));
  INV_X1    g580(.A(G99gat), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n765), .A2(new_n767), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n466), .A2(new_n782), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n781), .A2(new_n782), .B1(new_n783), .B2(new_n784), .ZN(G1338gat));
  NOR2_X1   g584(.A1(new_n352), .A2(G106gat), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n758), .A2(new_n662), .A3(new_n760), .A4(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  OAI21_X1  g587(.A(G106gat), .B1(new_n764), .B2(new_n352), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n765), .A2(new_n458), .A3(new_n767), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n761), .A2(new_n786), .B1(new_n791), .B2(G106gat), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n792), .B2(new_n788), .ZN(G1339gat));
  NAND3_X1  g592(.A1(new_n596), .A2(new_n688), .A3(new_n663), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n656), .A2(new_n650), .A3(new_n658), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n642), .A2(KEYINPUT54), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n646), .B1(new_n642), .B2(KEYINPUT54), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n647), .B1(new_n659), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n642), .A2(new_n796), .A3(KEYINPUT54), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n802), .A3(KEYINPUT55), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n799), .A2(new_n649), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n622), .A2(new_n612), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n611), .A2(new_n613), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n601), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n627), .A2(new_n807), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n804), .A2(new_n685), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n662), .A2(new_n627), .A3(new_n807), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n804), .B2(new_n688), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n809), .B1(new_n685), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n794), .B1(new_n812), .B2(new_n687), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n428), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n427), .ZN(new_n815));
  AOI21_X1  g614(.A(G113gat), .B1(new_n815), .B2(new_n628), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n813), .A2(new_n352), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n710), .A2(new_n397), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n817), .A2(new_n677), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n688), .A2(new_n250), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(G1340gat));
  AOI21_X1  g620(.A(G120gat), .B1(new_n815), .B2(new_n662), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n663), .A2(new_n252), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n819), .B2(new_n823), .ZN(G1341gat));
  XNOR2_X1  g623(.A(KEYINPUT68), .B(G127gat), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n525), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n815), .A2(new_n687), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n819), .A2(new_n826), .B1(new_n827), .B2(new_n825), .ZN(G1342gat));
  NAND3_X1  g627(.A1(new_n815), .A2(new_n245), .A3(new_n595), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT56), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT113), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n819), .A2(new_n595), .ZN(new_n832));
  OAI221_X1 g631(.A(new_n831), .B1(KEYINPUT56), .B2(new_n829), .C1(new_n245), .C2(new_n832), .ZN(G1343gat));
  NAND2_X1  g632(.A1(new_n799), .A2(KEYINPUT114), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n835), .B(new_n795), .C1(new_n797), .C2(new_n798), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n628), .A2(new_n649), .A3(new_n803), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n810), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n809), .B1(new_n839), .B2(new_n685), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n794), .B1(new_n840), .B2(new_n687), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT57), .B1(new_n842), .B2(new_n352), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n466), .A2(new_n818), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n813), .A2(new_n458), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n843), .B(new_n844), .C1(KEYINPUT57), .C2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(G141gat), .B1(new_n846), .B2(new_n688), .ZN(new_n847));
  INV_X1    g646(.A(new_n814), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n718), .A2(new_n352), .A3(new_n710), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n628), .A2(new_n302), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n847), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g652(.A(new_n850), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n304), .A3(new_n662), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n846), .A2(new_n663), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n304), .A2(KEYINPUT59), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT115), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT115), .B(new_n857), .C1(new_n846), .C2(new_n663), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n352), .B1(new_n841), .B2(KEYINPUT117), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n864), .B(new_n794), .C1(new_n840), .C2(new_n687), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT57), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n811), .A2(new_n685), .ZN(new_n867));
  INV_X1    g666(.A(new_n809), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n687), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR4_X1   g668(.A1(new_n525), .A2(new_n595), .A3(new_n628), .A4(new_n662), .ZN(new_n870));
  OAI211_X1 g669(.A(KEYINPUT57), .B(new_n458), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n813), .A2(KEYINPUT116), .A3(KEYINPUT57), .A4(new_n458), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n866), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n662), .A3(new_n844), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n862), .B1(new_n878), .B2(G148gat), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n855), .B1(new_n861), .B2(new_n879), .ZN(G1345gat));
  OAI21_X1  g679(.A(G155gat), .B1(new_n846), .B2(new_n525), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n854), .A2(new_n307), .A3(new_n687), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1346gat));
  NOR3_X1   g682(.A1(new_n846), .A2(new_n308), .A3(new_n685), .ZN(new_n884));
  AOI21_X1  g683(.A(G162gat), .B1(new_n854), .B2(new_n595), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(G1347gat));
  AND2_X1   g685(.A1(new_n813), .A2(new_n397), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n887), .A2(new_n710), .A3(new_n353), .ZN(new_n888));
  AOI21_X1  g687(.A(G169gat), .B1(new_n888), .B2(new_n628), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n425), .A2(new_n428), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n677), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n817), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n628), .A2(G169gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(G1348gat));
  INV_X1    g693(.A(new_n892), .ZN(new_n895));
  OAI21_X1  g694(.A(G176gat), .B1(new_n895), .B2(new_n663), .ZN(new_n896));
  INV_X1    g695(.A(G176gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n888), .A2(new_n897), .A3(new_n662), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1349gat));
  AOI21_X1  g698(.A(new_n225), .B1(new_n892), .B2(new_n687), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n525), .A2(new_n229), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n888), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(KEYINPUT60), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT60), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(KEYINPUT119), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n904), .A2(new_n906), .B1(new_n902), .B2(new_n907), .ZN(G1350gat));
  NAND3_X1  g707(.A1(new_n888), .A2(new_n239), .A3(new_n595), .ZN(new_n909));
  XOR2_X1   g708(.A(new_n909), .B(KEYINPUT120), .Z(new_n910));
  AOI21_X1  g709(.A(new_n239), .B1(new_n892), .B2(new_n595), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT61), .Z(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1351gat));
  NAND2_X1  g712(.A1(new_n466), .A2(new_n890), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT121), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n877), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G197gat), .B1(new_n916), .B2(new_n688), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n718), .A2(new_n352), .A3(new_n425), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n887), .A2(new_n919), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n920), .A2(G197gat), .A3(new_n688), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n918), .A3(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(G197gat), .ZN(new_n924));
  INV_X1    g723(.A(new_n915), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n876), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n924), .B1(new_n926), .B2(new_n628), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT122), .B1(new_n927), .B2(new_n921), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n923), .A2(new_n928), .ZN(G1352gat));
  XNOR2_X1  g728(.A(KEYINPUT123), .B(G204gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(new_n916), .B2(new_n663), .ZN(new_n931));
  INV_X1    g730(.A(new_n920), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(new_n662), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n934), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n931), .A2(new_n936), .ZN(G1353gat));
  OR3_X1    g736(.A1(new_n920), .A2(G211gat), .A3(new_n525), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n687), .B(new_n915), .C1(new_n866), .C2(new_n875), .ZN(new_n939));
  AND2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n939), .A2(KEYINPUT125), .A3(new_n940), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n943), .B(new_n944), .C1(KEYINPUT126), .C2(new_n945), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n945), .A2(KEYINPUT126), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n938), .B1(new_n946), .B2(new_n947), .ZN(G1354gat));
  OAI21_X1  g747(.A(G218gat), .B1(new_n916), .B2(new_n685), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n685), .A2(G218gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n920), .B2(new_n950), .ZN(G1355gat));
endmodule


