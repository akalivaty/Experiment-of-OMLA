

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U552 ( .A(KEYINPUT30), .B(KEYINPUT102), .ZN(n641) );
  XNOR2_X1 U553 ( .A(n642), .B(n641), .ZN(n643) );
  INV_X1 U554 ( .A(KEYINPUT29), .ZN(n690) );
  NOR2_X1 U555 ( .A1(n647), .A2(n646), .ZN(n649) );
  INV_X1 U556 ( .A(KEYINPUT104), .ZN(n698) );
  NOR2_X2 U557 ( .A1(n519), .A2(G2105), .ZN(n879) );
  NOR2_X1 U558 ( .A1(G651), .A2(n545), .ZN(n788) );
  NOR2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  XOR2_X1 U560 ( .A(KEYINPUT17), .B(n518), .Z(n880) );
  NAND2_X1 U561 ( .A1(n880), .A2(G137), .ZN(n527) );
  INV_X1 U562 ( .A(G2104), .ZN(n519) );
  NAND2_X1 U563 ( .A1(G101), .A2(n879), .ZN(n520) );
  XNOR2_X1 U564 ( .A(KEYINPUT23), .B(n520), .ZN(n525) );
  NAND2_X1 U565 ( .A1(n519), .A2(G2105), .ZN(n521) );
  XNOR2_X2 U566 ( .A(n521), .B(KEYINPUT65), .ZN(n884) );
  NAND2_X1 U567 ( .A1(G125), .A2(n884), .ZN(n523) );
  AND2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n883) );
  NAND2_X1 U569 ( .A1(G113), .A2(n883), .ZN(n522) );
  NAND2_X1 U570 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U571 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U572 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X2 U573 ( .A(KEYINPUT64), .B(n528), .Z(G160) );
  NAND2_X1 U574 ( .A1(G102), .A2(n879), .ZN(n530) );
  NAND2_X1 U575 ( .A1(G138), .A2(n880), .ZN(n529) );
  NAND2_X1 U576 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U577 ( .A(KEYINPUT92), .B(n531), .ZN(n535) );
  NAND2_X1 U578 ( .A1(G114), .A2(n883), .ZN(n533) );
  NAND2_X1 U579 ( .A1(G126), .A2(n884), .ZN(n532) );
  NAND2_X1 U580 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U581 ( .A1(n535), .A2(n534), .ZN(G164) );
  INV_X1 U582 ( .A(G651), .ZN(n544) );
  NOR2_X1 U583 ( .A1(G543), .A2(n544), .ZN(n536) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n536), .Z(n784) );
  XOR2_X1 U585 ( .A(KEYINPUT0), .B(G543), .Z(n545) );
  NAND2_X1 U586 ( .A1(G87), .A2(n545), .ZN(n537) );
  XNOR2_X1 U587 ( .A(n537), .B(KEYINPUT82), .ZN(n540) );
  NAND2_X1 U588 ( .A1(G74), .A2(G651), .ZN(n538) );
  XOR2_X1 U589 ( .A(KEYINPUT81), .B(n538), .Z(n539) );
  NAND2_X1 U590 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U591 ( .A1(n784), .A2(n541), .ZN(n543) );
  NAND2_X1 U592 ( .A1(n788), .A2(G49), .ZN(n542) );
  NAND2_X1 U593 ( .A1(n543), .A2(n542), .ZN(G288) );
  NOR2_X1 U594 ( .A1(n545), .A2(n544), .ZN(n787) );
  NAND2_X1 U595 ( .A1(n787), .A2(G73), .ZN(n547) );
  XNOR2_X1 U596 ( .A(KEYINPUT2), .B(KEYINPUT84), .ZN(n546) );
  XNOR2_X1 U597 ( .A(n547), .B(n546), .ZN(n554) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n782) );
  NAND2_X1 U599 ( .A1(G86), .A2(n782), .ZN(n549) );
  NAND2_X1 U600 ( .A1(G48), .A2(n788), .ZN(n548) );
  NAND2_X1 U601 ( .A1(n549), .A2(n548), .ZN(n552) );
  NAND2_X1 U602 ( .A1(G61), .A2(n784), .ZN(n550) );
  XNOR2_X1 U603 ( .A(KEYINPUT83), .B(n550), .ZN(n551) );
  NOR2_X1 U604 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U605 ( .A1(n554), .A2(n553), .ZN(G305) );
  NAND2_X1 U606 ( .A1(G63), .A2(n784), .ZN(n556) );
  NAND2_X1 U607 ( .A1(G51), .A2(n788), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U609 ( .A(n557), .B(KEYINPUT77), .ZN(n558) );
  XNOR2_X1 U610 ( .A(n558), .B(KEYINPUT6), .ZN(n565) );
  XNOR2_X1 U611 ( .A(KEYINPUT5), .B(KEYINPUT76), .ZN(n563) );
  NAND2_X1 U612 ( .A1(n782), .A2(G89), .ZN(n559) );
  XNOR2_X1 U613 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U614 ( .A1(G76), .A2(n787), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U616 ( .A(n563), .B(n562), .ZN(n564) );
  NAND2_X1 U617 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U618 ( .A(KEYINPUT7), .B(n566), .ZN(G168) );
  XNOR2_X1 U619 ( .A(KEYINPUT69), .B(KEYINPUT9), .ZN(n570) );
  NAND2_X1 U620 ( .A1(G90), .A2(n782), .ZN(n568) );
  NAND2_X1 U621 ( .A1(G77), .A2(n787), .ZN(n567) );
  NAND2_X1 U622 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U623 ( .A(n570), .B(n569), .ZN(n575) );
  NAND2_X1 U624 ( .A1(n788), .A2(G52), .ZN(n571) );
  XNOR2_X1 U625 ( .A(n571), .B(KEYINPUT68), .ZN(n573) );
  NAND2_X1 U626 ( .A1(G64), .A2(n784), .ZN(n572) );
  NAND2_X1 U627 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U628 ( .A1(n575), .A2(n574), .ZN(G171) );
  NAND2_X1 U629 ( .A1(G91), .A2(n782), .ZN(n577) );
  NAND2_X1 U630 ( .A1(G78), .A2(n787), .ZN(n576) );
  NAND2_X1 U631 ( .A1(n577), .A2(n576), .ZN(n580) );
  NAND2_X1 U632 ( .A1(n784), .A2(G65), .ZN(n578) );
  XOR2_X1 U633 ( .A(KEYINPUT70), .B(n578), .Z(n579) );
  NOR2_X1 U634 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U635 ( .A1(n788), .A2(G53), .ZN(n581) );
  NAND2_X1 U636 ( .A1(n582), .A2(n581), .ZN(G299) );
  NAND2_X1 U637 ( .A1(G88), .A2(n782), .ZN(n584) );
  NAND2_X1 U638 ( .A1(G75), .A2(n787), .ZN(n583) );
  NAND2_X1 U639 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U640 ( .A1(G62), .A2(n784), .ZN(n586) );
  NAND2_X1 U641 ( .A1(G50), .A2(n788), .ZN(n585) );
  NAND2_X1 U642 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U643 ( .A1(n588), .A2(n587), .ZN(G166) );
  INV_X1 U644 ( .A(G166), .ZN(G303) );
  XOR2_X1 U645 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U646 ( .A1(G60), .A2(n784), .ZN(n590) );
  NAND2_X1 U647 ( .A1(G47), .A2(n788), .ZN(n589) );
  NAND2_X1 U648 ( .A1(n590), .A2(n589), .ZN(n595) );
  NAND2_X1 U649 ( .A1(G85), .A2(n782), .ZN(n592) );
  NAND2_X1 U650 ( .A1(G72), .A2(n787), .ZN(n591) );
  NAND2_X1 U651 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U652 ( .A(KEYINPUT66), .B(n593), .ZN(n594) );
  NOR2_X1 U653 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U654 ( .A(n596), .B(KEYINPUT67), .ZN(G290) );
  NOR2_X1 U655 ( .A1(G164), .A2(G1384), .ZN(n630) );
  NAND2_X1 U656 ( .A1(G160), .A2(G40), .ZN(n597) );
  XOR2_X1 U657 ( .A(n597), .B(KEYINPUT93), .Z(n629) );
  NOR2_X1 U658 ( .A1(n630), .A2(n629), .ZN(n750) );
  XNOR2_X1 U659 ( .A(G2067), .B(KEYINPUT37), .ZN(n598) );
  XNOR2_X1 U660 ( .A(n598), .B(KEYINPUT94), .ZN(n748) );
  NAND2_X1 U661 ( .A1(G104), .A2(n879), .ZN(n600) );
  NAND2_X1 U662 ( .A1(G140), .A2(n880), .ZN(n599) );
  NAND2_X1 U663 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U664 ( .A(KEYINPUT34), .B(n601), .ZN(n606) );
  NAND2_X1 U665 ( .A1(G116), .A2(n883), .ZN(n603) );
  NAND2_X1 U666 ( .A1(G128), .A2(n884), .ZN(n602) );
  NAND2_X1 U667 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U668 ( .A(KEYINPUT35), .B(n604), .Z(n605) );
  NOR2_X1 U669 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U670 ( .A(KEYINPUT36), .B(n607), .ZN(n892) );
  NOR2_X1 U671 ( .A1(n748), .A2(n892), .ZN(n973) );
  NAND2_X1 U672 ( .A1(n750), .A2(n973), .ZN(n746) );
  INV_X1 U673 ( .A(n746), .ZN(n627) );
  NAND2_X1 U674 ( .A1(G95), .A2(n879), .ZN(n609) );
  NAND2_X1 U675 ( .A1(G107), .A2(n883), .ZN(n608) );
  NAND2_X1 U676 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U677 ( .A1(G131), .A2(n880), .ZN(n611) );
  NAND2_X1 U678 ( .A1(G119), .A2(n884), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n611), .A2(n610), .ZN(n612) );
  OR2_X1 U680 ( .A1(n613), .A2(n612), .ZN(n865) );
  XOR2_X1 U681 ( .A(KEYINPUT95), .B(G1991), .Z(n946) );
  AND2_X1 U682 ( .A1(n865), .A2(n946), .ZN(n624) );
  NAND2_X1 U683 ( .A1(G105), .A2(n879), .ZN(n614) );
  XOR2_X1 U684 ( .A(KEYINPUT38), .B(n614), .Z(n620) );
  NAND2_X1 U685 ( .A1(n883), .A2(G117), .ZN(n615) );
  XNOR2_X1 U686 ( .A(n615), .B(KEYINPUT96), .ZN(n617) );
  NAND2_X1 U687 ( .A1(G129), .A2(n884), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U689 ( .A(KEYINPUT97), .B(n618), .Z(n619) );
  NOR2_X1 U690 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n880), .A2(G141), .ZN(n621) );
  NAND2_X1 U692 ( .A1(n622), .A2(n621), .ZN(n875) );
  AND2_X1 U693 ( .A1(n875), .A2(G1996), .ZN(n623) );
  NOR2_X1 U694 ( .A1(n624), .A2(n623), .ZN(n971) );
  INV_X1 U695 ( .A(n750), .ZN(n625) );
  NOR2_X1 U696 ( .A1(n971), .A2(n625), .ZN(n743) );
  XNOR2_X1 U697 ( .A(KEYINPUT98), .B(n743), .ZN(n626) );
  NOR2_X1 U698 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n628), .B(KEYINPUT99), .ZN(n737) );
  NOR2_X1 U700 ( .A1(G1976), .A2(G288), .ZN(n997) );
  NAND2_X1 U701 ( .A1(n997), .A2(KEYINPUT33), .ZN(n632) );
  INV_X1 U702 ( .A(n629), .ZN(n631) );
  NAND2_X2 U703 ( .A1(n631), .A2(n630), .ZN(n705) );
  NAND2_X1 U704 ( .A1(G8), .A2(n705), .ZN(n730) );
  NOR2_X1 U705 ( .A1(n632), .A2(n730), .ZN(n634) );
  XOR2_X1 U706 ( .A(G1981), .B(G305), .Z(n1010) );
  INV_X1 U707 ( .A(n1010), .ZN(n633) );
  NOR2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U709 ( .A1(G1976), .A2(G288), .ZN(n1001) );
  INV_X1 U710 ( .A(n1001), .ZN(n635) );
  NOR2_X1 U711 ( .A1(n730), .A2(n635), .ZN(n636) );
  OR2_X1 U712 ( .A1(KEYINPUT33), .A2(n636), .ZN(n637) );
  AND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n722) );
  NOR2_X1 U714 ( .A1(G2084), .A2(n705), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G8), .A2(n639), .ZN(n704) );
  NOR2_X1 U716 ( .A1(G1966), .A2(n730), .ZN(n699) );
  NOR2_X1 U717 ( .A1(n639), .A2(n699), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n640), .A2(G8), .ZN(n642) );
  NOR2_X1 U719 ( .A1(G168), .A2(n643), .ZN(n647) );
  XNOR2_X1 U720 ( .A(G2078), .B(KEYINPUT25), .ZN(n948) );
  NOR2_X1 U721 ( .A1(n705), .A2(n948), .ZN(n645) );
  AND2_X1 U722 ( .A1(n705), .A2(G1961), .ZN(n644) );
  NOR2_X1 U723 ( .A1(n645), .A2(n644), .ZN(n692) );
  NOR2_X1 U724 ( .A1(G171), .A2(n692), .ZN(n646) );
  XNOR2_X1 U725 ( .A(KEYINPUT103), .B(KEYINPUT31), .ZN(n648) );
  XNOR2_X1 U726 ( .A(n649), .B(n648), .ZN(n697) );
  NAND2_X1 U727 ( .A1(G92), .A2(n782), .ZN(n651) );
  NAND2_X1 U728 ( .A1(G66), .A2(n784), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U730 ( .A1(G79), .A2(n787), .ZN(n653) );
  NAND2_X1 U731 ( .A1(G54), .A2(n788), .ZN(n652) );
  NAND2_X1 U732 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U733 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U734 ( .A(KEYINPUT15), .B(n656), .Z(n993) );
  INV_X1 U735 ( .A(n993), .ZN(n777) );
  NOR2_X1 U736 ( .A1(G2067), .A2(n705), .ZN(n658) );
  INV_X1 U737 ( .A(n705), .ZN(n680) );
  NOR2_X1 U738 ( .A1(n680), .A2(G1348), .ZN(n657) );
  NOR2_X1 U739 ( .A1(n658), .A2(n657), .ZN(n676) );
  NAND2_X1 U740 ( .A1(n777), .A2(n676), .ZN(n675) );
  INV_X1 U741 ( .A(G1996), .ZN(n954) );
  NOR2_X1 U742 ( .A1(n705), .A2(n954), .ZN(n659) );
  XOR2_X1 U743 ( .A(n659), .B(KEYINPUT26), .Z(n673) );
  AND2_X1 U744 ( .A1(n705), .A2(G1341), .ZN(n671) );
  NAND2_X1 U745 ( .A1(G56), .A2(n784), .ZN(n660) );
  XOR2_X1 U746 ( .A(KEYINPUT14), .B(n660), .Z(n668) );
  XOR2_X1 U747 ( .A(KEYINPUT12), .B(KEYINPUT72), .Z(n662) );
  NAND2_X1 U748 ( .A1(G81), .A2(n782), .ZN(n661) );
  XNOR2_X1 U749 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U750 ( .A(KEYINPUT71), .B(n663), .ZN(n665) );
  NAND2_X1 U751 ( .A1(n787), .A2(G68), .ZN(n664) );
  NAND2_X1 U752 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U753 ( .A(KEYINPUT13), .B(n666), .Z(n667) );
  NOR2_X1 U754 ( .A1(n668), .A2(n667), .ZN(n670) );
  NAND2_X1 U755 ( .A1(n788), .A2(G43), .ZN(n669) );
  NAND2_X1 U756 ( .A1(n670), .A2(n669), .ZN(n1007) );
  NOR2_X1 U757 ( .A1(n671), .A2(n1007), .ZN(n672) );
  AND2_X1 U758 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n675), .A2(n674), .ZN(n678) );
  OR2_X1 U760 ( .A1(n676), .A2(n777), .ZN(n677) );
  NAND2_X1 U761 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U762 ( .A(n679), .B(KEYINPUT101), .ZN(n685) );
  NAND2_X1 U763 ( .A1(n680), .A2(G2072), .ZN(n681) );
  XNOR2_X1 U764 ( .A(n681), .B(KEYINPUT27), .ZN(n683) );
  AND2_X1 U765 ( .A1(G1956), .A2(n705), .ZN(n682) );
  NOR2_X1 U766 ( .A1(n683), .A2(n682), .ZN(n686) );
  INV_X1 U767 ( .A(G299), .ZN(n800) );
  NAND2_X1 U768 ( .A1(n686), .A2(n800), .ZN(n684) );
  NAND2_X1 U769 ( .A1(n685), .A2(n684), .ZN(n689) );
  NOR2_X1 U770 ( .A1(n686), .A2(n800), .ZN(n687) );
  XOR2_X1 U771 ( .A(n687), .B(KEYINPUT28), .Z(n688) );
  NAND2_X1 U772 ( .A1(n689), .A2(n688), .ZN(n691) );
  XNOR2_X1 U773 ( .A(n691), .B(n690), .ZN(n695) );
  AND2_X1 U774 ( .A1(G171), .A2(n692), .ZN(n693) );
  XOR2_X1 U775 ( .A(KEYINPUT100), .B(n693), .Z(n694) );
  NAND2_X1 U776 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U777 ( .A1(n697), .A2(n696), .ZN(n709) );
  XNOR2_X1 U778 ( .A(n709), .B(n698), .ZN(n700) );
  NOR2_X1 U779 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U780 ( .A(KEYINPUT105), .B(n701), .ZN(n702) );
  INV_X1 U781 ( .A(n702), .ZN(n703) );
  NAND2_X1 U782 ( .A1(n704), .A2(n703), .ZN(n715) );
  NOR2_X1 U783 ( .A1(G1971), .A2(n730), .ZN(n707) );
  NOR2_X1 U784 ( .A1(G2090), .A2(n705), .ZN(n706) );
  NOR2_X1 U785 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U786 ( .A1(n708), .A2(G303), .ZN(n711) );
  NAND2_X1 U787 ( .A1(n709), .A2(G286), .ZN(n710) );
  NAND2_X1 U788 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U789 ( .A1(G8), .A2(n712), .ZN(n713) );
  XNOR2_X1 U790 ( .A(KEYINPUT32), .B(n713), .ZN(n714) );
  NAND2_X1 U791 ( .A1(n715), .A2(n714), .ZN(n728) );
  NOR2_X1 U792 ( .A1(G1971), .A2(G303), .ZN(n716) );
  NOR2_X1 U793 ( .A1(n997), .A2(n716), .ZN(n717) );
  XNOR2_X1 U794 ( .A(n717), .B(KEYINPUT106), .ZN(n719) );
  INV_X1 U795 ( .A(KEYINPUT33), .ZN(n718) );
  AND2_X1 U796 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U797 ( .A1(n728), .A2(n720), .ZN(n721) );
  NAND2_X1 U798 ( .A1(n722), .A2(n721), .ZN(n735) );
  NOR2_X1 U799 ( .A1(G2090), .A2(G303), .ZN(n723) );
  NAND2_X1 U800 ( .A1(G8), .A2(n723), .ZN(n726) );
  NOR2_X1 U801 ( .A1(G1981), .A2(G305), .ZN(n724) );
  XOR2_X1 U802 ( .A(n724), .B(KEYINPUT24), .Z(n725) );
  OR2_X1 U803 ( .A1(n730), .A2(n725), .ZN(n729) );
  AND2_X1 U804 ( .A1(n726), .A2(n729), .ZN(n727) );
  NAND2_X1 U805 ( .A1(n728), .A2(n727), .ZN(n733) );
  INV_X1 U806 ( .A(n729), .ZN(n731) );
  OR2_X1 U807 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U808 ( .A1(n733), .A2(n732), .ZN(n734) );
  AND2_X1 U809 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U810 ( .A1(n737), .A2(n736), .ZN(n739) );
  XNOR2_X1 U811 ( .A(G1986), .B(G290), .ZN(n1003) );
  NAND2_X1 U812 ( .A1(n1003), .A2(n750), .ZN(n738) );
  NAND2_X1 U813 ( .A1(n739), .A2(n738), .ZN(n753) );
  NOR2_X1 U814 ( .A1(G1996), .A2(n875), .ZN(n968) );
  NOR2_X1 U815 ( .A1(n946), .A2(n865), .ZN(n977) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n740) );
  NOR2_X1 U817 ( .A1(n977), .A2(n740), .ZN(n741) );
  XOR2_X1 U818 ( .A(KEYINPUT107), .B(n741), .Z(n742) );
  NOR2_X1 U819 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U820 ( .A1(n968), .A2(n744), .ZN(n745) );
  XNOR2_X1 U821 ( .A(KEYINPUT39), .B(n745), .ZN(n747) );
  NAND2_X1 U822 ( .A1(n747), .A2(n746), .ZN(n749) );
  NAND2_X1 U823 ( .A1(n748), .A2(n892), .ZN(n970) );
  NAND2_X1 U824 ( .A1(n749), .A2(n970), .ZN(n751) );
  NAND2_X1 U825 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n755) );
  XNOR2_X1 U827 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n754) );
  XNOR2_X1 U828 ( .A(n755), .B(n754), .ZN(G329) );
  AND2_X1 U829 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U830 ( .A1(G99), .A2(n879), .ZN(n757) );
  NAND2_X1 U831 ( .A1(G111), .A2(n883), .ZN(n756) );
  NAND2_X1 U832 ( .A1(n757), .A2(n756), .ZN(n760) );
  NAND2_X1 U833 ( .A1(n884), .A2(G123), .ZN(n758) );
  XOR2_X1 U834 ( .A(KEYINPUT18), .B(n758), .Z(n759) );
  NOR2_X1 U835 ( .A1(n760), .A2(n759), .ZN(n762) );
  NAND2_X1 U836 ( .A1(n880), .A2(G135), .ZN(n761) );
  NAND2_X1 U837 ( .A1(n762), .A2(n761), .ZN(n974) );
  XNOR2_X1 U838 ( .A(G2096), .B(n974), .ZN(n763) );
  OR2_X1 U839 ( .A1(G2100), .A2(n763), .ZN(G156) );
  INV_X1 U840 ( .A(G57), .ZN(G237) );
  NAND2_X1 U841 ( .A1(G7), .A2(G661), .ZN(n764) );
  XNOR2_X1 U842 ( .A(n764), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U843 ( .A(G223), .ZN(n828) );
  NAND2_X1 U844 ( .A1(n828), .A2(G567), .ZN(n765) );
  XOR2_X1 U845 ( .A(KEYINPUT11), .B(n765), .Z(G234) );
  INV_X1 U846 ( .A(n1007), .ZN(n766) );
  INV_X1 U847 ( .A(G860), .ZN(n794) );
  XNOR2_X1 U848 ( .A(KEYINPUT73), .B(n794), .ZN(n774) );
  NAND2_X1 U849 ( .A1(n766), .A2(n774), .ZN(G153) );
  NOR2_X1 U850 ( .A1(n993), .A2(G868), .ZN(n767) );
  XNOR2_X1 U851 ( .A(n767), .B(KEYINPUT74), .ZN(n769) );
  INV_X1 U852 ( .A(G868), .ZN(n807) );
  NOR2_X1 U853 ( .A1(n807), .A2(G171), .ZN(n768) );
  NOR2_X1 U854 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U855 ( .A(KEYINPUT75), .B(n770), .ZN(G284) );
  INV_X1 U856 ( .A(G171), .ZN(G301) );
  NOR2_X1 U857 ( .A1(G286), .A2(n807), .ZN(n772) );
  NOR2_X1 U858 ( .A1(G868), .A2(G299), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n772), .A2(n771), .ZN(G297) );
  INV_X1 U860 ( .A(G559), .ZN(n773) );
  NOR2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U862 ( .A1(n777), .A2(n775), .ZN(n776) );
  XOR2_X1 U863 ( .A(KEYINPUT16), .B(n776), .Z(G148) );
  NOR2_X1 U864 ( .A1(n777), .A2(n807), .ZN(n778) );
  XOR2_X1 U865 ( .A(KEYINPUT78), .B(n778), .Z(n779) );
  NOR2_X1 U866 ( .A1(G559), .A2(n779), .ZN(n781) );
  NOR2_X1 U867 ( .A1(G868), .A2(n1007), .ZN(n780) );
  NOR2_X1 U868 ( .A1(n781), .A2(n780), .ZN(G282) );
  NAND2_X1 U869 ( .A1(n782), .A2(G93), .ZN(n783) );
  XNOR2_X1 U870 ( .A(n783), .B(KEYINPUT80), .ZN(n786) );
  NAND2_X1 U871 ( .A1(G67), .A2(n784), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n792) );
  NAND2_X1 U873 ( .A1(G80), .A2(n787), .ZN(n790) );
  NAND2_X1 U874 ( .A1(G55), .A2(n788), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n790), .A2(n789), .ZN(n791) );
  OR2_X1 U876 ( .A1(n792), .A2(n791), .ZN(n808) );
  NAND2_X1 U877 ( .A1(G559), .A2(n993), .ZN(n793) );
  XOR2_X1 U878 ( .A(n1007), .B(n793), .Z(n804) );
  NAND2_X1 U879 ( .A1(n804), .A2(n794), .ZN(n795) );
  XNOR2_X1 U880 ( .A(KEYINPUT79), .B(n795), .ZN(n796) );
  XOR2_X1 U881 ( .A(n808), .B(n796), .Z(G145) );
  XOR2_X1 U882 ( .A(n808), .B(G288), .Z(n803) );
  XNOR2_X1 U883 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n798) );
  XNOR2_X1 U884 ( .A(G290), .B(G166), .ZN(n797) );
  XNOR2_X1 U885 ( .A(n798), .B(n797), .ZN(n799) );
  XNOR2_X1 U886 ( .A(n800), .B(n799), .ZN(n801) );
  XNOR2_X1 U887 ( .A(n801), .B(G305), .ZN(n802) );
  XNOR2_X1 U888 ( .A(n803), .B(n802), .ZN(n896) );
  XNOR2_X1 U889 ( .A(n804), .B(n896), .ZN(n805) );
  XNOR2_X1 U890 ( .A(KEYINPUT86), .B(n805), .ZN(n806) );
  NOR2_X1 U891 ( .A1(n807), .A2(n806), .ZN(n810) );
  NOR2_X1 U892 ( .A1(G868), .A2(n808), .ZN(n809) );
  NOR2_X1 U893 ( .A1(n810), .A2(n809), .ZN(G295) );
  NAND2_X1 U894 ( .A1(G2084), .A2(G2078), .ZN(n811) );
  XNOR2_X1 U895 ( .A(n811), .B(KEYINPUT87), .ZN(n812) );
  XNOR2_X1 U896 ( .A(n812), .B(KEYINPUT20), .ZN(n813) );
  NAND2_X1 U897 ( .A1(n813), .A2(G2090), .ZN(n814) );
  XNOR2_X1 U898 ( .A(n814), .B(KEYINPUT21), .ZN(n815) );
  XNOR2_X1 U899 ( .A(n815), .B(KEYINPUT88), .ZN(n816) );
  NAND2_X1 U900 ( .A1(n816), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U901 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U902 ( .A1(G69), .A2(G120), .ZN(n817) );
  NOR2_X1 U903 ( .A1(G237), .A2(n817), .ZN(n818) );
  NAND2_X1 U904 ( .A1(G108), .A2(n818), .ZN(n835) );
  NAND2_X1 U905 ( .A1(G567), .A2(n835), .ZN(n825) );
  XOR2_X1 U906 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n820) );
  NAND2_X1 U907 ( .A1(G132), .A2(G82), .ZN(n819) );
  XNOR2_X1 U908 ( .A(n820), .B(n819), .ZN(n821) );
  NOR2_X1 U909 ( .A1(n821), .A2(G218), .ZN(n822) );
  XNOR2_X1 U910 ( .A(KEYINPUT90), .B(n822), .ZN(n823) );
  NAND2_X1 U911 ( .A1(n823), .A2(G96), .ZN(n834) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n834), .ZN(n824) );
  NAND2_X1 U913 ( .A1(n825), .A2(n824), .ZN(n836) );
  NAND2_X1 U914 ( .A1(G483), .A2(G661), .ZN(n826) );
  NOR2_X1 U915 ( .A1(n836), .A2(n826), .ZN(n831) );
  NAND2_X1 U916 ( .A1(n831), .A2(G36), .ZN(n827) );
  XOR2_X1 U917 ( .A(KEYINPUT91), .B(n827), .Z(G176) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n828), .ZN(G217) );
  NAND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n829) );
  XOR2_X1 U920 ( .A(KEYINPUT110), .B(n829), .Z(n830) );
  NAND2_X1 U921 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U923 ( .A1(n832), .A2(n831), .ZN(n833) );
  XOR2_X1 U924 ( .A(KEYINPUT111), .B(n833), .Z(G188) );
  NOR2_X1 U925 ( .A1(n835), .A2(n834), .ZN(G325) );
  XOR2_X1 U926 ( .A(KEYINPUT112), .B(G325), .Z(G261) );
  INV_X1 U927 ( .A(n836), .ZN(G319) );
  XOR2_X1 U928 ( .A(G2100), .B(G2096), .Z(n838) );
  XNOR2_X1 U929 ( .A(KEYINPUT42), .B(G2678), .ZN(n837) );
  XNOR2_X1 U930 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U931 ( .A(KEYINPUT43), .B(G2090), .Z(n840) );
  XNOR2_X1 U932 ( .A(G2067), .B(G2072), .ZN(n839) );
  XNOR2_X1 U933 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U934 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U935 ( .A(G2084), .B(G2078), .ZN(n843) );
  XNOR2_X1 U936 ( .A(n844), .B(n843), .ZN(G227) );
  XOR2_X1 U937 ( .A(KEYINPUT114), .B(G1981), .Z(n846) );
  XNOR2_X1 U938 ( .A(G1956), .B(G1961), .ZN(n845) );
  XNOR2_X1 U939 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U940 ( .A(n847), .B(KEYINPUT41), .Z(n849) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U942 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U943 ( .A(G1976), .B(G1971), .Z(n851) );
  XNOR2_X1 U944 ( .A(G1986), .B(G1966), .ZN(n850) );
  XNOR2_X1 U945 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U946 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U947 ( .A(KEYINPUT113), .B(G2474), .ZN(n854) );
  XNOR2_X1 U948 ( .A(n855), .B(n854), .ZN(G229) );
  NAND2_X1 U949 ( .A1(G100), .A2(n879), .ZN(n857) );
  NAND2_X1 U950 ( .A1(G112), .A2(n883), .ZN(n856) );
  NAND2_X1 U951 ( .A1(n857), .A2(n856), .ZN(n862) );
  NAND2_X1 U952 ( .A1(G124), .A2(n884), .ZN(n858) );
  XNOR2_X1 U953 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U954 ( .A1(n880), .A2(G136), .ZN(n859) );
  NAND2_X1 U955 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U956 ( .A1(n862), .A2(n861), .ZN(G162) );
  XNOR2_X1 U957 ( .A(G162), .B(G160), .ZN(n863) );
  XNOR2_X1 U958 ( .A(n863), .B(n974), .ZN(n864) );
  XOR2_X1 U959 ( .A(n864), .B(KEYINPUT48), .Z(n867) );
  XOR2_X1 U960 ( .A(n865), .B(KEYINPUT46), .Z(n866) );
  XNOR2_X1 U961 ( .A(n867), .B(n866), .ZN(n878) );
  NAND2_X1 U962 ( .A1(G118), .A2(n883), .ZN(n869) );
  NAND2_X1 U963 ( .A1(G130), .A2(n884), .ZN(n868) );
  NAND2_X1 U964 ( .A1(n869), .A2(n868), .ZN(n874) );
  NAND2_X1 U965 ( .A1(G106), .A2(n879), .ZN(n871) );
  NAND2_X1 U966 ( .A1(G142), .A2(n880), .ZN(n870) );
  NAND2_X1 U967 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U968 ( .A(n872), .B(KEYINPUT45), .Z(n873) );
  NOR2_X1 U969 ( .A1(n874), .A2(n873), .ZN(n876) );
  XNOR2_X1 U970 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U971 ( .A(n878), .B(n877), .Z(n891) );
  NAND2_X1 U972 ( .A1(G103), .A2(n879), .ZN(n882) );
  NAND2_X1 U973 ( .A1(G139), .A2(n880), .ZN(n881) );
  NAND2_X1 U974 ( .A1(n882), .A2(n881), .ZN(n889) );
  NAND2_X1 U975 ( .A1(G115), .A2(n883), .ZN(n886) );
  NAND2_X1 U976 ( .A1(G127), .A2(n884), .ZN(n885) );
  NAND2_X1 U977 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U978 ( .A(KEYINPUT47), .B(n887), .Z(n888) );
  NOR2_X1 U979 ( .A1(n889), .A2(n888), .ZN(n981) );
  XNOR2_X1 U980 ( .A(G164), .B(n981), .ZN(n890) );
  XNOR2_X1 U981 ( .A(n891), .B(n890), .ZN(n893) );
  XNOR2_X1 U982 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U983 ( .A1(G37), .A2(n894), .ZN(G395) );
  XNOR2_X1 U984 ( .A(n993), .B(G171), .ZN(n895) );
  XNOR2_X1 U985 ( .A(n895), .B(G286), .ZN(n898) );
  XNOR2_X1 U986 ( .A(n1007), .B(n896), .ZN(n897) );
  XNOR2_X1 U987 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U988 ( .A1(G37), .A2(n899), .ZN(G397) );
  XOR2_X1 U989 ( .A(G2454), .B(G2430), .Z(n901) );
  XNOR2_X1 U990 ( .A(G2451), .B(G2446), .ZN(n900) );
  XNOR2_X1 U991 ( .A(n901), .B(n900), .ZN(n908) );
  XOR2_X1 U992 ( .A(G2443), .B(G2427), .Z(n903) );
  XNOR2_X1 U993 ( .A(G2438), .B(KEYINPUT109), .ZN(n902) );
  XNOR2_X1 U994 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U995 ( .A(n904), .B(G2435), .Z(n906) );
  XNOR2_X1 U996 ( .A(G1348), .B(G1341), .ZN(n905) );
  XNOR2_X1 U997 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U998 ( .A(n908), .B(n907), .ZN(n909) );
  NAND2_X1 U999 ( .A1(n909), .A2(G14), .ZN(n915) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n915), .ZN(n912) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1003 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1005 ( .A1(n914), .A2(n913), .ZN(G225) );
  XNOR2_X1 U1006 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  INV_X1 U1008 ( .A(G132), .ZN(G219) );
  INV_X1 U1009 ( .A(G120), .ZN(G236) );
  INV_X1 U1010 ( .A(G96), .ZN(G221) );
  INV_X1 U1011 ( .A(G82), .ZN(G220) );
  INV_X1 U1012 ( .A(G69), .ZN(G235) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(n915), .ZN(G401) );
  XOR2_X1 U1015 ( .A(G16), .B(KEYINPUT124), .Z(n940) );
  XNOR2_X1 U1016 ( .A(G1956), .B(G20), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(G1981), .B(G6), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n924) );
  XOR2_X1 U1019 ( .A(KEYINPUT126), .B(G4), .Z(n919) );
  XNOR2_X1 U1020 ( .A(G1348), .B(KEYINPUT59), .ZN(n918) );
  XNOR2_X1 U1021 ( .A(n919), .B(n918), .ZN(n922) );
  XOR2_X1 U1022 ( .A(KEYINPUT125), .B(G1341), .Z(n920) );
  XNOR2_X1 U1023 ( .A(G19), .B(n920), .ZN(n921) );
  NOR2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1026 ( .A(KEYINPUT60), .B(n925), .Z(n936) );
  XOR2_X1 U1027 ( .A(G1966), .B(G21), .Z(n927) );
  XOR2_X1 U1028 ( .A(G1961), .B(G5), .Z(n926) );
  NAND2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(G1971), .B(G22), .ZN(n929) );
  XNOR2_X1 U1031 ( .A(G23), .B(G1976), .ZN(n928) );
  NOR2_X1 U1032 ( .A1(n929), .A2(n928), .ZN(n931) );
  XOR2_X1 U1033 ( .A(G1986), .B(G24), .Z(n930) );
  NAND2_X1 U1034 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1035 ( .A(KEYINPUT58), .B(n932), .ZN(n933) );
  NOR2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(n937), .B(KEYINPUT127), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(n938), .B(KEYINPUT61), .ZN(n939) );
  NAND2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1041 ( .A1(G11), .A2(n941), .ZN(n966) );
  XOR2_X1 U1042 ( .A(G2090), .B(G35), .Z(n945) );
  XNOR2_X1 U1043 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n942) );
  XNOR2_X1 U1044 ( .A(n942), .B(G34), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(G2084), .B(n943), .ZN(n944) );
  NAND2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n962) );
  XOR2_X1 U1047 ( .A(G25), .B(n946), .Z(n959) );
  XNOR2_X1 U1048 ( .A(KEYINPUT117), .B(G2072), .ZN(n947) );
  XNOR2_X1 U1049 ( .A(n947), .B(G33), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(G27), .B(n948), .ZN(n949) );
  NAND2_X1 U1051 ( .A1(n949), .A2(G28), .ZN(n951) );
  XNOR2_X1 U1052 ( .A(G26), .B(G2067), .ZN(n950) );
  NOR2_X1 U1053 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1054 ( .A1(n953), .A2(n952), .ZN(n957) );
  XOR2_X1 U1055 ( .A(G32), .B(n954), .Z(n955) );
  XNOR2_X1 U1056 ( .A(KEYINPUT118), .B(n955), .ZN(n956) );
  NOR2_X1 U1057 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1059 ( .A(KEYINPUT53), .B(n960), .Z(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1061 ( .A1(G29), .A2(n963), .ZN(n964) );
  XOR2_X1 U1062 ( .A(KEYINPUT55), .B(n964), .Z(n965) );
  NOR2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n992) );
  XOR2_X1 U1064 ( .A(G2090), .B(G162), .Z(n967) );
  NOR2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1066 ( .A(KEYINPUT51), .B(n969), .Z(n988) );
  NAND2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G160), .B(G2084), .ZN(n975) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(n978), .B(KEYINPUT116), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n986) );
  XOR2_X1 U1074 ( .A(G2072), .B(n981), .Z(n983) );
  XOR2_X1 U1075 ( .A(G164), .B(G2078), .Z(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1077 ( .A(KEYINPUT50), .B(n984), .Z(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(KEYINPUT52), .B(n989), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n990), .A2(G29), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n1021) );
  XOR2_X1 U1083 ( .A(G16), .B(KEYINPUT56), .Z(n1018) );
  XOR2_X1 U1084 ( .A(G1348), .B(n993), .Z(n995) );
  XNOR2_X1 U1085 ( .A(G301), .B(G1961), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(KEYINPUT120), .B(n996), .ZN(n1006) );
  XOR2_X1 U1088 ( .A(n997), .B(KEYINPUT121), .Z(n999) );
  XOR2_X1 U1089 ( .A(G166), .B(G1971), .Z(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(KEYINPUT122), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1016) );
  XNOR2_X1 U1095 ( .A(G299), .B(G1956), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(n1007), .B(G1341), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(G1966), .B(G168), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(n1012), .B(KEYINPUT57), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1104 ( .A(KEYINPUT123), .B(n1019), .Z(n1020) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1022), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

