//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  NAND2_X1  g000(.A1(KEYINPUT18), .A2(G131), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT85), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT70), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G237), .ZN(new_n192));
  INV_X1    g006(.A(G237), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(KEYINPUT70), .ZN(new_n194));
  OAI211_X1 g008(.A(G214), .B(new_n190), .C1(new_n192), .C2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT85), .A2(G143), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n189), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n189), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(KEYINPUT70), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n191), .A2(G237), .ZN(new_n200));
  AOI21_X1  g014(.A(G953), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n198), .B1(new_n201), .B2(G214), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n188), .B1(new_n197), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT86), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI211_X1 g019(.A(KEYINPUT86), .B(new_n188), .C1(new_n197), .C2(new_n202), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n195), .A2(new_n189), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n201), .A2(G214), .B1(KEYINPUT85), .B2(G143), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n208), .B(new_n187), .C1(new_n209), .C2(new_n189), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT87), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n195), .A2(new_n196), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n198), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n214), .A2(KEYINPUT87), .A3(new_n187), .A4(new_n208), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G140), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G125), .ZN(new_n218));
  INV_X1    g032(.A(G125), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G140), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n207), .A2(new_n216), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(G131), .B1(new_n197), .B2(new_n202), .ZN(new_n225));
  INV_X1    g039(.A(G131), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n208), .B(new_n226), .C1(new_n209), .C2(new_n189), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT17), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT74), .B1(new_n218), .B2(KEYINPUT16), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n218), .A2(new_n220), .A3(KEYINPUT16), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT74), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT16), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n232), .A2(new_n233), .A3(new_n217), .A4(G125), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n235), .A2(new_n222), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT89), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n230), .A2(new_n231), .A3(G146), .A4(new_n234), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  OAI211_X1 g054(.A(KEYINPUT17), .B(G131), .C1(new_n197), .C2(new_n202), .ZN(new_n241));
  INV_X1    g055(.A(new_n239), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT89), .B1(new_n236), .B2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n229), .A2(new_n240), .A3(new_n241), .A4(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(G113), .B(G122), .ZN(new_n245));
  INV_X1    g059(.A(G104), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(KEYINPUT88), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n224), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT90), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT90), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n224), .A2(new_n251), .A3(new_n244), .A4(new_n248), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT91), .ZN(new_n254));
  AOI211_X1 g068(.A(new_n254), .B(new_n247), .C1(new_n224), .C2(new_n244), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n224), .A2(new_n244), .ZN(new_n257));
  INV_X1    g071(.A(new_n247), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n254), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n253), .A2(new_n256), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G902), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT92), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT91), .B1(new_n257), .B2(new_n258), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(new_n255), .ZN(new_n267));
  AOI21_X1  g081(.A(G902), .B1(new_n267), .B2(new_n253), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT92), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n265), .A2(G475), .A3(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(KEYINPUT9), .B(G234), .Z(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(G217), .A3(new_n190), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G116), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G122), .ZN(new_n275));
  OR2_X1    g089(.A1(KEYINPUT66), .A2(G116), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT66), .A2(G116), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n275), .B1(new_n278), .B2(G122), .ZN(new_n279));
  XOR2_X1   g093(.A(KEYINPUT93), .B(G107), .Z(new_n280));
  OR2_X1    g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  XNOR2_X1  g096(.A(G128), .B(G143), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n279), .A2(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G143), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT13), .B1(new_n285), .B2(G128), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT94), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G128), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G143), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n285), .A2(KEYINPUT13), .A3(G128), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n290), .B(new_n291), .C1(new_n286), .C2(KEYINPUT94), .ZN(new_n292));
  OAI21_X1  g106(.A(G134), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n281), .A2(new_n284), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT95), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n281), .A2(new_n284), .A3(KEYINPUT95), .A4(new_n293), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT14), .ZN(new_n299));
  OAI21_X1  g113(.A(G107), .B1(new_n275), .B2(new_n299), .ZN(new_n300));
  OR2_X1    g114(.A1(new_n279), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n283), .B(new_n282), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n279), .A2(new_n300), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n273), .B1(new_n298), .B2(new_n305), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n272), .B(new_n304), .C1(new_n296), .C2(new_n297), .ZN(new_n307));
  OR2_X1    g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT96), .ZN(new_n309));
  INV_X1    g123(.A(G478), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(KEYINPUT15), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n308), .A2(new_n309), .A3(new_n262), .A4(new_n312), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n309), .B(new_n262), .C1(new_n306), .C2(new_n307), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n311), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT97), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n225), .A2(new_n227), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n221), .B(KEYINPUT19), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n242), .B1(new_n319), .B2(new_n222), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n224), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n258), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n253), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT20), .ZN(new_n325));
  INV_X1    g139(.A(G475), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .A4(new_n262), .ZN(new_n327));
  XOR2_X1   g141(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n328));
  AOI22_X1  g142(.A1(new_n250), .A2(new_n252), .B1(new_n258), .B2(new_n322), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(new_n262), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n270), .A2(new_n317), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G221), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n271), .B2(new_n262), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n222), .A2(G143), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n285), .A2(G146), .ZN(new_n339));
  AOI21_X1  g153(.A(G128), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n285), .A2(KEYINPUT1), .A3(G146), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n337), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT1), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n338), .A2(new_n339), .A3(new_n344), .A4(G128), .ZN(new_n345));
  XNOR2_X1  g159(.A(G143), .B(G146), .ZN(new_n346));
  OAI211_X1 g160(.A(KEYINPUT78), .B(new_n341), .C1(new_n346), .C2(G128), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G101), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n246), .A2(G107), .ZN(new_n350));
  INV_X1    g164(.A(G107), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(KEYINPUT3), .A3(G104), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT3), .B1(new_n351), .B2(G104), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n349), .B(new_n350), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n351), .B2(G104), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n351), .A2(G104), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n246), .A2(KEYINPUT77), .A3(G107), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G101), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n348), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n341), .B1(new_n346), .B2(G128), .ZN(new_n365));
  INV_X1    g179(.A(new_n345), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(new_n364), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n363), .A2(new_n364), .B1(new_n368), .B2(new_n362), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT11), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n282), .B2(G137), .ZN(new_n371));
  INV_X1    g185(.A(G137), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(KEYINPUT11), .A3(G134), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n282), .A2(G137), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G131), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n371), .A2(new_n373), .A3(new_n226), .A4(new_n374), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G101), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(KEYINPUT4), .A3(new_n355), .ZN(new_n382));
  NAND2_X1  g196(.A1(KEYINPUT0), .A2(G128), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n338), .A2(new_n339), .A3(new_n383), .ZN(new_n384));
  XOR2_X1   g198(.A(KEYINPUT0), .B(G128), .Z(new_n385));
  OAI21_X1  g199(.A(new_n384), .B1(new_n385), .B2(new_n346), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n380), .A2(new_n387), .A3(G101), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n382), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n369), .A2(new_n379), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n355), .A2(new_n361), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n367), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n363), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT12), .B1(new_n393), .B2(new_n378), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT12), .ZN(new_n395));
  AOI211_X1 g209(.A(new_n395), .B(new_n379), .C1(new_n363), .C2(new_n392), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n390), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT79), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT79), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n390), .B(new_n399), .C1(new_n396), .C2(new_n394), .ZN(new_n400));
  XNOR2_X1  g214(.A(G110), .B(G140), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n190), .A2(G227), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n398), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n369), .A2(new_n379), .A3(new_n389), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n379), .B1(new_n369), .B2(new_n389), .ZN(new_n407));
  OR3_X1    g221(.A1(new_n406), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(G469), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n390), .B(new_n403), .C1(new_n394), .C2(new_n396), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G469), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(new_n262), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(new_n262), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n336), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n333), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT24), .B(G110), .ZN(new_n421));
  INV_X1    g235(.A(G119), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(G128), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n289), .A2(G119), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n421), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT23), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n289), .A2(G119), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT73), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n423), .B2(KEYINPUT23), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n427), .A2(KEYINPUT73), .A3(new_n426), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n425), .B1(new_n432), .B2(G110), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n242), .B2(new_n236), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n421), .B1(new_n423), .B2(new_n424), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n432), .B2(G110), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n221), .A2(new_n222), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n239), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n434), .A2(KEYINPUT75), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT22), .B(G137), .ZN(new_n441));
  INV_X1    g255(.A(G234), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n334), .A2(new_n442), .A3(G953), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n441), .B(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT75), .B1(new_n434), .B2(new_n439), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI211_X1 g261(.A(KEYINPUT75), .B(new_n444), .C1(new_n434), .C2(new_n439), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n262), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT25), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n446), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n440), .A3(new_n444), .ZN(new_n453));
  INV_X1    g267(.A(new_n448), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(KEYINPUT25), .A3(new_n262), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G217), .B1(new_n442), .B2(G902), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n458), .B(KEYINPUT72), .Z(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n262), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n461), .B(KEYINPUT76), .Z(new_n462));
  NAND2_X1  g276(.A1(new_n455), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n201), .A2(G210), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(G101), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT71), .B(KEYINPUT28), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  XOR2_X1   g285(.A(KEYINPUT2), .B(G113), .Z(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT67), .ZN(new_n474));
  AND2_X1   g288(.A1(KEYINPUT66), .A2(G116), .ZN(new_n475));
  NOR2_X1   g289(.A1(KEYINPUT66), .A2(G116), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n474), .B(G119), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT68), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n422), .B1(new_n276), .B2(new_n277), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT67), .B1(new_n422), .B2(G116), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n477), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G119), .B1(new_n475), .B2(new_n476), .ZN(new_n483));
  INV_X1    g297(.A(new_n480), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n478), .B1(new_n485), .B2(new_n477), .ZN(new_n486));
  OAI211_X1 g300(.A(KEYINPUT69), .B(new_n473), .C1(new_n482), .C2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n480), .B1(new_n278), .B2(G119), .ZN(new_n488));
  INV_X1    g302(.A(new_n477), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT68), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n472), .B1(new_n490), .B2(new_n481), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n485), .A2(new_n472), .A3(new_n477), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT69), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n487), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g309(.A1(KEYINPUT0), .A2(G128), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n338), .A2(new_n339), .B1(new_n496), .B2(new_n383), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n338), .A2(new_n339), .A3(new_n383), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT64), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT64), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n500), .B(new_n384), .C1(new_n385), .C2(new_n346), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n378), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n372), .A2(KEYINPUT65), .A3(G134), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT65), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(new_n282), .B2(G137), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n372), .A2(G134), .ZN(new_n506));
  OAI211_X1 g320(.A(G131), .B(new_n503), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n507), .A2(new_n377), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n338), .A2(new_n339), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n289), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n341), .A3(new_n345), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n502), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n495), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n511), .A2(new_n508), .B1(new_n378), .B2(new_n386), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n487), .B(new_n515), .C1(new_n491), .C2(new_n494), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n471), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT28), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n469), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n515), .A2(KEYINPUT30), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n495), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(new_n468), .A3(new_n516), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT31), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT31), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n525), .A2(new_n528), .A3(new_n468), .A4(new_n516), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n521), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(G472), .A2(G902), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n530), .A2(KEYINPUT32), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT32), .B1(new_n530), .B2(new_n531), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n517), .A2(new_n520), .A3(new_n469), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n468), .B1(new_n525), .B2(new_n516), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT29), .ZN(new_n537));
  INV_X1    g351(.A(new_n515), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n495), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n516), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT28), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n519), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n468), .A2(KEYINPUT29), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n262), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(G472), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n464), .B1(new_n534), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(G210), .B1(G237), .B2(G902), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(G110), .B(G122), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n382), .A2(new_n388), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n473), .B1(new_n482), .B2(new_n486), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n493), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n551), .B1(new_n553), .B2(new_n487), .ZN(new_n554));
  INV_X1    g368(.A(new_n492), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n490), .A2(KEYINPUT5), .A3(new_n481), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n274), .A2(KEYINPUT5), .A3(G119), .ZN(new_n557));
  INV_X1    g371(.A(G113), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI211_X1 g373(.A(new_n555), .B(new_n391), .C1(new_n556), .C2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n550), .B1(new_n554), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n551), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n495), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n555), .B1(new_n556), .B2(new_n559), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n362), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n549), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n561), .A2(new_n566), .A3(KEYINPUT6), .ZN(new_n567));
  INV_X1    g381(.A(G224), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(G953), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT80), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n510), .A2(new_n219), .A3(new_n341), .A4(new_n345), .ZN(new_n572));
  OAI211_X1 g386(.A(G125), .B(new_n384), .C1(new_n385), .C2(new_n346), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n573), .A2(new_n571), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n570), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n574), .A2(new_n576), .A3(new_n569), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT6), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n581), .B(new_n550), .C1(new_n554), .C2(new_n560), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n567), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT82), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n549), .B(KEYINPUT8), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n488), .A2(new_n489), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n477), .B(KEYINPUT5), .C1(new_n479), .C2(new_n480), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n586), .A2(new_n472), .B1(new_n587), .B2(new_n559), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n585), .B1(new_n588), .B2(new_n391), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n391), .B2(new_n564), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n575), .A2(new_n577), .A3(KEYINPUT7), .A4(new_n570), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n572), .A2(new_n573), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT81), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT7), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n569), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n593), .B2(new_n594), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n584), .B1(new_n590), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n597), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n579), .B2(KEYINPUT7), .ZN(new_n601));
  AOI211_X1 g415(.A(new_n555), .B(new_n362), .C1(new_n556), .C2(new_n559), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n601), .B(KEYINPUT82), .C1(new_n602), .C2(new_n589), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n599), .A2(new_n603), .A3(new_n566), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n262), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n548), .B1(new_n583), .B2(new_n605), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n591), .B(new_n597), .C1(new_n602), .C2(new_n589), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n495), .A2(new_n562), .B1(new_n564), .B2(new_n362), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n607), .A2(new_n584), .B1(new_n608), .B2(new_n549), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n609), .B2(new_n603), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n567), .A2(new_n580), .A3(new_n582), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n547), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n606), .A2(KEYINPUT83), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n547), .B1(new_n610), .B2(new_n611), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT83), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n190), .A2(G952), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(G234), .B2(G237), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT21), .B(G898), .Z(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(G234), .A2(G237), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(G902), .A3(G953), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n618), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(G214), .B1(G237), .B2(G902), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n613), .A2(new_n616), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n420), .A2(new_n546), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G101), .ZN(G3));
  NAND2_X1  g444(.A1(new_n527), .A2(new_n529), .ZN(new_n631));
  INV_X1    g445(.A(new_n516), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n553), .A2(new_n487), .B1(new_n512), .B2(new_n502), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n470), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n468), .B1(new_n634), .B2(new_n519), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n531), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(G472), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n530), .B2(new_n262), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT98), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n640), .B1(KEYINPUT98), .B2(new_n639), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n410), .A2(new_n418), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n457), .A2(new_n459), .B1(new_n462), .B2(new_n455), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n336), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(G475), .B1(new_n268), .B2(KEYINPUT92), .ZN(new_n646));
  AOI211_X1 g460(.A(new_n264), .B(G902), .C1(new_n267), .C2(new_n253), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n332), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n304), .B1(new_n296), .B2(new_n297), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n649), .A2(KEYINPUT99), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT33), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n308), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n306), .A2(new_n307), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(KEYINPUT33), .A3(new_n650), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(G478), .A3(new_n262), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n310), .B1(new_n653), .B2(G902), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n648), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n624), .B(new_n626), .C1(new_n606), .C2(new_n612), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n645), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT34), .B(G104), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G6));
  INV_X1    g478(.A(KEYINPUT97), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n316), .B(new_n665), .ZN(new_n666));
  OR3_X1    g480(.A1(new_n329), .A2(new_n328), .A3(new_n330), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n331), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n270), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n645), .A2(new_n670), .A3(new_n661), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  NAND2_X1  g487(.A1(new_n434), .A2(new_n439), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n444), .A2(KEYINPUT36), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n462), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n457), .B2(new_n459), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n641), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n420), .A2(new_n628), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  INV_X1    g497(.A(new_n618), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n622), .A2(G900), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n270), .A2(new_n666), .A3(new_n668), .A4(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n418), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n335), .B1(new_n688), .B2(new_n409), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT32), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n636), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n530), .A2(KEYINPUT32), .A3(new_n531), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n545), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n626), .B1(new_n606), .B2(new_n612), .ZN(new_n694));
  INV_X1    g508(.A(new_n679), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n689), .A2(new_n693), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n687), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n289), .ZN(G30));
  NAND2_X1  g512(.A1(new_n613), .A2(new_n616), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n317), .B1(new_n270), .B2(new_n332), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n625), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT101), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n525), .A2(new_n516), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n468), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n706), .B(new_n262), .C1(new_n468), .C2(new_n540), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G472), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n704), .B1(new_n534), .B2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n691), .A2(new_n692), .A3(new_n704), .A4(new_n708), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NOR4_X1   g526(.A1(new_n701), .A2(new_n703), .A3(new_n695), .A4(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n686), .B(KEYINPUT39), .Z(new_n716));
  NOR2_X1   g530(.A1(new_n419), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT40), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n713), .A2(new_n714), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n285), .ZN(G45));
  NAND3_X1  g536(.A1(new_n648), .A2(new_n658), .A3(new_n686), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n696), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n222), .ZN(G48));
  NAND2_X1  g539(.A1(new_n693), .A2(new_n643), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n414), .B1(new_n413), .B2(new_n262), .ZN(new_n727));
  AOI211_X1 g541(.A(G469), .B(G902), .C1(new_n411), .C2(new_n412), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n727), .A2(new_n728), .A3(new_n335), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n660), .A2(new_n661), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT41), .B(G113), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NAND2_X1  g548(.A1(new_n606), .A2(new_n612), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n625), .A3(new_n729), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n726), .A2(new_n736), .A3(new_n624), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n670), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  NOR4_X1   g553(.A1(new_n727), .A2(new_n728), .A3(new_n624), .A4(new_n335), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n693), .A2(new_n694), .A3(new_n740), .A4(new_n695), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n333), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n422), .ZN(G21));
  INV_X1    g557(.A(new_n531), .ZN(new_n744));
  INV_X1    g558(.A(new_n631), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n542), .A2(new_n469), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n639), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n643), .A2(new_n729), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n624), .ZN(new_n751));
  INV_X1    g565(.A(new_n612), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n751), .B(new_n625), .C1(new_n752), .C2(new_n614), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n702), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G122), .ZN(G24));
  NOR3_X1   g570(.A1(new_n679), .A2(new_n639), .A3(new_n747), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n648), .A2(new_n658), .A3(new_n686), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n736), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n219), .ZN(G27));
  INV_X1    g574(.A(KEYINPUT103), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT42), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n626), .B1(new_n613), .B2(new_n616), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n546), .A2(new_n763), .A3(new_n689), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n762), .B1(new_n764), .B2(new_n723), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n761), .A2(KEYINPUT42), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n766), .B1(new_n764), .B2(new_n723), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  NAND2_X1  g585(.A1(new_n699), .A2(new_n625), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n419), .ZN(new_n773));
  INV_X1    g587(.A(new_n687), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT104), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n773), .A2(new_n774), .A3(new_n775), .A4(new_n546), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT104), .B1(new_n764), .B2(new_n687), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  AND2_X1   g593(.A1(new_n405), .A2(new_n408), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(KEYINPUT45), .ZN(new_n781));
  OAI21_X1  g595(.A(G469), .B1(new_n780), .B2(KEYINPUT45), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n416), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n728), .B1(new_n784), .B2(KEYINPUT46), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n785), .B1(KEYINPUT46), .B2(new_n784), .ZN(new_n786));
  INV_X1    g600(.A(new_n716), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(new_n336), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n326), .B1(new_n263), .B2(new_n264), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n789), .A2(new_n269), .B1(new_n331), .B2(new_n327), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n658), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT43), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n641), .A3(new_n695), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n772), .B(new_n788), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  NAND2_X1  g612(.A1(new_n786), .A2(new_n336), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT105), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n801), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n802), .B1(new_n799), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NOR4_X1   g620(.A1(new_n723), .A2(new_n772), .A3(new_n643), .A4(new_n693), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G140), .ZN(G42));
  NOR3_X1   g623(.A1(new_n772), .A2(new_n684), .A3(new_n730), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n643), .A3(new_n712), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n617), .B1(new_n812), .B2(new_n660), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n464), .A2(new_n639), .A3(new_n747), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n793), .A2(new_n618), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n793), .A2(new_n546), .A3(new_n810), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(KEYINPUT115), .B2(KEYINPUT48), .ZN(new_n817));
  NAND2_X1  g631(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n816), .A2(KEYINPUT115), .A3(KEYINPUT48), .ZN(new_n820));
  OAI221_X1 g634(.A(new_n813), .B1(new_n736), .B2(new_n815), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n727), .A2(new_n728), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n335), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n803), .B2(new_n805), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n701), .A2(new_n626), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n730), .A2(KEYINPUT50), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n824), .A2(new_n763), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n815), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n825), .A2(new_n729), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT50), .B1(new_n815), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n793), .A2(new_n757), .A3(new_n810), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n812), .A2(new_n790), .A3(new_n657), .A4(new_n656), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT114), .B1(new_n828), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n821), .B1(new_n834), .B2(KEYINPUT51), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n696), .B1(new_n723), .B2(new_n687), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n759), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT112), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n648), .A2(new_n735), .A3(new_n625), .A4(new_n666), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n336), .B(new_n686), .C1(new_n410), .C2(new_n418), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n691), .A2(new_n692), .A3(new_n708), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT101), .ZN(new_n844));
  AOI211_X1 g658(.A(new_n695), .B(new_n842), .C1(new_n844), .C2(new_n710), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n839), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n842), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n847), .B(new_n679), .C1(new_n709), .C2(new_n711), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n848), .A2(KEYINPUT112), .A3(new_n840), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n838), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT52), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n841), .A2(new_n845), .A3(new_n839), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT112), .B1(new_n848), .B2(new_n840), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n855), .A3(new_n838), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n789), .A2(new_n269), .B1(new_n331), .B2(new_n667), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT109), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT109), .B1(new_n313), .B2(new_n315), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n686), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n857), .A2(new_n763), .A3(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n863), .A2(KEYINPUT111), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n693), .A2(new_n689), .A3(new_n695), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n865), .B1(new_n863), .B2(KEYINPUT111), .ZN(new_n866));
  INV_X1    g680(.A(new_n773), .ZN(new_n867));
  OAI22_X1  g681(.A1(new_n864), .A2(new_n866), .B1(new_n758), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n851), .A2(new_n856), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n736), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n546), .A3(new_n751), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n546), .A2(new_n661), .A3(new_n729), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n872), .A2(new_n669), .B1(new_n873), .B2(new_n659), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n814), .A2(new_n661), .A3(new_n729), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n648), .A2(new_n666), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n875), .A2(new_n876), .B1(new_n333), .B2(new_n741), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT108), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n333), .ZN(new_n879));
  INV_X1    g693(.A(new_n741), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n879), .A2(new_n880), .B1(new_n702), .B2(new_n754), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT108), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n881), .A2(new_n732), .A3(new_n882), .A4(new_n738), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n768), .A2(new_n769), .B1(new_n776), .B2(new_n777), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT110), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n628), .A2(new_n790), .A3(new_n886), .A4(new_n860), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n860), .B(new_n332), .C1(new_n646), .C2(new_n647), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n613), .A2(new_n616), .A3(new_n627), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT110), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n887), .A2(new_n890), .A3(new_n645), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n645), .A2(new_n660), .A3(new_n628), .ZN(new_n892));
  AND4_X1   g706(.A1(new_n629), .A2(new_n891), .A3(new_n681), .A4(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n884), .A2(new_n885), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n836), .B1(new_n870), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n891), .A2(new_n629), .A3(new_n681), .A4(new_n892), .ZN(new_n897));
  NOR4_X1   g711(.A1(new_n897), .A2(new_n836), .A3(new_n874), .A4(new_n877), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n868), .B1(new_n850), .B2(KEYINPUT52), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n898), .A2(new_n899), .A3(new_n856), .A4(new_n885), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n895), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n897), .B1(new_n878), .B2(new_n883), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n899), .A2(new_n902), .A3(new_n856), .A4(new_n885), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT113), .B1(new_n903), .B2(new_n836), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n854), .A2(new_n855), .A3(new_n838), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n855), .B1(new_n854), .B2(new_n838), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n905), .A2(new_n906), .A3(new_n868), .ZN(new_n907));
  INV_X1    g721(.A(new_n894), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT113), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .A4(KEYINPUT53), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n904), .A2(new_n895), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n901), .B1(new_n911), .B2(KEYINPUT54), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n835), .B(new_n912), .C1(KEYINPUT51), .C2(new_n834), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(G952), .B2(G953), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n644), .A2(new_n626), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT106), .ZN(new_n916));
  INV_X1    g730(.A(new_n791), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n822), .B(KEYINPUT49), .Z(new_n918));
  NOR3_X1   g732(.A1(new_n918), .A2(new_n709), .A3(new_n711), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n916), .A2(new_n701), .A3(new_n917), .A4(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT107), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n914), .A2(new_n921), .ZN(G75));
  NOR2_X1   g736(.A1(new_n190), .A2(G952), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n895), .A2(new_n900), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(G210), .A3(G902), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n567), .A2(new_n582), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(new_n580), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(new_n583), .ZN(new_n928));
  XNOR2_X1  g742(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n928), .B(new_n929), .Z(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(KEYINPUT56), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n923), .B1(new_n925), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT117), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT56), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n924), .A2(KEYINPUT117), .A3(G210), .A4(G902), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT118), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n937), .A2(new_n938), .A3(new_n930), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n937), .B2(new_n930), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n932), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT119), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g757(.A(KEYINPUT119), .B(new_n932), .C1(new_n939), .C2(new_n940), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(G51));
  XNOR2_X1  g759(.A(new_n924), .B(KEYINPUT54), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n416), .B(KEYINPUT57), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n948), .A2(KEYINPUT120), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(KEYINPUT120), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n949), .A2(new_n413), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n924), .A2(G902), .A3(new_n783), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n923), .B1(new_n951), .B2(new_n952), .ZN(G54));
  AND4_X1   g767(.A1(KEYINPUT58), .A2(new_n924), .A3(G475), .A4(G902), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n954), .A2(new_n324), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(new_n324), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n955), .A2(new_n956), .A3(new_n923), .ZN(G60));
  INV_X1    g771(.A(new_n655), .ZN(new_n958));
  NAND2_X1  g772(.A1(G478), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT59), .Z(new_n960));
  NOR2_X1   g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n923), .B1(new_n946), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n960), .ZN(new_n963));
  NOR4_X1   g777(.A1(new_n870), .A2(new_n894), .A3(KEYINPUT113), .A4(new_n836), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT53), .B1(new_n907), .B2(new_n908), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n896), .B1(new_n966), .B2(new_n904), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n963), .B1(new_n967), .B2(new_n901), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT121), .B1(new_n968), .B2(new_n958), .ZN(new_n969));
  OAI211_X1 g783(.A(KEYINPUT121), .B(new_n958), .C1(new_n912), .C2(new_n960), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n962), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT122), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g788(.A(KEYINPUT122), .B(new_n962), .C1(new_n969), .C2(new_n971), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(G63));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT60), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n895), .B2(new_n900), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n923), .B1(new_n979), .B2(new_n676), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n455), .B2(new_n979), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g796(.A(new_n190), .B1(new_n619), .B2(G224), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT123), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n902), .A2(G953), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n983), .A2(new_n984), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n926), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(G898), .B2(new_n190), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT124), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n988), .B(new_n991), .ZN(G69));
  NOR2_X1   g806(.A1(new_n190), .A2(G900), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n788), .A2(new_n726), .A3(new_n840), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n994), .A2(new_n759), .A3(new_n837), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n797), .A2(new_n808), .A3(new_n885), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n993), .B1(new_n996), .B2(new_n190), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT125), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n523), .A2(new_n524), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(new_n319), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n997), .A2(new_n998), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n999), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n838), .B1(new_n719), .B2(new_n720), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT62), .Z(new_n1006));
  NAND2_X1  g820(.A1(new_n659), .A2(new_n888), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1007), .A2(new_n546), .A3(new_n717), .A4(new_n763), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1006), .A2(new_n797), .A3(new_n808), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n190), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n1001), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1004), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1012), .B1(new_n1004), .B2(new_n1011), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1014), .A2(new_n1015), .ZN(G72));
  XNOR2_X1  g830(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n638), .A2(new_n262), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n902), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1019), .B1(new_n996), .B2(new_n1020), .ZN(new_n1021));
  AOI211_X1 g835(.A(new_n468), .B(new_n705), .C1(new_n1021), .C2(KEYINPUT127), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1022), .B1(KEYINPUT127), .B2(new_n1021), .ZN(new_n1023));
  INV_X1    g837(.A(new_n526), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n911), .B(new_n1019), .C1(new_n1024), .C2(new_n536), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1019), .B1(new_n1009), .B2(new_n1020), .ZN(new_n1026));
  INV_X1    g840(.A(new_n706), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n923), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AND3_X1   g842(.A1(new_n1023), .A2(new_n1025), .A3(new_n1028), .ZN(G57));
endmodule


