//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT8), .Z(new_n190));
  OR2_X1    g004(.A1(KEYINPUT2), .A2(G113), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT2), .A2(G113), .ZN(new_n192));
  NAND2_X1  g006(.A1(G116), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(G116), .A2(G119), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n191), .B(new_n192), .C1(new_n194), .C2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT5), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n198), .B1(new_n194), .B2(new_n195), .ZN(new_n199));
  INV_X1    g013(.A(G116), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT66), .A3(new_n193), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n197), .B1(new_n199), .B2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n197), .A2(new_n201), .A3(G116), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT83), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n197), .A2(new_n201), .A3(KEYINPUT83), .A4(G116), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(G113), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n196), .B1(new_n204), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G107), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G104), .ZN(new_n214));
  OAI21_X1  g028(.A(G101), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT3), .B1(new_n211), .B2(G107), .ZN(new_n216));
  AOI21_X1  g030(.A(G101), .B1(new_n211), .B2(G107), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(new_n213), .A3(G104), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n210), .A2(new_n221), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n215), .A2(new_n220), .A3(new_n196), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT5), .B1(new_n194), .B2(new_n195), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n224), .A2(new_n207), .A3(G113), .A4(new_n208), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n190), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g042(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(G143), .B(G146), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(G128), .ZN(new_n232));
  INV_X1    g046(.A(G125), .ZN(new_n233));
  INV_X1    g047(.A(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G143), .ZN(new_n235));
  INV_X1    g049(.A(G143), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G146), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n241));
  INV_X1    g055(.A(new_n237), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n232), .A2(new_n233), .A3(new_n240), .A4(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n235), .A2(new_n237), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT0), .B(G128), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n231), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G125), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G953), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G224), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n252), .A2(KEYINPUT7), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n244), .A2(new_n249), .A3(new_n253), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT86), .B1(new_n227), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n190), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n215), .A2(new_n220), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n194), .A2(new_n195), .A3(new_n198), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT66), .B1(new_n202), .B2(new_n193), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT5), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n207), .A2(G113), .A3(new_n208), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n260), .B1(new_n265), .B2(new_n196), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n223), .A2(new_n225), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n259), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT86), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n244), .A2(new_n249), .A3(new_n253), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n253), .B1(new_n244), .B2(new_n249), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n268), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n265), .A2(new_n223), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n211), .A2(G107), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n216), .A2(new_n219), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G101), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n191), .A2(new_n192), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n199), .A2(new_n203), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n196), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT4), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n276), .A2(new_n282), .A3(G101), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n278), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n274), .A2(new_n284), .A3(new_n189), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n258), .A2(new_n273), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT87), .ZN(new_n287));
  INV_X1    g101(.A(G902), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n287), .B1(new_n286), .B2(new_n288), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n274), .A2(new_n284), .ZN(new_n292));
  INV_X1    g106(.A(new_n189), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT6), .A3(new_n285), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n252), .B(KEYINPUT84), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n250), .B(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT6), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n292), .A2(new_n298), .A3(new_n293), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n295), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n300), .B(KEYINPUT85), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n188), .B1(new_n291), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT88), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n210), .A2(new_n221), .B1(new_n223), .B2(new_n225), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n255), .B(new_n256), .C1(new_n304), .C2(new_n190), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n285), .B1(new_n305), .B2(KEYINPUT86), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n269), .B1(new_n268), .B2(new_n272), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n288), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT87), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT85), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n300), .B(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(new_n187), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n302), .A2(new_n303), .A3(new_n314), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n311), .A2(KEYINPUT88), .A3(new_n313), .A4(new_n187), .ZN(new_n316));
  INV_X1    g130(.A(G234), .ZN(new_n317));
  INV_X1    g131(.A(G237), .ZN(new_n318));
  OAI211_X1 g132(.A(G952), .B(new_n251), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(KEYINPUT95), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT68), .B(G953), .ZN(new_n322));
  AOI211_X1 g136(.A(new_n288), .B(new_n322), .C1(G234), .C2(G237), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT21), .B(G898), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G214), .B1(G237), .B2(G902), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n326), .B(KEYINPUT82), .Z(new_n327));
  NOR2_X1   g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n315), .A2(new_n316), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n322), .A2(G221), .A3(G234), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n330), .A2(KEYINPUT73), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT22), .B(G137), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(KEYINPUT73), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n332), .B1(new_n331), .B2(new_n333), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n201), .B2(G128), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n239), .A2(KEYINPUT23), .A3(G119), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n339), .B(new_n340), .C1(G119), .C2(new_n239), .ZN(new_n341));
  XNOR2_X1  g155(.A(G119), .B(G128), .ZN(new_n342));
  XOR2_X1   g156(.A(KEYINPUT24), .B(G110), .Z(new_n343));
  AOI22_X1  g157(.A1(new_n341), .A2(G110), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G125), .B(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT16), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT16), .ZN(new_n347));
  INV_X1    g161(.A(G140), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(G125), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(G146), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(G146), .B1(new_n346), .B2(new_n349), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n344), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n354));
  OAI22_X1  g168(.A1(new_n341), .A2(G110), .B1(new_n342), .B2(new_n343), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n345), .A2(new_n234), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n350), .A3(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n353), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n354), .B1(new_n353), .B2(new_n357), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n337), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n336), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n334), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n353), .A2(new_n357), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n362), .B1(KEYINPUT74), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(G217), .B1(new_n317), .B2(G902), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n288), .ZN(new_n366));
  XOR2_X1   g180(.A(new_n366), .B(KEYINPUT75), .Z(new_n367));
  NAND3_X1  g181(.A1(new_n360), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT76), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n360), .A2(new_n364), .A3(KEYINPUT76), .A4(new_n367), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT25), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n360), .A2(new_n364), .A3(new_n373), .A4(new_n288), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n360), .A2(new_n288), .A3(new_n364), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n365), .B1(new_n375), .B2(KEYINPUT25), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n372), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT67), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n248), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT11), .ZN(new_n381));
  INV_X1    g195(.A(G134), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n381), .B1(new_n382), .B2(G137), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(G137), .ZN(new_n384));
  INV_X1    g198(.A(G137), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(KEYINPUT11), .A3(G134), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G131), .ZN(new_n388));
  INV_X1    g202(.A(G131), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n383), .A2(new_n386), .A3(new_n389), .A4(new_n384), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n246), .B(KEYINPUT67), .C1(new_n231), .C2(new_n247), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n380), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n232), .A2(new_n240), .A3(new_n243), .ZN(new_n394));
  INV_X1    g208(.A(new_n384), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n382), .A2(G137), .ZN(new_n396));
  OAI21_X1  g210(.A(G131), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n390), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n281), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n393), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT28), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT70), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n393), .A2(new_n398), .A3(KEYINPUT70), .A4(new_n399), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n393), .A2(new_n398), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n281), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT71), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT71), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n411), .A3(new_n281), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n407), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n403), .B1(new_n413), .B2(KEYINPUT28), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT26), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n251), .A2(KEYINPUT68), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT68), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G953), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n416), .A2(new_n418), .A3(G210), .A4(new_n318), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT27), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT27), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n322), .A2(new_n421), .A3(G210), .A4(new_n318), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n415), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n420), .A2(new_n422), .A3(new_n415), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(G101), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G101), .ZN(new_n427));
  INV_X1    g241(.A(new_n425), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n427), .B1(new_n428), .B2(new_n423), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT29), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(G902), .B1(new_n414), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT64), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n248), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n246), .B(KEYINPUT64), .C1(new_n231), .C2(new_n247), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n391), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n398), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n400), .A2(new_n401), .B1(new_n438), .B2(new_n281), .ZN(new_n439));
  INV_X1    g253(.A(new_n430), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n393), .A2(new_n398), .A3(KEYINPUT28), .A4(new_n399), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n393), .A2(KEYINPUT30), .A3(new_n398), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT30), .B1(new_n437), .B2(new_n398), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n444), .A2(new_n445), .A3(new_n399), .ZN(new_n446));
  INV_X1    g260(.A(new_n400), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n430), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT69), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n443), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n431), .B1(new_n442), .B2(KEYINPUT69), .ZN(new_n451));
  OAI22_X1  g265(.A1(new_n433), .A2(KEYINPUT72), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n413), .A2(KEYINPUT28), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n402), .A3(new_n432), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n288), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT72), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G472), .B1(new_n452), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n439), .A2(new_n441), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n430), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT30), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n438), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n393), .A2(new_n398), .A3(KEYINPUT30), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n281), .A3(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n400), .A2(new_n426), .A3(new_n429), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n464), .A2(KEYINPUT31), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT31), .B1(new_n464), .B2(new_n465), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(G472), .A2(G902), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT32), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT32), .B1(new_n468), .B2(new_n469), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n378), .B1(new_n458), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT9), .B(G234), .ZN(new_n476));
  OAI21_X1  g290(.A(G221), .B1(new_n476), .B2(G902), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT81), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n322), .A2(G227), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(G140), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT77), .B(G110), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n278), .A2(new_n380), .A3(new_n392), .A4(new_n283), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n388), .A2(new_n390), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n236), .A2(KEYINPUT1), .A3(G146), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n238), .B2(new_n239), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n232), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT10), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n489), .A2(new_n260), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n490), .B1(new_n394), .B2(new_n260), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n485), .B(new_n486), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT78), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n260), .A3(new_n490), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n239), .A2(new_n238), .B1(new_n241), .B2(new_n242), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n221), .B1(new_n232), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n496), .B1(new_n498), .B2(new_n490), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n499), .A2(KEYINPUT78), .A3(new_n486), .A4(new_n485), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n394), .A2(new_n260), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n221), .B1(new_n232), .B2(new_n488), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n391), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT79), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT12), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n489), .A2(new_n260), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n497), .A2(new_n221), .A3(new_n232), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n486), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT79), .B1(new_n510), .B2(KEYINPUT12), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(KEYINPUT12), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n507), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n501), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT80), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT80), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n501), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n484), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n483), .B1(new_n495), .B2(new_n500), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n499), .A2(new_n485), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n391), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n479), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n517), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n516), .B1(new_n501), .B2(new_n513), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n483), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(KEYINPUT81), .A3(new_n522), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n528), .A3(G469), .ZN(new_n529));
  INV_X1    g343(.A(G469), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n519), .A2(new_n513), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n484), .B1(new_n501), .B2(new_n521), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n530), .B(new_n288), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(G469), .A2(G902), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n478), .B1(new_n529), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n416), .A2(new_n418), .A3(G214), .A4(new_n318), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n236), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n322), .A2(G143), .A3(G214), .A4(new_n318), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G131), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT89), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT89), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n540), .A2(new_n544), .A3(G131), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n538), .A2(new_n539), .A3(new_n389), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n542), .A2(new_n543), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n351), .A2(new_n352), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n544), .B1(new_n540), .B2(G131), .ZN(new_n549));
  AOI211_X1 g363(.A(KEYINPUT89), .B(new_n389), .C1(new_n538), .C2(new_n539), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT17), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n547), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G113), .B(G122), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(new_n211), .ZN(new_n554));
  AND2_X1   g368(.A1(KEYINPUT18), .A2(G131), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n540), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n348), .A2(G125), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n233), .A2(G140), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(G146), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n356), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n540), .B2(new_n555), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n552), .A2(new_n554), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n554), .B1(new_n552), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n288), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G475), .ZN(new_n568));
  NOR2_X1   g382(.A1(G475), .A2(G902), .ZN(new_n569));
  XOR2_X1   g383(.A(new_n569), .B(KEYINPUT91), .Z(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n552), .A2(new_n554), .A3(new_n564), .ZN(new_n572));
  INV_X1    g386(.A(new_n554), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n345), .B(KEYINPUT19), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT90), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n234), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n345), .A2(KEYINPUT19), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n234), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT90), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n576), .A2(new_n580), .A3(new_n350), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n549), .A2(new_n550), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(new_n546), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n573), .B1(new_n583), .B2(new_n563), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n571), .B1(new_n572), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n572), .A2(new_n584), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT92), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT20), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT92), .ZN(new_n590));
  AND4_X1   g404(.A1(new_n590), .A2(new_n586), .A3(new_n588), .A4(new_n570), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n568), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G478), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(KEYINPUT15), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT93), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n200), .A2(G122), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n595), .B1(new_n596), .B2(KEYINPUT14), .ZN(new_n597));
  INV_X1    g411(.A(G122), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G116), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT14), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n600), .A2(new_n200), .A3(KEYINPUT93), .A4(G122), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n596), .A2(KEYINPUT14), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n597), .A2(new_n599), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(G107), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n599), .A2(new_n596), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n213), .ZN(new_n606));
  XNOR2_X1  g420(.A(G128), .B(G143), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(G134), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n382), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n604), .B(new_n606), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n605), .B(new_n213), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT13), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n236), .A3(G128), .ZN(new_n614));
  OAI211_X1 g428(.A(G134), .B(new_n614), .C1(new_n608), .C2(new_n613), .ZN(new_n615));
  INV_X1    g429(.A(new_n609), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n612), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(G217), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n476), .A2(new_n619), .A3(G953), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n611), .A2(new_n617), .A3(new_n620), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT94), .B1(new_n624), .B2(new_n288), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT94), .ZN(new_n626));
  AOI211_X1 g440(.A(new_n626), .B(G902), .C1(new_n622), .C2(new_n623), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n594), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n624), .B(new_n288), .C1(KEYINPUT15), .C2(new_n593), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n592), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n329), .A2(new_n475), .A3(new_n536), .A4(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  AOI21_X1  g447(.A(new_n440), .B1(new_n439), .B2(new_n441), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT31), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n400), .A2(new_n426), .A3(new_n429), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n635), .B1(new_n446), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT31), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n634), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(G472), .B1(new_n639), .B2(G902), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n377), .A2(new_n470), .A3(new_n640), .ZN(new_n641));
  AOI211_X1 g455(.A(new_n478), .B(new_n641), .C1(new_n529), .C2(new_n535), .ZN(new_n642));
  INV_X1    g456(.A(new_n327), .ZN(new_n643));
  INV_X1    g457(.A(new_n325), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n291), .A2(new_n301), .A3(new_n188), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n187), .B1(new_n311), .B2(new_n313), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n643), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  OR2_X1    g461(.A1(new_n625), .A2(new_n627), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n624), .B(KEYINPUT33), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n593), .A2(G902), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n648), .A2(new_n593), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n592), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n642), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT34), .B(G104), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  NAND2_X1  g471(.A1(new_n302), .A2(new_n314), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n585), .A2(new_n588), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n585), .A2(new_n588), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n630), .B(new_n568), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n658), .A2(new_n643), .A3(new_n662), .A4(new_n644), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n642), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NAND2_X1  g480(.A1(new_n376), .A2(new_n374), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n362), .A2(KEYINPUT36), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n363), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n367), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n640), .A2(new_n470), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n329), .A2(new_n536), .A3(new_n631), .A4(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n323), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(KEYINPUT96), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(KEYINPUT96), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n321), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n661), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n536), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n327), .B1(new_n302), .B2(new_n314), .ZN(new_n685));
  INV_X1    g499(.A(G472), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n448), .A2(new_n449), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n451), .B1(new_n687), .B2(new_n442), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n455), .B2(new_n456), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n686), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n472), .ZN(new_n692));
  INV_X1    g506(.A(new_n469), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n471), .B1(new_n639), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n685), .B(new_n671), .C1(new_n691), .C2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n684), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n239), .ZN(G30));
  INV_X1    g512(.A(KEYINPUT99), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n682), .B(KEYINPUT39), .Z(new_n700));
  AND2_X1   g514(.A1(new_n536), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n699), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(KEYINPUT99), .A3(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT98), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n464), .A2(new_n400), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n440), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n710), .B(new_n288), .C1(new_n440), .C2(new_n413), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G472), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT97), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n474), .ZN(new_n714));
  INV_X1    g528(.A(new_n586), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n590), .B1(new_n572), .B2(new_n584), .ZN(new_n716));
  OAI22_X1  g530(.A1(new_n715), .A2(new_n571), .B1(new_n716), .B2(KEYINPUT20), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n587), .A2(new_n588), .A3(new_n585), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n717), .A2(new_n718), .B1(G475), .B2(new_n567), .ZN(new_n719));
  INV_X1    g533(.A(new_n630), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AND4_X1   g535(.A1(new_n643), .A2(new_n714), .A3(new_n672), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n315), .A2(new_n316), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT38), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n315), .A2(KEYINPUT38), .A3(new_n316), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n708), .B1(new_n722), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n722), .A2(new_n727), .A3(new_n708), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n704), .B(new_n707), .C1(new_n728), .C2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G143), .ZN(G45));
  NAND2_X1  g546(.A1(new_n529), .A2(new_n535), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n719), .A2(new_n651), .A3(new_n682), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n477), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n696), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n234), .ZN(G48));
  NAND2_X1  g551(.A1(new_n501), .A2(new_n521), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n738), .A2(new_n483), .B1(new_n519), .B2(new_n513), .ZN(new_n739));
  OAI21_X1  g553(.A(G469), .B1(new_n739), .B2(G902), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n477), .A3(new_n533), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT100), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT100), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n740), .A2(new_n743), .A3(new_n533), .A4(new_n477), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n742), .A2(KEYINPUT101), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT101), .B1(new_n742), .B2(new_n744), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n654), .B(new_n475), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT102), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n742), .A2(new_n744), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT101), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n742), .A2(KEYINPUT101), .A3(new_n744), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(KEYINPUT102), .A3(new_n475), .A4(new_n654), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n749), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g570(.A(KEYINPUT41), .B(G113), .Z(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT103), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n756), .B(new_n758), .ZN(G15));
  OAI211_X1 g573(.A(new_n663), .B(new_n475), .C1(new_n745), .C2(new_n746), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G116), .ZN(G18));
  AOI21_X1  g575(.A(new_n672), .B1(new_n458), .B2(new_n474), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n742), .A2(new_n744), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n592), .A2(new_n325), .A3(new_n630), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n762), .A2(new_n763), .A3(new_n685), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G119), .ZN(G21));
  NAND2_X1  g580(.A1(new_n468), .A2(new_n288), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n637), .A2(new_n638), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n414), .B2(new_n440), .ZN(new_n769));
  AOI22_X1  g583(.A1(G472), .A2(new_n767), .B1(new_n769), .B2(new_n469), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(new_n377), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n644), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n752), .B2(new_n753), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT104), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n721), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT104), .B1(new_n719), .B2(new_n720), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n685), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G122), .ZN(G24));
  INV_X1    g594(.A(KEYINPUT105), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n781), .B1(new_n770), .B2(new_n671), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n769), .A2(new_n469), .ZN(new_n783));
  AND4_X1   g597(.A1(new_n781), .A2(new_n783), .A3(new_n671), .A4(new_n640), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n734), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n685), .A2(new_n744), .A3(new_n742), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT106), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n685), .A2(new_n744), .A3(new_n742), .ZN(new_n788));
  INV_X1    g602(.A(new_n682), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n592), .A2(new_n652), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n783), .A2(new_n671), .A3(new_n640), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT105), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n770), .A2(new_n781), .A3(new_n671), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT106), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n788), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n787), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G125), .ZN(G27));
  AOI21_X1  g612(.A(new_n327), .B1(new_n315), .B2(new_n316), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT42), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n790), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n533), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n534), .B(KEYINPUT107), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n527), .A2(G469), .A3(new_n522), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n478), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n799), .A2(new_n801), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n473), .A2(KEYINPUT108), .A3(KEYINPUT109), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT108), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n810), .B1(new_n694), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n692), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT109), .B1(new_n473), .B2(KEYINPUT108), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n694), .A2(new_n811), .A3(new_n810), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n472), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n813), .A2(new_n458), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT110), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n817), .A2(new_n818), .A3(new_n377), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n818), .B1(new_n817), .B2(new_n377), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n808), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n475), .A2(new_n799), .A3(new_n734), .A4(new_n806), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n800), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G131), .ZN(G33));
  NAND4_X1  g639(.A1(new_n475), .A2(new_n799), .A3(new_n683), .A4(new_n806), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G134), .ZN(G36));
  OAI21_X1  g641(.A(KEYINPUT43), .B1(new_n592), .B2(new_n651), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT43), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n719), .A2(new_n829), .A3(new_n652), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n673), .A2(new_n671), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(KEYINPUT44), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n799), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT112), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT45), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n518), .A2(new_n479), .A3(new_n523), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT81), .B1(new_n527), .B2(new_n522), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n527), .A2(KEYINPUT45), .A3(new_n522), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(G469), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n803), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT111), .B1(new_n843), .B2(KEYINPUT46), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n802), .B1(new_n843), .B2(KEYINPUT46), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT111), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT46), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n524), .A2(new_n528), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n841), .B1(new_n848), .B2(new_n836), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n846), .B(new_n847), .C1(new_n849), .C2(new_n803), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n844), .A2(new_n845), .A3(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n851), .A2(new_n477), .A3(new_n700), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n831), .A2(new_n832), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n835), .B(new_n852), .C1(KEYINPUT44), .C2(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(G137), .ZN(G39));
  NAND2_X1  g669(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n851), .A2(new_n477), .A3(new_n856), .ZN(new_n857));
  XOR2_X1   g671(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n851), .B2(new_n477), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n691), .A2(new_n790), .A3(new_n695), .A4(new_n377), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n799), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(G140), .ZN(G42));
  INV_X1    g677(.A(new_n727), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n714), .A2(new_n378), .A3(new_n327), .A4(new_n478), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n592), .A2(new_n651), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n740), .A2(new_n533), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT49), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n864), .A2(new_n865), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n632), .A2(new_n765), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n760), .A2(new_n675), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n641), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n733), .A2(new_n477), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n315), .A2(new_n316), .A3(new_n328), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT114), .B1(new_n719), .B2(new_n651), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT114), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n592), .A2(new_n880), .A3(new_n652), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n879), .B(new_n881), .C1(new_n592), .C2(new_n720), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n778), .A2(new_n773), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n756), .A2(new_n872), .A3(new_n874), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n630), .A2(new_n682), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n885), .B(new_n568), .C1(new_n660), .C2(new_n659), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n762), .A2(new_n799), .A3(new_n536), .A4(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n794), .A2(new_n799), .A3(new_n806), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n826), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n817), .A2(new_n377), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT110), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n817), .A2(new_n818), .A3(new_n377), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n807), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n823), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n891), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n884), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n696), .B1(new_n684), .B2(new_n735), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n714), .A2(new_n806), .A3(new_n672), .A4(new_n789), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n777), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n797), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT52), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n899), .B1(new_n796), .B2(new_n787), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(KEYINPUT52), .A3(new_n902), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n898), .A2(KEYINPUT115), .A3(KEYINPUT53), .A4(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT52), .B1(new_n906), .B2(new_n902), .ZN(new_n911));
  AND4_X1   g725(.A1(KEYINPUT52), .A2(new_n900), .A3(new_n797), .A4(new_n902), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n890), .B1(new_n821), .B2(new_n823), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n642), .A2(new_n882), .A3(new_n329), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n644), .B(new_n771), .C1(new_n745), .C2(new_n746), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(new_n777), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n917), .A2(new_n873), .A3(new_n871), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n914), .A2(new_n918), .A3(new_n756), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n910), .B1(new_n913), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n909), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n884), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n908), .A2(new_n922), .A3(KEYINPUT53), .A4(new_n914), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT115), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n870), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n920), .A2(KEYINPUT116), .A3(new_n923), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT116), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n928), .B(new_n910), .C1(new_n913), .C2(new_n919), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT54), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n831), .A2(new_n321), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n792), .A2(new_n793), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n799), .A2(new_n763), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n799), .B2(new_n763), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n931), .B(new_n932), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n714), .A2(new_n378), .A3(new_n320), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n592), .A2(new_n652), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n937), .B(new_n938), .C1(new_n934), .C2(new_n935), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n315), .A2(KEYINPUT38), .A3(new_n316), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT38), .B1(new_n315), .B2(new_n316), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n742), .A2(new_n327), .A3(new_n744), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n771), .A2(new_n828), .A3(new_n830), .A4(new_n321), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n942), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n742), .A2(new_n327), .A3(new_n744), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n725), .A2(new_n726), .A3(new_n950), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n951), .A2(new_n941), .A3(new_n947), .ZN(new_n952));
  OAI21_X1  g766(.A(KEYINPUT119), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n946), .A2(new_n942), .A3(new_n948), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n941), .B1(new_n951), .B2(new_n947), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT119), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n940), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(KEYINPUT121), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT121), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n940), .A2(new_n953), .A3(new_n960), .A4(new_n957), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n867), .A2(new_n478), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n857), .B2(new_n859), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n948), .A2(new_n799), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT117), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n959), .A2(new_n961), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT51), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(G952), .ZN(new_n970));
  AOI211_X1 g784(.A(new_n970), .B(G953), .C1(new_n948), .C2(new_n788), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n937), .B1(new_n934), .B2(new_n935), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n831), .A2(new_n321), .ZN(new_n973));
  INV_X1    g787(.A(new_n935), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n799), .A2(new_n763), .A3(new_n933), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n893), .A2(new_n894), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT48), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n976), .B2(new_n977), .ZN(new_n980));
  OAI221_X1 g794(.A(new_n971), .B1(new_n653), .B2(new_n972), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n968), .B1(new_n954), .B2(new_n955), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n940), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n981), .B1(new_n966), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n969), .A2(new_n984), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n926), .A2(new_n930), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n970), .A2(new_n251), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT122), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n869), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(KEYINPUT123), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT123), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n991), .B(new_n869), .C1(new_n986), .C2(new_n988), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(G75));
  NAND2_X1  g807(.A1(new_n927), .A2(new_n929), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n994), .A2(new_n288), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(G210), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT56), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n295), .A2(new_n299), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(new_n297), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT55), .Z(new_n1000));
  AND3_X1   g814(.A1(new_n996), .A2(new_n997), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1000), .B1(new_n996), .B2(new_n997), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n322), .A2(G952), .ZN(new_n1003));
  NOR3_X1   g817(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(G51));
  XNOR2_X1  g818(.A(new_n803), .B(KEYINPUT57), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n994), .A2(new_n870), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1005), .B1(new_n1006), .B2(new_n930), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1007), .B1(new_n532), .B2(new_n531), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n995), .A2(new_n849), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1003), .B1(new_n1008), .B2(new_n1009), .ZN(G54));
  NAND3_X1  g824(.A1(new_n995), .A2(KEYINPUT58), .A3(G475), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n1011), .A2(new_n715), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1011), .A2(new_n715), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1012), .A2(new_n1013), .A3(new_n1003), .ZN(G60));
  OR2_X1    g828(.A1(new_n926), .A2(new_n930), .ZN(new_n1015));
  NAND2_X1  g829(.A1(G478), .A2(G902), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT59), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n649), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n649), .B(new_n1017), .C1(new_n1006), .C2(new_n930), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1003), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1018), .A2(new_n1021), .ZN(G63));
  NAND2_X1  g836(.A1(new_n360), .A2(new_n364), .ZN(new_n1023));
  NAND2_X1  g837(.A1(G217), .A2(G902), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(KEYINPUT60), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1023), .B1(new_n994), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1025), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n927), .A2(new_n669), .A3(new_n929), .A4(new_n1027), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1026), .A2(new_n1020), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(KEYINPUT61), .B1(new_n1028), .B2(KEYINPUT124), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1029), .B(new_n1030), .ZN(G66));
  INV_X1    g845(.A(G224), .ZN(new_n1032));
  OAI21_X1  g846(.A(G953), .B1(new_n324), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(new_n322), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1033), .B1(new_n922), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g849(.A(G898), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n998), .B1(new_n1036), .B2(new_n1034), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1035), .B(new_n1037), .Z(G69));
  AOI21_X1  g852(.A(new_n322), .B1(G227), .B2(G900), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n701), .A2(new_n475), .A3(new_n799), .A4(new_n882), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g855(.A(KEYINPUT62), .B1(new_n731), .B2(new_n906), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n731), .A2(KEYINPUT62), .A3(new_n906), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n862), .A2(new_n854), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1034), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n444), .A2(new_n445), .ZN(new_n1049));
  XNOR2_X1  g863(.A(new_n1049), .B(new_n574), .ZN(new_n1050));
  XNOR2_X1  g864(.A(new_n1050), .B(KEYINPUT125), .ZN(new_n1051));
  OAI21_X1  g865(.A(KEYINPUT126), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g866(.A(new_n1044), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1040), .B1(new_n1053), .B2(new_n1042), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n322), .B1(new_n1054), .B2(new_n1046), .ZN(new_n1055));
  INV_X1    g869(.A(KEYINPUT126), .ZN(new_n1056));
  INV_X1    g870(.A(new_n1051), .ZN(new_n1057));
  NAND3_X1  g871(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1052), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1034), .A2(G900), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n852), .A2(new_n778), .A3(new_n977), .ZN(new_n1061));
  AND3_X1   g875(.A1(new_n824), .A2(new_n826), .A3(new_n906), .ZN(new_n1062));
  NAND4_X1  g876(.A1(new_n862), .A2(new_n854), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  OAI211_X1 g877(.A(new_n1050), .B(new_n1060), .C1(new_n1063), .C2(new_n1034), .ZN(new_n1064));
  INV_X1    g878(.A(KEYINPUT127), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g880(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n1039), .B1(new_n1059), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g882(.A(new_n1039), .ZN(new_n1069));
  AOI211_X1 g883(.A(new_n1069), .B(new_n1066), .C1(new_n1052), .C2(new_n1058), .ZN(new_n1070));
  NOR2_X1   g884(.A1(new_n1068), .A2(new_n1070), .ZN(G72));
  NAND2_X1  g885(.A1(G472), .A2(G902), .ZN(new_n1072));
  XOR2_X1   g886(.A(new_n1072), .B(KEYINPUT63), .Z(new_n1073));
  OAI21_X1  g887(.A(new_n1073), .B1(new_n1063), .B2(new_n884), .ZN(new_n1074));
  NOR2_X1   g888(.A1(new_n709), .A2(new_n440), .ZN(new_n1075));
  NAND2_X1  g889(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g890(.A1(new_n1076), .A2(new_n1020), .ZN(new_n1077));
  NAND3_X1  g891(.A1(new_n1045), .A2(new_n1047), .A3(new_n922), .ZN(new_n1078));
  AOI21_X1  g892(.A(new_n710), .B1(new_n1078), .B2(new_n1073), .ZN(new_n1079));
  NAND2_X1  g893(.A1(new_n921), .A2(new_n925), .ZN(new_n1080));
  NAND2_X1  g894(.A1(new_n710), .A2(new_n1073), .ZN(new_n1081));
  NOR2_X1   g895(.A1(new_n1081), .A2(new_n1075), .ZN(new_n1082));
  AOI211_X1 g896(.A(new_n1077), .B(new_n1079), .C1(new_n1080), .C2(new_n1082), .ZN(G57));
endmodule


