

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592;

  INV_X1 U325 ( .A(KEYINPUT101), .ZN(n472) );
  XNOR2_X1 U326 ( .A(n438), .B(n437), .ZN(n439) );
  NAND2_X1 U327 ( .A1(n481), .A2(n480), .ZN(n491) );
  NAND2_X1 U328 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U329 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U330 ( .A(n442), .B(n441), .ZN(n562) );
  NAND2_X1 U331 ( .A1(n532), .A2(n541), .ZN(n293) );
  XOR2_X1 U332 ( .A(n347), .B(n346), .Z(n294) );
  NOR2_X1 U333 ( .A1(n369), .A2(n576), .ZN(n370) );
  XNOR2_X1 U334 ( .A(n430), .B(n339), .ZN(n340) );
  XOR2_X1 U335 ( .A(G148GAT), .B(G78GAT), .Z(n430) );
  XNOR2_X1 U336 ( .A(n341), .B(n340), .ZN(n343) );
  XNOR2_X1 U337 ( .A(n547), .B(n472), .ZN(n473) );
  XNOR2_X1 U338 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n309) );
  XNOR2_X1 U339 ( .A(n428), .B(n427), .ZN(n434) );
  XNOR2_X1 U340 ( .A(n309), .B(KEYINPUT74), .ZN(n338) );
  XNOR2_X1 U341 ( .A(n495), .B(KEYINPUT37), .ZN(n496) );
  XNOR2_X1 U342 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U343 ( .A(n330), .B(n329), .ZN(n332) );
  XNOR2_X1 U344 ( .A(n497), .B(n496), .ZN(n521) );
  XNOR2_X1 U345 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n441) );
  XNOR2_X1 U346 ( .A(n440), .B(n439), .ZN(n476) );
  INV_X1 U347 ( .A(G190GAT), .ZN(n461) );
  XNOR2_X1 U348 ( .A(n499), .B(KEYINPUT38), .ZN(n508) );
  XNOR2_X1 U349 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U350 ( .A(n464), .B(n463), .ZN(G1351GAT) );
  INV_X1 U351 ( .A(KEYINPUT64), .ZN(n420) );
  XOR2_X1 U352 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n296) );
  XNOR2_X1 U353 ( .A(KEYINPUT84), .B(KEYINPUT12), .ZN(n295) );
  XNOR2_X1 U354 ( .A(n296), .B(n295), .ZN(n308) );
  XOR2_X1 U355 ( .A(G211GAT), .B(G155GAT), .Z(n298) );
  XNOR2_X1 U356 ( .A(G8GAT), .B(G127GAT), .ZN(n297) );
  XNOR2_X1 U357 ( .A(n298), .B(n297), .ZN(n306) );
  XOR2_X1 U358 ( .A(G78GAT), .B(KEYINPUT81), .Z(n300) );
  XNOR2_X1 U359 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n299) );
  XNOR2_X1 U360 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U361 ( .A(G64GAT), .B(G71GAT), .Z(n302) );
  XNOR2_X1 U362 ( .A(G22GAT), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U363 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U364 ( .A(n304), .B(n303), .Z(n305) );
  XNOR2_X1 U365 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n313) );
  XOR2_X1 U367 ( .A(G1GAT), .B(G15GAT), .Z(n354) );
  XOR2_X1 U368 ( .A(n338), .B(n354), .Z(n311) );
  NAND2_X1 U369 ( .A1(G231GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n313), .B(n312), .ZN(n570) );
  XNOR2_X1 U372 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n314) );
  XNOR2_X1 U373 ( .A(n314), .B(G29GAT), .ZN(n315) );
  XOR2_X1 U374 ( .A(n315), .B(KEYINPUT8), .Z(n317) );
  XNOR2_X1 U375 ( .A(G43GAT), .B(G50GAT), .ZN(n316) );
  XNOR2_X1 U376 ( .A(n317), .B(n316), .ZN(n367) );
  XOR2_X1 U377 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n319) );
  XNOR2_X1 U378 ( .A(KEYINPUT79), .B(KEYINPUT67), .ZN(n318) );
  XNOR2_X1 U379 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n367), .B(n320), .ZN(n334) );
  XOR2_X1 U381 ( .A(G162GAT), .B(G218GAT), .Z(n429) );
  XNOR2_X1 U382 ( .A(G106GAT), .B(G92GAT), .ZN(n322) );
  XNOR2_X1 U383 ( .A(G99GAT), .B(G85GAT), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n322), .B(n321), .ZN(n323) );
  INV_X1 U385 ( .A(n323), .ZN(n350) );
  NAND2_X1 U386 ( .A1(n429), .A2(n350), .ZN(n326) );
  INV_X1 U387 ( .A(n429), .ZN(n324) );
  NAND2_X1 U388 ( .A1(n324), .A2(n323), .ZN(n325) );
  NAND2_X1 U389 ( .A1(n326), .A2(n325), .ZN(n330) );
  AND2_X1 U390 ( .A1(G232GAT), .A2(G233GAT), .ZN(n328) );
  INV_X1 U391 ( .A(KEYINPUT9), .ZN(n327) );
  XOR2_X1 U392 ( .A(G190GAT), .B(G134GAT), .Z(n453) );
  XNOR2_X1 U393 ( .A(n453), .B(KEYINPUT10), .ZN(n331) );
  XNOR2_X1 U394 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n334), .B(n333), .ZN(n559) );
  XOR2_X1 U396 ( .A(KEYINPUT80), .B(n559), .Z(n541) );
  XOR2_X1 U397 ( .A(KEYINPUT36), .B(KEYINPUT105), .Z(n335) );
  XNOR2_X1 U398 ( .A(n541), .B(n335), .ZN(n493) );
  NAND2_X1 U399 ( .A1(n570), .A2(n493), .ZN(n336) );
  XNOR2_X1 U400 ( .A(n336), .B(KEYINPUT45), .ZN(n337) );
  XNOR2_X1 U401 ( .A(KEYINPUT65), .B(n337), .ZN(n352) );
  XOR2_X1 U402 ( .A(G120GAT), .B(G71GAT), .Z(n454) );
  XOR2_X1 U403 ( .A(n338), .B(n454), .Z(n341) );
  NAND2_X1 U404 ( .A1(G230GAT), .A2(G233GAT), .ZN(n339) );
  XOR2_X1 U405 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U407 ( .A(KEYINPUT76), .B(KEYINPUT33), .Z(n345) );
  XNOR2_X1 U408 ( .A(KEYINPUT75), .B(KEYINPUT77), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U410 ( .A(G64GAT), .B(G204GAT), .Z(n349) );
  XNOR2_X1 U411 ( .A(G176GAT), .B(KEYINPUT78), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n381) );
  XNOR2_X1 U413 ( .A(n350), .B(n381), .ZN(n351) );
  XOR2_X1 U414 ( .A(n294), .B(n351), .Z(n582) );
  NAND2_X1 U415 ( .A1(n352), .A2(n582), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n353), .B(KEYINPUT115), .ZN(n368) );
  XOR2_X1 U417 ( .A(G141GAT), .B(G22GAT), .Z(n427) );
  XOR2_X1 U418 ( .A(n427), .B(n354), .Z(n356) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U420 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U421 ( .A(G169GAT), .B(G8GAT), .Z(n391) );
  XOR2_X1 U422 ( .A(n357), .B(n391), .Z(n365) );
  XOR2_X1 U423 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n359) );
  XNOR2_X1 U424 ( .A(G113GAT), .B(G197GAT), .ZN(n358) );
  XNOR2_X1 U425 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U426 ( .A(KEYINPUT72), .B(KEYINPUT69), .Z(n361) );
  XNOR2_X1 U427 ( .A(KEYINPUT71), .B(KEYINPUT30), .ZN(n360) );
  XNOR2_X1 U428 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n576) );
  XOR2_X1 U432 ( .A(KEYINPUT73), .B(n576), .Z(n465) );
  NAND2_X1 U433 ( .A1(n368), .A2(n465), .ZN(n376) );
  XNOR2_X1 U434 ( .A(n582), .B(KEYINPUT41), .ZN(n510) );
  INV_X1 U435 ( .A(n510), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(KEYINPUT46), .ZN(n371) );
  NOR2_X1 U437 ( .A1(n570), .A2(n371), .ZN(n372) );
  NAND2_X1 U438 ( .A1(n372), .A2(n559), .ZN(n374) );
  XOR2_X1 U439 ( .A(KEYINPUT114), .B(KEYINPUT47), .Z(n373) );
  XNOR2_X1 U440 ( .A(n374), .B(n373), .ZN(n375) );
  NAND2_X1 U441 ( .A1(n376), .A2(n375), .ZN(n378) );
  INV_X1 U442 ( .A(KEYINPUT48), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n548) );
  XOR2_X1 U444 ( .A(G183GAT), .B(KEYINPUT17), .Z(n380) );
  XNOR2_X1 U445 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n379) );
  XNOR2_X1 U446 ( .A(n380), .B(n379), .ZN(n449) );
  XNOR2_X1 U447 ( .A(n449), .B(n381), .ZN(n389) );
  XOR2_X1 U448 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n387) );
  XOR2_X1 U449 ( .A(G92GAT), .B(G218GAT), .Z(n383) );
  XNOR2_X1 U450 ( .A(G36GAT), .B(G190GAT), .ZN(n382) );
  XNOR2_X1 U451 ( .A(n383), .B(n382), .ZN(n385) );
  XNOR2_X1 U452 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n384), .B(G211GAT), .ZN(n436) );
  XNOR2_X1 U454 ( .A(n385), .B(n436), .ZN(n386) );
  XNOR2_X1 U455 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U457 ( .A(n391), .B(n390), .Z(n393) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n393), .B(n392), .ZN(n524) );
  NOR2_X1 U460 ( .A1(n548), .A2(n524), .ZN(n395) );
  XNOR2_X1 U461 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n418) );
  XOR2_X1 U463 ( .A(KEYINPUT3), .B(KEYINPUT94), .Z(n397) );
  XNOR2_X1 U464 ( .A(KEYINPUT93), .B(G155GAT), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U466 ( .A(KEYINPUT2), .B(n398), .Z(n438) );
  XOR2_X1 U467 ( .A(KEYINPUT5), .B(G148GAT), .Z(n400) );
  NAND2_X1 U468 ( .A1(G225GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U470 ( .A(KEYINPUT4), .B(n401), .ZN(n416) );
  XOR2_X1 U471 ( .A(G57GAT), .B(KEYINPUT1), .Z(n403) );
  XNOR2_X1 U472 ( .A(G141GAT), .B(KEYINPUT6), .ZN(n402) );
  XNOR2_X1 U473 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U474 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n405) );
  XNOR2_X1 U475 ( .A(G1GAT), .B(G120GAT), .ZN(n404) );
  XNOR2_X1 U476 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U477 ( .A(n407), .B(n406), .Z(n414) );
  XOR2_X1 U478 ( .A(G162GAT), .B(G85GAT), .Z(n411) );
  XOR2_X1 U479 ( .A(G127GAT), .B(KEYINPUT0), .Z(n409) );
  XNOR2_X1 U480 ( .A(G113GAT), .B(KEYINPUT85), .ZN(n408) );
  XNOR2_X1 U481 ( .A(n409), .B(n408), .ZN(n450) );
  XNOR2_X1 U482 ( .A(n450), .B(G134GAT), .ZN(n410) );
  XNOR2_X1 U483 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U484 ( .A(G29GAT), .B(n412), .ZN(n413) );
  XNOR2_X1 U485 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U486 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U487 ( .A(n438), .B(n417), .ZN(n546) );
  NAND2_X1 U488 ( .A1(n418), .A2(n546), .ZN(n419) );
  XNOR2_X1 U489 ( .A(n420), .B(n419), .ZN(n575) );
  XOR2_X1 U490 ( .A(KEYINPUT92), .B(G106GAT), .Z(n422) );
  XNOR2_X1 U491 ( .A(G50GAT), .B(G204GAT), .ZN(n421) );
  XNOR2_X1 U492 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U493 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n424) );
  XNOR2_X1 U494 ( .A(KEYINPUT90), .B(KEYINPUT95), .ZN(n423) );
  XNOR2_X1 U495 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U496 ( .A(n426), .B(n425), .Z(n428) );
  XOR2_X1 U497 ( .A(n430), .B(n429), .Z(n432) );
  NAND2_X1 U498 ( .A1(G228GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U499 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U500 ( .A(n435), .B(KEYINPUT23), .Z(n440) );
  XNOR2_X1 U501 ( .A(n436), .B(KEYINPUT91), .ZN(n437) );
  NAND2_X1 U502 ( .A1(n575), .A2(n476), .ZN(n442) );
  XOR2_X1 U503 ( .A(KEYINPUT88), .B(KEYINPUT86), .Z(n444) );
  XNOR2_X1 U504 ( .A(KEYINPUT20), .B(KEYINPUT87), .ZN(n443) );
  XNOR2_X1 U505 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U506 ( .A(KEYINPUT89), .B(G176GAT), .Z(n446) );
  XNOR2_X1 U507 ( .A(G169GAT), .B(G15GAT), .ZN(n445) );
  XNOR2_X1 U508 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U509 ( .A(n448), .B(n447), .Z(n452) );
  XNOR2_X1 U510 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U511 ( .A(n452), .B(n451), .ZN(n458) );
  XOR2_X1 U512 ( .A(n454), .B(n453), .Z(n456) );
  NAND2_X1 U513 ( .A1(G227GAT), .A2(G233GAT), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U515 ( .A(n458), .B(n457), .Z(n460) );
  XNOR2_X1 U516 ( .A(G43GAT), .B(G99GAT), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n460), .B(n459), .ZN(n561) );
  INV_X1 U518 ( .A(n561), .ZN(n532) );
  OR2_X1 U519 ( .A1(n562), .A2(n293), .ZN(n464) );
  XOR2_X1 U520 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n462) );
  INV_X1 U521 ( .A(n465), .ZN(n563) );
  AND2_X1 U522 ( .A1(n582), .A2(n563), .ZN(n498) );
  INV_X1 U523 ( .A(n570), .ZN(n586) );
  NOR2_X1 U524 ( .A1(n541), .A2(n586), .ZN(n466) );
  XNOR2_X1 U525 ( .A(KEYINPUT16), .B(n466), .ZN(n482) );
  OR2_X1 U526 ( .A1(n561), .A2(n524), .ZN(n467) );
  NAND2_X1 U527 ( .A1(n467), .A2(n476), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT102), .ZN(n469) );
  XOR2_X1 U529 ( .A(KEYINPUT25), .B(n469), .Z(n474) );
  NOR2_X1 U530 ( .A1(n476), .A2(n532), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n470), .B(KEYINPUT26), .ZN(n574) );
  XOR2_X1 U532 ( .A(n524), .B(KEYINPUT27), .Z(n471) );
  XNOR2_X1 U533 ( .A(KEYINPUT100), .B(n471), .ZN(n478) );
  NAND2_X1 U534 ( .A1(n574), .A2(n478), .ZN(n547) );
  NAND2_X1 U535 ( .A1(n475), .A2(n546), .ZN(n481) );
  XNOR2_X1 U536 ( .A(KEYINPUT28), .B(KEYINPUT68), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(n528) );
  NAND2_X1 U538 ( .A1(n478), .A2(n528), .ZN(n479) );
  NOR2_X1 U539 ( .A1(n546), .A2(n479), .ZN(n533) );
  NAND2_X1 U540 ( .A1(n561), .A2(n533), .ZN(n480) );
  AND2_X1 U541 ( .A1(n482), .A2(n491), .ZN(n511) );
  NAND2_X1 U542 ( .A1(n498), .A2(n511), .ZN(n489) );
  NOR2_X1 U543 ( .A1(n546), .A2(n489), .ZN(n483) );
  XOR2_X1 U544 ( .A(KEYINPUT34), .B(n483), .Z(n484) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n484), .ZN(G1324GAT) );
  NOR2_X1 U546 ( .A1(n524), .A2(n489), .ZN(n485) );
  XOR2_X1 U547 ( .A(G8GAT), .B(n485), .Z(G1325GAT) );
  NOR2_X1 U548 ( .A1(n561), .A2(n489), .ZN(n487) );
  XNOR2_X1 U549 ( .A(KEYINPUT35), .B(KEYINPUT103), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U551 ( .A(G15GAT), .B(n488), .Z(G1326GAT) );
  NOR2_X1 U552 ( .A1(n528), .A2(n489), .ZN(n490) );
  XOR2_X1 U553 ( .A(G22GAT), .B(n490), .Z(G1327GAT) );
  NAND2_X1 U554 ( .A1(n491), .A2(n586), .ZN(n492) );
  XOR2_X1 U555 ( .A(KEYINPUT106), .B(n492), .Z(n494) );
  BUF_X1 U556 ( .A(n493), .Z(n590) );
  NAND2_X1 U557 ( .A1(n494), .A2(n590), .ZN(n497) );
  XOR2_X1 U558 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n495) );
  NAND2_X1 U559 ( .A1(n521), .A2(n498), .ZN(n499) );
  NOR2_X1 U560 ( .A1(n546), .A2(n508), .ZN(n503) );
  XOR2_X1 U561 ( .A(KEYINPUT104), .B(KEYINPUT109), .Z(n501) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NOR2_X1 U565 ( .A1(n524), .A2(n508), .ZN(n504) );
  XOR2_X1 U566 ( .A(KEYINPUT110), .B(n504), .Z(n505) );
  XNOR2_X1 U567 ( .A(G36GAT), .B(n505), .ZN(G1329GAT) );
  NOR2_X1 U568 ( .A1(n561), .A2(n508), .ZN(n506) );
  XOR2_X1 U569 ( .A(KEYINPUT40), .B(n506), .Z(n507) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NOR2_X1 U571 ( .A1(n508), .A2(n528), .ZN(n509) );
  XOR2_X1 U572 ( .A(G50GAT), .B(n509), .Z(G1331GAT) );
  AND2_X1 U573 ( .A1(n576), .A2(n510), .ZN(n520) );
  NAND2_X1 U574 ( .A1(n520), .A2(n511), .ZN(n517) );
  NOR2_X1 U575 ( .A1(n546), .A2(n517), .ZN(n513) );
  XNOR2_X1 U576 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  NOR2_X1 U579 ( .A1(n524), .A2(n517), .ZN(n515) );
  XOR2_X1 U580 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U581 ( .A1(n561), .A2(n517), .ZN(n516) );
  XOR2_X1 U582 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U583 ( .A1(n528), .A2(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(KEYINPUT112), .ZN(n529) );
  NOR2_X1 U588 ( .A1(n529), .A2(n546), .ZN(n523) );
  XOR2_X1 U589 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U590 ( .A1(n524), .A2(n529), .ZN(n525) );
  XOR2_X1 U591 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  XNOR2_X1 U592 ( .A(G99GAT), .B(KEYINPUT113), .ZN(n527) );
  NOR2_X1 U593 ( .A1(n561), .A2(n529), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(G1338GAT) );
  NOR2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(n530), .Z(n531) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U599 ( .A1(n548), .A2(n534), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n542), .A2(n563), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n535), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n537) );
  NAND2_X1 U603 ( .A1(n542), .A2(n510), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(n538), .ZN(G1341GAT) );
  NAND2_X1 U606 ( .A1(n570), .A2(n542), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n539), .B(KEYINPUT50), .ZN(n540) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n544) );
  NAND2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U612 ( .A(G134GAT), .B(n545), .Z(G1343GAT) );
  INV_X1 U613 ( .A(n546), .ZN(n550) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n558) );
  NOR2_X1 U616 ( .A1(n576), .A2(n558), .ZN(n551) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n551), .Z(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT118), .B(n552), .ZN(G1344GAT) );
  NOR2_X1 U619 ( .A1(n558), .A2(n369), .ZN(n556) );
  XOR2_X1 U620 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n554) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U624 ( .A1(n586), .A2(n558), .ZN(n557) );
  XOR2_X1 U625 ( .A(G155GAT), .B(n557), .Z(G1346GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n565) );
  NOR2_X2 U629 ( .A1(n562), .A2(n561), .ZN(n566) );
  BUF_X1 U630 ( .A(n566), .Z(n571) );
  NAND2_X1 U631 ( .A1(n563), .A2(n571), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n568) );
  NAND2_X1 U634 ( .A1(n566), .A2(n510), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(n569), .ZN(G1349GAT) );
  XOR2_X1 U637 ( .A(G183GAT), .B(KEYINPUT123), .Z(n573) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1350GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n588) );
  NOR2_X1 U641 ( .A1(n576), .A2(n588), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(KEYINPUT125), .B(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n588), .ZN(n584) );
  XNOR2_X1 U648 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(G204GAT), .B(n585), .Z(G1353GAT) );
  NOR2_X1 U651 ( .A1(n586), .A2(n588), .ZN(n587) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n587), .Z(G1354GAT) );
  INV_X1 U653 ( .A(n588), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(KEYINPUT62), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

