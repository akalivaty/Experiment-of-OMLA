//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT68), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G113gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G120gat), .ZN(new_n209));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G113gat), .Z(new_n210));
  AOI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(G120gat), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n211), .A2(KEYINPUT67), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(KEYINPUT67), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n207), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G113gat), .B(G120gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n203), .B1(KEYINPUT1), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT27), .B(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(new_n220), .B(KEYINPUT28), .Z(new_n221));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(G169gat), .ZN(new_n223));
  INV_X1    g022(.A(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(KEYINPUT26), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n225), .A2(KEYINPUT26), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n221), .A2(new_n222), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n222), .A2(KEYINPUT24), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(new_n226), .ZN(new_n232));
  INV_X1    g031(.A(G183gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n219), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(KEYINPUT24), .A3(new_n222), .ZN(new_n235));
  NOR2_X1   g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT23), .B1(new_n236), .B2(KEYINPUT64), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT23), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n225), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n232), .A2(new_n235), .A3(new_n237), .A4(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT25), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n241), .A2(new_n242), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n244), .B1(new_n243), .B2(new_n245), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n217), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n214), .A2(new_n216), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n243), .A2(new_n245), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT65), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n250), .A2(new_n252), .A3(new_n246), .A4(new_n230), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G227gat), .ZN(new_n255));
  INV_X1    g054(.A(G233gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT34), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n249), .A2(new_n257), .A3(new_n253), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT32), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT33), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G15gat), .B(G43gat), .Z(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT69), .ZN(new_n266));
  XOR2_X1   g065(.A(G71gat), .B(G99gat), .Z(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n262), .A2(new_n264), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT34), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n270), .A3(new_n258), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n268), .B(KEYINPUT70), .Z(new_n272));
  OAI211_X1 g071(.A(new_n261), .B(KEYINPUT32), .C1(new_n263), .C2(new_n272), .ZN(new_n273));
  AND4_X1   g072(.A1(new_n260), .A2(new_n269), .A3(new_n271), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n260), .A2(new_n271), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n269), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n276), .B1(new_n269), .B2(new_n273), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n275), .B(KEYINPUT72), .C1(new_n277), .C2(new_n278), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n274), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT75), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(new_n287), .B2(new_n285), .ZN(new_n288));
  XOR2_X1   g087(.A(G141gat), .B(G148gat), .Z(new_n289));
  INV_X1    g088(.A(KEYINPUT76), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n289), .A2(new_n290), .B1(KEYINPUT2), .B2(new_n285), .ZN(new_n291));
  XNOR2_X1  g090(.A(G141gat), .B(G148gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT76), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n288), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  OR3_X1    g093(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n292), .B1(new_n285), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n214), .A2(new_n297), .A3(new_n216), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT4), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT3), .B1(new_n294), .B2(new_n296), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT3), .ZN(new_n302));
  INV_X1    g101(.A(new_n296), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n291), .A2(new_n293), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n302), .B(new_n303), .C1(new_n304), .C2(new_n288), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n250), .A2(new_n301), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n214), .A2(new_n297), .A3(KEYINPUT4), .A4(new_n216), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n300), .A2(new_n306), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n307), .ZN(new_n310));
  INV_X1    g109(.A(new_n298), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n297), .B1(new_n214), .B2(new_n216), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT5), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT5), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n309), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G1gat), .B(G29gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(KEYINPUT0), .ZN(new_n320));
  XNOR2_X1  g119(.A(G57gat), .B(G85gat), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n320), .B(new_n321), .Z(new_n322));
  AOI21_X1  g121(.A(KEYINPUT6), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n317), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n316), .B1(new_n309), .B2(new_n313), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n322), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(KEYINPUT6), .A3(new_n327), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G197gat), .B(G204gat), .ZN(new_n332));
  INV_X1    g131(.A(G211gat), .ZN(new_n333));
  INV_X1    g132(.A(G218gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n332), .B1(KEYINPUT22), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G211gat), .B(G218gat), .Z(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n340), .B(KEYINPUT73), .Z(new_n341));
  NAND3_X1  g140(.A1(new_n252), .A2(new_n246), .A3(new_n230), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n230), .A2(new_n251), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(new_n340), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n339), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n340), .B1(new_n345), .B2(KEYINPUT29), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n342), .A2(new_n341), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n338), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(G8gat), .B(G36gat), .Z(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT74), .ZN(new_n353));
  XNOR2_X1  g152(.A(G64gat), .B(G92gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n355), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n347), .A2(new_n350), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(KEYINPUT30), .A3(new_n358), .ZN(new_n359));
  OR2_X1    g158(.A1(new_n358), .A2(KEYINPUT30), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n331), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G78gat), .B(G106gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT31), .B(G50gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(KEYINPUT78), .B(G22gat), .Z(new_n368));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n338), .B1(new_n305), .B2(new_n343), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n338), .A2(new_n343), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n297), .B1(new_n302), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n369), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G228gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(new_n256), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  OAI221_X1 g175(.A(new_n369), .B1(new_n374), .B2(new_n256), .C1(new_n370), .C2(new_n372), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n368), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT79), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n376), .A2(new_n377), .A3(new_n368), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n378), .B2(KEYINPUT79), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n367), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n376), .A2(new_n377), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G22gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n385), .A2(new_n366), .A3(new_n381), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n283), .A2(new_n363), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT35), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n269), .A2(new_n273), .B1(new_n260), .B2(new_n271), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n274), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT82), .B(KEYINPUT35), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n387), .A2(new_n391), .A3(new_n361), .A4(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n322), .B(KEYINPUT80), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n315), .A2(new_n317), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT81), .B1(new_n323), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n322), .B1(new_n324), .B2(new_n325), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n395), .A2(new_n397), .A3(KEYINPUT81), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n330), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n393), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n281), .A2(new_n282), .ZN(new_n404));
  INV_X1    g203(.A(new_n274), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(KEYINPUT36), .A3(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n391), .A2(KEYINPUT36), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n329), .A2(new_n330), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n387), .B1(new_n410), .B2(new_n361), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n355), .B1(new_n351), .B2(KEYINPUT37), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT38), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n344), .A2(new_n346), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(new_n339), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n348), .A2(new_n349), .A3(new_n339), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT37), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n413), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n419), .A2(new_n358), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT37), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n347), .B2(new_n350), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT38), .B1(new_n412), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n401), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n306), .A2(new_n300), .A3(new_n308), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n310), .ZN(new_n426));
  OR2_X1    g225(.A1(new_n426), .A2(KEYINPUT39), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n311), .A2(new_n312), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n426), .B(KEYINPUT39), .C1(new_n310), .C2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n394), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n427), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT40), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n427), .A2(new_n429), .A3(KEYINPUT40), .A4(new_n430), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n395), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n387), .B1(new_n435), .B2(new_n361), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n411), .B1(new_n424), .B2(new_n437), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n389), .A2(new_n403), .B1(new_n409), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G22gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G15gat), .ZN(new_n441));
  INV_X1    g240(.A(G15gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(G22gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT87), .ZN(new_n445));
  INV_X1    g244(.A(G1gat), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT87), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n441), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n445), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT88), .ZN(new_n450));
  AOI21_X1  g249(.A(G8gat), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n446), .A2(KEYINPUT16), .ZN(new_n452));
  INV_X1    g251(.A(new_n448), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n447), .B1(new_n441), .B2(new_n443), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n449), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n455), .B(new_n449), .C1(new_n450), .C2(G8gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT17), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT83), .ZN(new_n461));
  INV_X1    g260(.A(G50gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(G43gat), .ZN(new_n463));
  INV_X1    g262(.A(G43gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G50gat), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n461), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n465), .A3(new_n461), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(KEYINPUT15), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT14), .ZN(new_n470));
  INV_X1    g269(.A(G29gat), .ZN(new_n471));
  INV_X1    g270(.A(G36gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n473), .A2(new_n474), .B1(G29gat), .B2(G36gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n464), .A2(G50gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT86), .B(G50gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(new_n478), .B2(new_n464), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n469), .B(new_n475), .C1(new_n479), .C2(KEYINPUT15), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n468), .A2(KEYINPUT15), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(new_n466), .ZN(new_n482));
  INV_X1    g281(.A(new_n474), .ZN(new_n483));
  NOR3_X1   g282(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT84), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G29gat), .A2(G36gat), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT84), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n473), .A2(new_n487), .A3(new_n474), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT85), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n482), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n490), .B1(new_n482), .B2(new_n489), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n460), .B(new_n480), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n488), .A2(new_n486), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n487), .B1(new_n473), .B2(new_n474), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT85), .B1(new_n497), .B2(new_n469), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n489), .A3(new_n490), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n460), .B1(new_n500), .B2(new_n480), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n459), .B1(new_n494), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G229gat), .A2(G233gat), .ZN(new_n503));
  INV_X1    g302(.A(new_n459), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n480), .B1(new_n491), .B2(new_n492), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT18), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n505), .B(new_n459), .Z(new_n509));
  XOR2_X1   g308(.A(new_n503), .B(KEYINPUT13), .Z(new_n510));
  AOI22_X1  g309(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n505), .A2(KEYINPUT17), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n504), .B1(new_n513), .B2(new_n493), .ZN(new_n514));
  INV_X1    g313(.A(new_n503), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n459), .B1(new_n500), .B2(new_n480), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n512), .B1(new_n517), .B2(KEYINPUT18), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n502), .A2(KEYINPUT18), .A3(new_n503), .A4(new_n506), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(KEYINPUT89), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n511), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G113gat), .B(G141gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT11), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(new_n223), .ZN(new_n524));
  INV_X1    g323(.A(G197gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT12), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n519), .A2(KEYINPUT89), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n493), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n516), .B1(new_n530), .B2(new_n459), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n531), .A2(new_n512), .A3(KEYINPUT18), .A4(new_n503), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n527), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n511), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n439), .A2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n539));
  AOI21_X1  g338(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT92), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G64gat), .ZN(new_n543));
  OR3_X1    g342(.A1(new_n543), .A2(KEYINPUT90), .A3(G57gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(G57gat), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT90), .B1(new_n543), .B2(G57gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(G71gat), .A2(G78gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(G71gat), .A2(G78gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT91), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT91), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n552), .A3(new_n549), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n542), .A2(new_n547), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n549), .B(new_n548), .C1(new_n555), .C2(new_n540), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT21), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT93), .Z(new_n561));
  XNOR2_X1  g360(.A(new_n559), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G127gat), .B(G155gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n562), .A2(new_n563), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n539), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n566), .ZN(new_n568));
  INV_X1    g367(.A(new_n539), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n554), .A2(KEYINPUT94), .A3(new_n556), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT94), .B1(new_n554), .B2(new_n556), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT21), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n459), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n459), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n567), .A2(new_n570), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G183gat), .B(G211gat), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  INV_X1    g384(.A(G85gat), .ZN(new_n586));
  INV_X1    g385(.A(G92gat), .ZN(new_n587));
  AOI22_X1  g386(.A1(KEYINPUT8), .A2(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT99), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n584), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G99gat), .B(G106gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n593), .B(new_n584), .C1(new_n590), .C2(new_n591), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n530), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT41), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n597), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n601), .B1(new_n602), .B2(new_n505), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n598), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n598), .B2(new_n603), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT97), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n599), .A2(new_n600), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT95), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT96), .ZN(new_n611));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n608), .A2(new_n613), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n580), .B1(new_n577), .B2(new_n579), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n557), .A2(KEYINPUT100), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n554), .A2(new_n619), .A3(new_n556), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n597), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n595), .A2(new_n557), .A3(KEYINPUT100), .A4(new_n596), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT10), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT10), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n624), .A2(new_n573), .A3(new_n574), .ZN(new_n625));
  INV_X1    g424(.A(G230gat), .ZN(new_n626));
  OAI22_X1  g425(.A1(new_n623), .A2(new_n625), .B1(new_n626), .B2(new_n256), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n256), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n621), .A2(new_n622), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(G176gat), .B(G204gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n627), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT101), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n633), .B1(new_n627), .B2(new_n629), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI211_X1 g436(.A(KEYINPUT101), .B(new_n633), .C1(new_n627), .C2(new_n629), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR4_X1   g438(.A1(new_n581), .A2(new_n616), .A3(new_n617), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n538), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n410), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(new_n446), .ZN(G1324gat));
  NAND3_X1  g442(.A1(new_n538), .A2(new_n362), .A3(new_n640), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(G8gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT42), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT16), .B(G8gat), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  MUX2_X1   g447(.A(new_n646), .B(KEYINPUT42), .S(new_n648), .Z(G1325gat));
  OAI21_X1  g448(.A(G15gat), .B1(new_n641), .B2(new_n409), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n391), .A2(new_n442), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n650), .B1(new_n641), .B2(new_n651), .ZN(G1326gat));
  NOR2_X1   g451(.A1(new_n641), .A2(new_n387), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT43), .B(G22gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  NOR2_X1   g454(.A1(new_n581), .A2(new_n617), .ZN(new_n656));
  INV_X1    g455(.A(new_n616), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n656), .A2(new_n657), .A3(new_n639), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n538), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n659), .A2(G29gat), .A3(new_n410), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(KEYINPUT45), .Z(new_n661));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n439), .B2(new_n657), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT35), .ZN(new_n664));
  INV_X1    g463(.A(new_n386), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n378), .A2(KEYINPUT79), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n666), .A2(new_n379), .A3(new_n381), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n665), .B1(new_n667), .B2(new_n367), .ZN(new_n668));
  AOI211_X1 g467(.A(new_n274), .B(new_n668), .C1(new_n281), .C2(new_n282), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n664), .B1(new_n669), .B2(new_n363), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n407), .B1(new_n283), .B2(KEYINPUT36), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n423), .B(new_n358), .C1(new_n412), .C2(new_n418), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n672), .A2(new_n396), .A3(new_n400), .ZN(new_n673));
  OAI22_X1  g472(.A1(new_n673), .A2(new_n436), .B1(new_n363), .B2(new_n387), .ZN(new_n674));
  OAI22_X1  g473(.A1(new_n670), .A2(new_n402), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(KEYINPUT44), .A3(new_n616), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n533), .A2(new_n511), .A3(new_n534), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n534), .B1(new_n533), .B2(new_n511), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n528), .A2(KEYINPUT102), .A3(new_n535), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n656), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n627), .A2(new_n629), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n632), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(KEYINPUT101), .A3(new_n634), .ZN(new_n687));
  INV_X1    g486(.A(new_n638), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n683), .A2(new_n684), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT103), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n663), .A2(new_n676), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n663), .A2(new_n676), .A3(KEYINPUT104), .A4(new_n691), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n694), .A2(new_n331), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n661), .B1(new_n471), .B2(new_n696), .ZN(G1328gat));
  NOR3_X1   g496(.A1(new_n659), .A2(G36gat), .A3(new_n361), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT46), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n694), .A2(new_n362), .A3(new_n695), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n700), .B2(new_n472), .ZN(G1329gat));
  INV_X1    g500(.A(new_n391), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n659), .A2(G43gat), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n694), .A2(new_n671), .A3(new_n695), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(G43gat), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n692), .A2(new_n409), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n464), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  OAI22_X1  g508(.A1(new_n705), .A2(KEYINPUT47), .B1(new_n707), .B2(new_n709), .ZN(G1330gat));
  XNOR2_X1  g509(.A(new_n659), .B(KEYINPUT105), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n387), .A2(new_n478), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n478), .B1(new_n692), .B2(new_n387), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(KEYINPUT48), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n694), .A2(new_n668), .A3(new_n695), .ZN(new_n716));
  AOI22_X1  g515(.A1(new_n716), .A2(new_n478), .B1(new_n711), .B2(new_n712), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n717), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g517(.A1(new_n683), .A2(new_n684), .A3(new_n616), .A4(new_n689), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n675), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n331), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n362), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  AND2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n725), .B2(new_n724), .ZN(G1333gat));
  OAI21_X1  g527(.A(G71gat), .B1(new_n720), .B2(new_n409), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n702), .A2(G71gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n720), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1334gat));
  NAND2_X1  g532(.A1(new_n721), .A2(new_n668), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT107), .B(G78gat), .Z(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1335gat));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n674), .A2(new_n671), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n402), .B1(new_n388), .B2(KEYINPUT35), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n738), .B(new_n616), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n683), .A2(KEYINPUT108), .A3(new_n656), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT108), .B1(new_n683), .B2(new_n656), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n738), .B1(new_n675), .B2(new_n616), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n737), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT110), .B1(new_n439), .B2(new_n657), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n748), .A2(KEYINPUT51), .A3(new_n744), .A4(new_n741), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n689), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n410), .A2(G85gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n744), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n689), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n663), .A2(new_n676), .A3(new_n331), .A4(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n586), .B1(new_n755), .B2(new_n756), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n752), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n752), .A2(new_n759), .A3(KEYINPUT111), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(G1336gat));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765));
  AOI21_X1  g564(.A(G92gat), .B1(new_n750), .B2(new_n362), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n663), .A2(new_n676), .ZN(new_n767));
  INV_X1    g566(.A(new_n754), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n769), .A2(G92gat), .A3(new_n362), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n765), .B1(new_n766), .B2(new_n771), .ZN(new_n772));
  AOI211_X1 g571(.A(new_n361), .B(new_n689), .C1(new_n747), .C2(new_n749), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n770), .B(KEYINPUT52), .C1(new_n773), .C2(G92gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(G1337gat));
  AOI21_X1  g574(.A(G99gat), .B1(new_n750), .B2(new_n391), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n671), .A2(G99gat), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n769), .B2(new_n777), .ZN(G1338gat));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  AOI21_X1  g578(.A(G106gat), .B1(new_n750), .B2(new_n668), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n769), .A2(G106gat), .A3(new_n668), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n779), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n387), .B(new_n689), .C1(new_n747), .C2(new_n749), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n781), .B(KEYINPUT53), .C1(new_n784), .C2(G106gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1339gat));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787));
  INV_X1    g586(.A(new_n526), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n531), .A2(new_n503), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n509), .A2(new_n510), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n535), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n787), .B1(new_n792), .B2(new_n689), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n639), .A2(KEYINPUT112), .A3(new_n535), .A4(new_n791), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n621), .A2(new_n622), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT10), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n625), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n628), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n633), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n798), .A2(new_n799), .A3(new_n628), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(new_n627), .A3(KEYINPUT54), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n634), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT55), .B1(new_n802), .B2(new_n804), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n680), .A2(new_n681), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n616), .B1(new_n795), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n792), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n809), .A2(new_n812), .A3(new_n616), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n684), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n640), .A2(new_n682), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n410), .A2(new_n362), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n819), .A2(new_n668), .A3(new_n702), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n537), .ZN(new_n822));
  INV_X1    g621(.A(new_n669), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT113), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n683), .A2(new_n210), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(G1340gat));
  OAI21_X1  g626(.A(G120gat), .B1(new_n821), .B2(new_n689), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n689), .A2(G120gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n828), .B1(new_n825), .B2(new_n829), .ZN(G1341gat));
  NAND2_X1  g629(.A1(new_n820), .A2(new_n656), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n684), .A2(G127gat), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n831), .A2(G127gat), .B1(new_n824), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT114), .ZN(G1342gat));
  NOR4_X1   g633(.A1(new_n819), .A2(G134gat), .A3(new_n823), .A4(new_n657), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT56), .ZN(new_n836));
  OAI21_X1  g635(.A(G134gat), .B1(new_n821), .B2(new_n657), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1343gat));
  NOR3_X1   g637(.A1(new_n671), .A2(new_n410), .A3(new_n362), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n387), .B1(new_n815), .B2(new_n816), .ZN(new_n840));
  XNOR2_X1  g639(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n802), .A2(new_n845), .A3(new_n804), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n845), .B1(new_n802), .B2(new_n804), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n806), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n807), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n536), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n812), .A2(new_n639), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n616), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n684), .B1(new_n853), .B2(new_n814), .ZN(new_n854));
  AOI211_X1 g653(.A(new_n844), .B(new_n387), .C1(new_n854), .C2(new_n816), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n839), .B1(new_n843), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(G141gat), .B1(new_n856), .B2(new_n537), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n671), .A2(new_n387), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n537), .A2(G141gat), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n817), .A2(new_n818), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n857), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n683), .B(new_n839), .C1(new_n843), .C2(new_n855), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n863), .A2(new_n864), .A3(G141gat), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n863), .B2(G141gat), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n861), .B(KEYINPUT118), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n862), .B1(new_n868), .B2(new_n858), .ZN(G1344gat));
  NOR4_X1   g668(.A1(new_n410), .A2(new_n362), .A3(G148gat), .A4(new_n689), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n817), .A2(new_n859), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n689), .ZN(new_n872));
  INV_X1    g671(.A(G148gat), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n872), .A2(KEYINPUT59), .A3(new_n873), .ZN(new_n874));
  XOR2_X1   g673(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n875));
  AOI211_X1 g674(.A(new_n387), .B(new_n841), .C1(new_n815), .C2(new_n816), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n640), .A2(new_n537), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n854), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n878), .B2(new_n668), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n639), .B(new_n839), .C1(new_n876), .C2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n875), .B1(new_n880), .B2(G148gat), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n871), .B1(new_n874), .B2(new_n881), .ZN(G1345gat));
  INV_X1    g681(.A(G155gat), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n856), .A2(new_n883), .A3(new_n684), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n819), .A2(new_n387), .A3(new_n671), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n656), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(KEYINPUT120), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(G155gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(KEYINPUT120), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(G1346gat));
  OAI21_X1  g689(.A(G162gat), .B1(new_n856), .B2(new_n657), .ZN(new_n891));
  INV_X1    g690(.A(G162gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n885), .A2(new_n892), .A3(new_n616), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(G1347gat));
  NOR2_X1   g693(.A1(new_n823), .A2(new_n361), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n895), .A2(KEYINPUT121), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n331), .B1(new_n895), .B2(KEYINPUT121), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n896), .A2(new_n817), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(G169gat), .B1(new_n898), .B2(new_n683), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n331), .A2(new_n361), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n391), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n387), .B1(new_n901), .B2(KEYINPUT122), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(KEYINPUT122), .B2(new_n901), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n903), .A2(new_n817), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n537), .A2(new_n223), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(G1348gat));
  NAND3_X1  g705(.A1(new_n898), .A2(new_n224), .A3(new_n639), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n904), .A2(new_n639), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n224), .ZN(G1349gat));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(KEYINPUT60), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n233), .B1(new_n904), .B2(new_n656), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n656), .A2(new_n218), .ZN(new_n913));
  AOI211_X1 g712(.A(new_n911), .B(new_n912), .C1(new_n898), .C2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n910), .A2(KEYINPUT60), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n914), .B(new_n915), .ZN(G1350gat));
  NAND2_X1  g715(.A1(new_n904), .A2(new_n616), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G190gat), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n918), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT61), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n918), .B(KEYINPUT124), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n898), .A2(new_n219), .A3(new_n616), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n921), .A2(new_n924), .A3(new_n925), .ZN(G1351gat));
  AND3_X1   g725(.A1(new_n840), .A2(new_n409), .A3(new_n900), .ZN(new_n927));
  AOI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n683), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n409), .A2(new_n929), .A3(new_n900), .ZN(new_n930));
  INV_X1    g729(.A(new_n900), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT125), .B1(new_n671), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n817), .A2(new_n668), .A3(new_n842), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n803), .A2(new_n627), .A3(KEYINPUT54), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n632), .B1(new_n627), .B2(KEYINPUT54), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT116), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n846), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n807), .B1(new_n806), .B2(new_n938), .ZN(new_n939));
  AOI22_X1  g738(.A1(new_n939), .A2(new_n536), .B1(new_n639), .B2(new_n812), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n813), .B1(new_n940), .B2(new_n616), .ZN(new_n941));
  AOI22_X1  g740(.A1(new_n941), .A2(new_n684), .B1(new_n537), .B2(new_n640), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n844), .B1(new_n942), .B2(new_n387), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n933), .B1(new_n934), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n537), .A2(new_n525), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n928), .B1(new_n944), .B2(new_n945), .ZN(G1352gat));
  INV_X1    g745(.A(G204gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n927), .A2(new_n947), .A3(new_n639), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT62), .Z(new_n949));
  AOI211_X1 g748(.A(new_n689), .B(new_n933), .C1(new_n934), .C2(new_n943), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n947), .B2(new_n950), .ZN(G1353gat));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n952));
  INV_X1    g751(.A(new_n933), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n656), .B(new_n953), .C1(new_n876), .C2(new_n879), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955));
  OAI21_X1  g754(.A(G211gat), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT126), .B1(new_n944), .B2(new_n656), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n952), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(KEYINPUT127), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n960), .B(new_n952), .C1(new_n956), .C2(new_n957), .ZN(new_n961));
  OR3_X1    g760(.A1(new_n956), .A2(new_n957), .A3(new_n952), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n927), .A2(new_n333), .A3(new_n656), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1354gat));
  NAND3_X1  g764(.A1(new_n927), .A2(new_n334), .A3(new_n616), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n944), .A2(new_n616), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(new_n334), .ZN(G1355gat));
endmodule


