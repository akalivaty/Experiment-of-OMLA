//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT32), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT70), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT2), .B(G113), .Z(new_n192));
  XNOR2_X1  g006(.A(G116), .B(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT2), .B(G113), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G116), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n195), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n194), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  OAI22_X1  g016(.A1(new_n202), .A2(G137), .B1(KEYINPUT65), .B2(KEYINPUT11), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT66), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G134), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n209), .A2(new_n211), .A3(new_n212), .A4(new_n204), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT11), .A2(G134), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n215), .B1(new_n216), .B2(G137), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n210), .A2(KEYINPUT67), .A3(KEYINPUT11), .A4(G134), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n210), .A2(G134), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(G131), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n214), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n220), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n211), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G131), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT64), .A2(G146), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(G143), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n228), .A2(G143), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G128), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n231), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT68), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n231), .A2(new_n238), .A3(new_n233), .A4(new_n235), .ZN(new_n239));
  AND2_X1   g053(.A1(KEYINPUT64), .A2(G146), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT64), .A2(G146), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n244));
  OAI21_X1  g058(.A(G128), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n228), .A2(G143), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n240), .A2(new_n241), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(G143), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n237), .A2(new_n239), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n201), .B1(new_n226), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  NOR2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n248), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n232), .B1(new_n247), .B2(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n251), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n214), .A2(new_n219), .A3(new_n223), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G131), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n257), .B1(new_n259), .B2(new_n222), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n191), .B1(new_n250), .B2(new_n260), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n248), .A2(new_n253), .B1(new_n255), .B2(new_n251), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n206), .A2(new_n213), .B1(new_n217), .B2(new_n218), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(new_n223), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n214), .A2(new_n219), .A3(new_n221), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n245), .A2(new_n248), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n238), .B1(new_n255), .B2(new_n235), .ZN(new_n269));
  INV_X1    g083(.A(new_n239), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n264), .A2(new_n221), .B1(G131), .B2(new_n224), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n267), .A2(new_n273), .A3(KEYINPUT70), .A4(new_n201), .ZN(new_n274));
  INV_X1    g088(.A(G237), .ZN(new_n275));
  INV_X1    g089(.A(G953), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(G210), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n277), .B(KEYINPUT27), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT26), .B(G101), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n261), .A2(new_n274), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT69), .B1(new_n226), .B2(new_n249), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n271), .A2(new_n285), .A3(new_n272), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n286), .A3(new_n267), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT30), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n194), .A2(new_n200), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n267), .A2(new_n273), .A3(KEYINPUT30), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT31), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n261), .A2(new_n274), .A3(KEYINPUT71), .A4(new_n280), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n283), .A2(new_n292), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n250), .A2(new_n260), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(KEYINPUT28), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n287), .A2(new_n290), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(new_n261), .A3(new_n274), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n299), .B2(KEYINPUT28), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n280), .B(KEYINPUT72), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n295), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n292), .A2(new_n294), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n293), .B1(new_n304), .B2(new_n283), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n190), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n267), .A2(new_n273), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n290), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n261), .A3(new_n274), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT28), .ZN(new_n310));
  INV_X1    g124(.A(new_n297), .ZN(new_n311));
  INV_X1    g125(.A(new_n280), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G902), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT29), .B1(new_n300), .B2(new_n302), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n261), .A2(new_n274), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n292), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n312), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n317), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G472), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n306), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n283), .A2(new_n292), .A3(new_n294), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT31), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n327), .B(new_n295), .C1(new_n300), .C2(new_n302), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT32), .B1(new_n328), .B2(new_n187), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT73), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT9), .B(G234), .ZN(new_n331));
  OAI21_X1  g145(.A(G221), .B1(new_n331), .B2(G902), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n332), .B(KEYINPUT78), .Z(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n246), .A2(KEYINPUT1), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n231), .A2(new_n233), .B1(new_n336), .B2(G128), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n269), .B2(new_n270), .ZN(new_n339));
  INV_X1    g153(.A(G104), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(G107), .ZN(new_n341));
  NAND2_X1  g155(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n341), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G101), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n340), .A2(G107), .ZN(new_n347));
  OAI22_X1  g161(.A1(new_n340), .A2(G107), .B1(KEYINPUT79), .B2(KEYINPUT3), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n345), .A2(new_n346), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G107), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G104), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n347), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G101), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n339), .A2(KEYINPUT81), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n337), .B1(new_n237), .B2(new_n239), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n349), .A2(new_n353), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT10), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n265), .A2(new_n266), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n363));
  OR2_X1    g177(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n351), .B1(new_n364), .B2(new_n342), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n348), .A2(new_n347), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n363), .B(G101), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n370), .A2(KEYINPUT80), .A3(new_n363), .A4(G101), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(G101), .B1(new_n365), .B2(new_n366), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(KEYINPUT4), .A3(new_n349), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n262), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n354), .A2(KEYINPUT10), .ZN(new_n376));
  OAI22_X1  g190(.A1(new_n372), .A2(new_n375), .B1(new_n376), .B2(new_n249), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n360), .A2(new_n362), .A3(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(G110), .B(G140), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n276), .A2(G227), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n379), .B(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n335), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT81), .B1(new_n339), .B2(new_n354), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n357), .A2(new_n356), .A3(new_n358), .ZN(new_n384));
  OAI22_X1  g198(.A1(new_n383), .A2(new_n384), .B1(new_n271), .B2(new_n354), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(KEYINPUT12), .A3(new_n362), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT12), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n237), .A2(new_n239), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n388), .A2(new_n268), .A3(new_n358), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n355), .B2(new_n359), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n387), .B1(new_n390), .B2(new_n361), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT10), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(new_n383), .B2(new_n384), .ZN(new_n394));
  INV_X1    g208(.A(new_n375), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n369), .A2(new_n371), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n358), .A2(new_n393), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n395), .A2(new_n396), .B1(new_n271), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n361), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n381), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(KEYINPUT82), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n382), .A2(new_n392), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n362), .B1(new_n360), .B2(new_n377), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n381), .ZN(new_n405));
  AOI211_X1 g219(.A(G469), .B(G902), .C1(new_n402), .C2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n378), .A2(new_n381), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n403), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n378), .B1(new_n386), .B2(new_n391), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n408), .B(G469), .C1(new_n400), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(G469), .A2(G902), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n334), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n193), .A2(KEYINPUT5), .ZN(new_n414));
  INV_X1    g228(.A(G113), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT5), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n197), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n194), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n358), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n374), .A2(new_n290), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n421), .B1(new_n372), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G122), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n424), .B(new_n421), .C1(new_n372), .C2(new_n422), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(KEYINPUT6), .A3(new_n427), .ZN(new_n428));
  OR2_X1    g242(.A1(KEYINPUT74), .A2(G125), .ZN(new_n429));
  NAND2_X1  g243(.A1(KEYINPUT74), .A2(G125), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n262), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n249), .B2(new_n431), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n276), .A2(G224), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(KEYINPUT83), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n433), .B(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n365), .A2(new_n366), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n363), .B1(new_n437), .B2(new_n346), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n201), .B1(new_n438), .B2(new_n373), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n420), .B1(new_n439), .B2(new_n396), .ZN(new_n440));
  OR3_X1    g254(.A1(new_n440), .A2(KEYINPUT6), .A3(new_n424), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n428), .A2(new_n436), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n358), .A2(new_n419), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(new_n420), .B2(KEYINPUT84), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT84), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n358), .A2(new_n419), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n424), .B(KEYINPUT8), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n447), .A2(new_n448), .B1(new_n440), .B2(new_n424), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n434), .A2(KEYINPUT7), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n431), .B1(new_n388), .B2(new_n268), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n254), .A2(new_n256), .A3(new_n431), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n432), .B(new_n450), .C1(new_n431), .C2(new_n249), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(G902), .B1(new_n449), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G210), .B1(G237), .B2(G902), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n442), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT85), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n442), .A2(new_n457), .ZN(new_n462));
  INV_X1    g276(.A(new_n458), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n442), .A2(new_n457), .A3(KEYINPUT85), .A4(new_n458), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n461), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G214), .B1(G237), .B2(G902), .ZN(new_n467));
  INV_X1    g281(.A(G217), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n331), .A2(new_n468), .A3(G953), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G128), .B(G143), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n242), .A2(G128), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n473), .B(G134), .C1(new_n474), .C2(new_n472), .ZN(new_n475));
  XNOR2_X1  g289(.A(G116), .B(G122), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(new_n350), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n471), .A2(new_n202), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n350), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n234), .A2(G143), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n474), .A2(new_n481), .A3(new_n202), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n202), .B1(new_n474), .B2(new_n481), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n196), .A2(G122), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n350), .B1(new_n486), .B2(KEYINPUT14), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT14), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n476), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT90), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G122), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G116), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n485), .A2(new_n493), .A3(new_n488), .ZN(new_n494));
  OAI21_X1  g308(.A(G107), .B1(new_n485), .B2(new_n488), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT90), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n484), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT91), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n479), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n483), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n500), .A2(new_n478), .B1(new_n350), .B2(new_n476), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n490), .B1(new_n487), .B2(new_n489), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT90), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n501), .B(new_n498), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n470), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT91), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n508), .A2(new_n504), .A3(new_n479), .A4(new_n469), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(KEYINPUT92), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n511), .B(new_n470), .C1(new_n499), .C2(new_n505), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n510), .A2(KEYINPUT93), .A3(new_n316), .A4(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G478), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n513), .A2(new_n515), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n275), .A2(new_n276), .A3(G214), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(new_n242), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G131), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n519), .B(G143), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n263), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT16), .ZN(new_n526));
  AND2_X1   g340(.A1(KEYINPUT74), .A2(G125), .ZN(new_n527));
  NOR2_X1   g341(.A1(KEYINPUT74), .A2(G125), .ZN(new_n528));
  OAI21_X1  g342(.A(G140), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(G125), .A2(G140), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n526), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(KEYINPUT16), .A2(G140), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n431), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n228), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n431), .A2(new_n533), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n530), .B1(new_n431), .B2(G140), .ZN(new_n537));
  OAI211_X1 g351(.A(G146), .B(new_n536), .C1(new_n537), .C2(new_n526), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n520), .A2(KEYINPUT17), .A3(G131), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n525), .A2(new_n535), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(G113), .B(G122), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(new_n340), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n537), .A2(G146), .ZN(new_n543));
  XNOR2_X1  g357(.A(G125), .B(G140), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n247), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(KEYINPUT18), .A2(G131), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(KEYINPUT87), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n522), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT86), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT18), .B(G131), .C1(new_n522), .C2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n520), .A2(KEYINPUT86), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n546), .B(new_n549), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n540), .A2(new_n542), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n542), .B1(new_n540), .B2(new_n553), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n316), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT88), .B(G475), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n276), .A2(G952), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(G234), .B2(G237), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  XOR2_X1   g376(.A(KEYINPUT21), .B(G898), .Z(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT94), .ZN(new_n564));
  NAND2_X1  g378(.A1(G234), .A2(G237), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n565), .A2(G902), .A3(G953), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n562), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n521), .A2(new_n523), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n537), .A2(KEYINPUT19), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT19), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n544), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n247), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(new_n573), .A3(new_n538), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n553), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n542), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n554), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT20), .ZN(new_n579));
  NOR2_X1   g393(.A1(G475), .A2(G902), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n579), .B1(new_n578), .B2(new_n580), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n559), .B(new_n568), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n466), .A2(new_n467), .A3(new_n518), .A4(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n413), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT22), .B(G137), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n276), .A2(G221), .A3(G234), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n535), .A2(new_n538), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n198), .A2(G128), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n234), .A2(KEYINPUT23), .A3(G119), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n198), .A2(G128), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(KEYINPUT23), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G110), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT24), .B(G110), .Z(new_n598));
  XNOR2_X1  g412(.A(G119), .B(G128), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n592), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT75), .B(G110), .ZN(new_n604));
  OAI22_X1  g418(.A1(new_n596), .A2(new_n604), .B1(new_n598), .B2(new_n599), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n538), .A2(new_n545), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n591), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n606), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n601), .B1(new_n535), .B2(new_n538), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT76), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT76), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n603), .A2(new_n611), .A3(new_n606), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n607), .B1(new_n613), .B2(new_n591), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT77), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n468), .B1(G234), .B2(new_n316), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(G902), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT25), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n619), .B1(new_n614), .B2(G902), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n590), .B1(new_n610), .B2(new_n612), .ZN(new_n621));
  OAI211_X1 g435(.A(KEYINPUT25), .B(new_n316), .C1(new_n621), .C2(new_n607), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n616), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n187), .B1(new_n303), .B2(new_n305), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n189), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT73), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n287), .A2(new_n290), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT28), .B1(new_n630), .B2(new_n319), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n631), .A2(new_n311), .A3(new_n302), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(new_n322), .A3(new_n313), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n315), .A2(new_n316), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(G472), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n628), .A2(new_n629), .A3(new_n306), .A4(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n330), .A2(new_n587), .A3(new_n626), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G101), .ZN(G3));
  AOI21_X1  g453(.A(new_n324), .B1(new_n328), .B2(new_n316), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n627), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n642), .A2(new_n625), .A3(new_n413), .ZN(new_n643));
  INV_X1    g457(.A(new_n467), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n462), .B2(new_n463), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n467), .A2(KEYINPUT95), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n459), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n462), .A2(KEYINPUT95), .A3(new_n467), .A4(new_n463), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n583), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n651), .A2(new_n581), .B1(new_n557), .B2(new_n558), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT33), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n510), .A2(new_n653), .A3(new_n512), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT96), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n510), .A2(KEYINPUT96), .A3(new_n653), .A4(new_n512), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n506), .A2(KEYINPUT33), .A3(new_n509), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n514), .A2(G902), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n510), .A2(new_n316), .A3(new_n512), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n514), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n652), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n650), .A2(new_n568), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT97), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n643), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT34), .B(G104), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  INV_X1    g483(.A(new_n652), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n518), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n650), .A2(new_n568), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n643), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT35), .B(G107), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G9));
  INV_X1    g489(.A(new_n617), .ZN(new_n676));
  OR3_X1    g490(.A1(new_n613), .A2(KEYINPUT36), .A3(new_n591), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n613), .B1(KEYINPUT36), .B2(new_n591), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n623), .B2(new_n616), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n303), .ZN(new_n682));
  AOI21_X1  g496(.A(G902), .B1(new_n682), .B2(new_n327), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n627), .B(new_n681), .C1(new_n683), .C2(new_n324), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT98), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n641), .A2(KEYINPUT98), .A3(new_n627), .A4(new_n681), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n687), .A3(new_n587), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT37), .B(G110), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G12));
  AOI21_X1  g504(.A(new_n680), .B1(new_n648), .B2(new_n649), .ZN(new_n691));
  AOI21_X1  g505(.A(KEYINPUT12), .B1(new_n385), .B2(new_n362), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n390), .A2(new_n387), .A3(new_n361), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n399), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n694), .A2(new_n381), .B1(new_n407), .B2(new_n403), .ZN(new_n695));
  OAI21_X1  g509(.A(G469), .B1(new_n695), .B2(G902), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n401), .A2(new_n392), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT82), .B1(new_n399), .B2(new_n400), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n405), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(G469), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n700), .A3(new_n316), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n691), .A2(new_n334), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(G900), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n561), .B1(new_n566), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n652), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n518), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n330), .A2(new_n703), .A3(new_n637), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G128), .ZN(G30));
  XNOR2_X1  g524(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n466), .B(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n518), .A2(new_n652), .ZN(new_n713));
  AND4_X1   g527(.A1(new_n467), .A2(new_n712), .A3(new_n680), .A4(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n324), .B1(new_n309), .B2(new_n301), .ZN(new_n715));
  AOI22_X1  g529(.A1(new_n326), .A2(new_n715), .B1(G472), .B2(G902), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT100), .ZN(new_n717));
  INV_X1    g531(.A(new_n306), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n717), .A2(new_n329), .A3(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n333), .B1(new_n696), .B2(new_n701), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n705), .B(KEYINPUT39), .Z(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n723), .A2(KEYINPUT40), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(KEYINPUT40), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n714), .A2(new_n720), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G143), .ZN(G45));
  AOI211_X1 g541(.A(new_n705), .B(new_n652), .C1(new_n661), .C2(new_n663), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n721), .A2(new_n691), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n330), .A3(new_n637), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  AND3_X1   g545(.A1(new_n330), .A2(new_n626), .A3(new_n637), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n701), .A2(KEYINPUT101), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n700), .B1(new_n699), .B2(new_n316), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI211_X1 g549(.A(KEYINPUT101), .B(new_n700), .C1(new_n699), .C2(new_n316), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n333), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n732), .A2(new_n666), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT41), .B(G113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  NAND3_X1  g555(.A1(new_n732), .A2(new_n672), .A3(new_n738), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G116), .ZN(G18));
  NAND2_X1  g557(.A1(new_n330), .A2(new_n637), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n334), .B(new_n650), .C1(new_n735), .C2(new_n736), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT102), .ZN(new_n747));
  INV_X1    g561(.A(new_n734), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(KEYINPUT101), .A3(new_n701), .ZN(new_n749));
  INV_X1    g563(.A(new_n736), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT102), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n752), .A3(new_n334), .A4(new_n650), .ZN(new_n753));
  INV_X1    g567(.A(new_n518), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n754), .A2(new_n680), .A3(new_n584), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n745), .A2(new_n747), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G119), .ZN(G21));
  INV_X1    g571(.A(new_n295), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n310), .A2(new_n311), .ZN(new_n759));
  AOI22_X1  g573(.A1(KEYINPUT31), .A2(new_n326), .B1(new_n759), .B2(new_n301), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT103), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n302), .B1(new_n310), .B2(new_n311), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT103), .B1(new_n305), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n188), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n713), .A2(new_n568), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n766), .A2(new_n626), .A3(new_n641), .A4(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT104), .B1(new_n769), .B2(new_n746), .ZN(new_n770));
  INV_X1    g584(.A(new_n650), .ZN(new_n771));
  AOI211_X1 g585(.A(new_n333), .B(new_n771), .C1(new_n749), .C2(new_n750), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n765), .A2(new_n640), .A3(new_n625), .A4(new_n767), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT104), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G122), .ZN(G24));
  NAND2_X1  g591(.A1(new_n664), .A2(new_n706), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n765), .A2(new_n778), .A3(new_n640), .A4(new_n680), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n747), .A2(new_n753), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G125), .ZN(G27));
  NOR2_X1   g595(.A1(new_n325), .A2(new_n329), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n625), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n645), .A2(new_n461), .A3(new_n465), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT106), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT106), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n645), .A2(new_n461), .A3(new_n786), .A4(new_n465), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n411), .B(KEYINPUT105), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n410), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n334), .B1(new_n406), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n788), .A2(new_n791), .A3(new_n778), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n783), .A2(KEYINPUT42), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT107), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT42), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n330), .A2(new_n626), .A3(new_n637), .ZN(new_n796));
  INV_X1    g610(.A(new_n788), .ZN(new_n797));
  INV_X1    g611(.A(new_n791), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n728), .A3(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n794), .B(new_n795), .C1(new_n796), .C2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n792), .A2(new_n626), .A3(new_n330), .A4(new_n637), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n794), .B1(new_n802), .B2(new_n795), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n793), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G131), .ZN(G33));
  NOR3_X1   g619(.A1(new_n744), .A2(new_n518), .A3(new_n707), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n788), .A2(new_n791), .A3(new_n625), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G134), .ZN(G36));
  NAND2_X1  g623(.A1(new_n642), .A2(new_n681), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n661), .A2(new_n663), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n652), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n812), .A2(KEYINPUT43), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(KEYINPUT43), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT44), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n810), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n816), .B1(new_n810), .B2(new_n815), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n797), .A3(new_n818), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(KEYINPUT109), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(KEYINPUT109), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n695), .A2(KEYINPUT45), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n695), .A2(KEYINPUT45), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(G469), .A3(new_n823), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n824), .A2(new_n789), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT108), .B1(new_n825), .B2(KEYINPUT46), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n406), .B1(new_n825), .B2(KEYINPUT46), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OR3_X1    g642(.A1(new_n825), .A2(KEYINPUT108), .A3(KEYINPUT46), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n333), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n820), .A2(new_n722), .A3(new_n821), .A4(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G137), .ZN(G39));
  INV_X1    g646(.A(KEYINPUT47), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n830), .B1(KEYINPUT110), .B2(new_n833), .ZN(new_n834));
  NOR4_X1   g648(.A1(new_n745), .A2(new_n626), .A3(new_n778), .A4(new_n788), .ZN(new_n835));
  XNOR2_X1  g649(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n834), .B(new_n835), .C1(new_n830), .C2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(G140), .ZN(G42));
  NAND3_X1  g652(.A1(new_n813), .A2(new_n561), .A3(new_n814), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n765), .A2(new_n640), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n626), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n737), .A2(new_n333), .A3(new_n467), .A4(new_n712), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g662(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n737), .A2(new_n333), .A3(new_n788), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n843), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n681), .A3(new_n844), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n626), .A2(new_n851), .A3(new_n561), .A4(new_n719), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n652), .A3(new_n663), .A4(new_n661), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n850), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n834), .B1(new_n830), .B2(new_n836), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n751), .A2(new_n333), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n797), .A3(new_n846), .ZN(new_n860));
  NOR2_X1   g674(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n846), .A2(new_n861), .A3(new_n847), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n856), .A2(new_n860), .A3(KEYINPUT51), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n788), .B(new_n845), .C1(new_n857), .C2(new_n858), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n850), .A2(new_n862), .A3(new_n853), .A4(new_n855), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n846), .A2(new_n747), .A3(new_n753), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n854), .A2(new_n664), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n560), .B(KEYINPUT118), .Z(new_n870));
  NAND3_X1  g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n852), .A2(new_n783), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n872), .A2(KEYINPUT48), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(KEYINPUT48), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n863), .A2(new_n867), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n413), .A2(new_n625), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n466), .A2(new_n467), .A3(new_n568), .ZN(new_n878));
  INV_X1    g692(.A(new_n664), .ZN(new_n879));
  INV_X1    g693(.A(new_n671), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n877), .A2(new_n881), .A3(new_n627), .A4(new_n641), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n688), .A2(new_n638), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT113), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n688), .A2(new_n638), .A3(KEYINPUT113), .A4(new_n882), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n518), .A2(new_n652), .A3(new_n706), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT114), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n797), .A2(new_n889), .A3(new_n721), .ZN(new_n890));
  INV_X1    g704(.A(new_n844), .ZN(new_n891));
  OAI22_X1  g705(.A1(new_n890), .A2(new_n744), .B1(new_n891), .B2(new_n799), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n892), .A2(new_n681), .B1(new_n806), .B2(new_n807), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n804), .A2(new_n887), .A3(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n709), .A2(new_n730), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n650), .A2(new_n713), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n681), .A2(new_n705), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n720), .A2(new_n798), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n895), .A2(new_n780), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT52), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT52), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n895), .A2(new_n780), .A3(new_n898), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n894), .A2(new_n903), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n732), .B(new_n738), .C1(new_n666), .C2(new_n672), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n776), .A2(new_n905), .A3(new_n756), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT112), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT112), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n776), .A2(new_n905), .A3(new_n756), .A4(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n914));
  INV_X1    g728(.A(new_n906), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n904), .A2(KEYINPUT53), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(KEYINPUT115), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT53), .B1(new_n904), .B2(new_n910), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n894), .A2(new_n903), .A3(new_n912), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n919), .B1(new_n910), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g735(.A(KEYINPUT115), .B(new_n917), .C1(new_n921), .C2(new_n914), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n876), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(G952), .A2(G953), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n737), .A2(KEYINPUT49), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n626), .A2(new_n334), .A3(new_n467), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT111), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NOR4_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n712), .A4(new_n812), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n737), .A2(KEYINPUT49), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n719), .A3(new_n931), .ZN(new_n932));
  OAI22_X1  g746(.A1(new_n923), .A2(new_n924), .B1(new_n925), .B2(new_n932), .ZN(G75));
  NAND2_X1  g747(.A1(new_n907), .A2(new_n909), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n934), .A2(new_n894), .A3(new_n903), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n916), .B1(KEYINPUT53), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n936), .A2(G210), .A3(G902), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n428), .A2(new_n441), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n436), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT55), .Z(new_n940));
  XOR2_X1   g754(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n941));
  NAND3_X1  g755(.A1(new_n937), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n276), .A2(G952), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n316), .B1(new_n913), .B2(new_n916), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT56), .B1(new_n946), .B2(G210), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT119), .B1(new_n947), .B2(new_n940), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT56), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n940), .B1(new_n937), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT119), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n945), .B1(new_n948), .B2(new_n952), .ZN(G51));
  XOR2_X1   g767(.A(new_n789), .B(KEYINPUT57), .Z(new_n954));
  INV_X1    g768(.A(new_n917), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n914), .B1(new_n913), .B2(new_n916), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n699), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n946), .A2(G469), .A3(new_n823), .A4(new_n822), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n943), .B1(new_n958), .B2(new_n959), .ZN(G54));
  NAND3_X1  g774(.A1(new_n946), .A2(KEYINPUT58), .A3(G475), .ZN(new_n961));
  INV_X1    g775(.A(new_n578), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n963), .A2(new_n964), .A3(new_n943), .ZN(G60));
  NAND2_X1  g779(.A1(new_n658), .A2(new_n659), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT121), .Z(new_n967));
  NAND2_X1  g781(.A1(G478), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT59), .Z(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n955), .B2(new_n956), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n944), .ZN(new_n972));
  INV_X1    g786(.A(new_n969), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n918), .A2(new_n922), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n972), .B1(new_n974), .B2(new_n967), .ZN(G63));
  NAND2_X1  g789(.A1(new_n677), .A2(new_n678), .ZN(new_n976));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT123), .ZN(new_n978));
  XOR2_X1   g792(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(new_n980));
  NOR4_X1   g794(.A1(new_n894), .A2(new_n903), .A3(new_n912), .A4(new_n906), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n976), .B(new_n980), .C1(new_n919), .C2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT124), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n936), .A2(KEYINPUT124), .A3(new_n976), .A4(new_n980), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT125), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(KEYINPUT61), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n944), .B1(new_n987), .B2(KEYINPUT61), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n980), .B1(new_n919), .B2(new_n981), .ZN(new_n990));
  INV_X1    g804(.A(new_n615), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n986), .A2(new_n988), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n988), .B1(new_n986), .B2(new_n992), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(G66));
  AOI21_X1  g809(.A(new_n276), .B1(new_n564), .B2(G224), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n910), .A2(new_n887), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n997), .B2(new_n276), .ZN(new_n998));
  INV_X1    g812(.A(G898), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n938), .B1(new_n999), .B2(G953), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n998), .B(new_n1000), .ZN(G69));
  NAND2_X1  g815(.A1(new_n289), .A2(new_n291), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n570), .A2(new_n572), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT126), .Z(new_n1004));
  XNOR2_X1  g818(.A(new_n1002), .B(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n895), .A2(new_n780), .A3(new_n726), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT62), .Z(new_n1007));
  AOI211_X1 g821(.A(new_n788), .B(new_n723), .C1(new_n879), .C2(new_n880), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n732), .ZN(new_n1009));
  AND4_X1   g823(.A1(new_n831), .A2(new_n1007), .A3(new_n837), .A4(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1005), .B1(new_n1010), .B2(G953), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n276), .A2(G900), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT127), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n830), .A2(new_n722), .A3(new_n783), .A4(new_n896), .ZN(new_n1014));
  AND4_X1   g828(.A1(new_n780), .A2(new_n1014), .A3(new_n808), .A4(new_n895), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1015), .A2(new_n804), .A3(new_n831), .A4(new_n837), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1013), .B1(new_n1016), .B2(new_n276), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1011), .B1(new_n1017), .B2(new_n1005), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n276), .B1(G227), .B2(G900), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1018), .B(new_n1019), .ZN(G72));
  NAND2_X1  g834(.A1(G472), .A2(G902), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT63), .Z(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  AOI211_X1 g837(.A(new_n1023), .B(new_n921), .C1(new_n326), .C2(new_n322), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1022), .B1(new_n1016), .B2(new_n997), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n321), .A2(new_n280), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n943), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n997), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1023), .B1(new_n1010), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n321), .A2(new_n280), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1024), .A2(new_n1031), .ZN(G57));
endmodule


