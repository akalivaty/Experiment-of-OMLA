//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  XOR2_X1   g009(.A(KEYINPUT67), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G219), .A3(G221), .A4(G220), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2104), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n457), .A2(G2105), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G101), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G137), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n460), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  NAND2_X1  g046(.A1(new_n457), .A2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(new_n461), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n475), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  NAND4_X1  g058(.A1(new_n472), .A2(new_n474), .A3(G138), .A4(new_n461), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n460), .A2(new_n486), .A3(G138), .A4(new_n461), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n472), .A2(new_n474), .A3(G126), .A4(G2105), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n492), .A3(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n489), .A2(KEYINPUT68), .A3(new_n493), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n488), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT69), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n488), .A2(new_n496), .A3(new_n500), .A4(new_n497), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  XOR2_X1   g078(.A(KEYINPUT70), .B(G651), .Z(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G651), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n505), .A2(G543), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n503), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT70), .B(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n507), .B1(new_n511), .B2(new_n506), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT71), .A3(G50), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  OAI21_X1  g091(.A(G543), .B1(new_n516), .B2(KEYINPUT72), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(new_n513), .A3(KEYINPUT5), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n510), .B(new_n515), .C1(new_n504), .C2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n517), .A2(new_n519), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n512), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n505), .A2(KEYINPUT73), .A3(new_n507), .A4(new_n520), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n525), .A2(new_n526), .A3(G88), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n522), .A2(new_n527), .ZN(G166));
  AND2_X1   g103(.A1(new_n525), .A2(new_n526), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G89), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT74), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT74), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n532), .A2(KEYINPUT7), .A3(new_n533), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(G51), .B2(new_n514), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n530), .A2(new_n540), .ZN(G168));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n524), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n514), .A2(G52), .B1(new_n511), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n525), .A2(new_n526), .ZN(new_n546));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(new_n529), .A2(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n524), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n514), .A2(G43), .B1(new_n511), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  INV_X1    g137(.A(G91), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT75), .B1(new_n546), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n525), .A2(new_n526), .A3(new_n565), .A4(G91), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n524), .B(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT9), .B1(new_n508), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n514), .A2(new_n575), .A3(G53), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n572), .A2(G651), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n567), .A2(new_n577), .ZN(G299));
  NAND2_X1  g153(.A1(new_n530), .A2(new_n540), .ZN(G286));
  INV_X1    g154(.A(G166), .ZN(G303));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n581));
  INV_X1    g156(.A(G87), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n546), .B2(new_n582), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n520), .A2(G74), .ZN(new_n584));
  AOI22_X1  g159(.A1(G651), .A2(new_n584), .B1(new_n514), .B2(G49), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n529), .A2(KEYINPUT77), .A3(G87), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(new_n529), .A2(G86), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n520), .A2(G61), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT78), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n504), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(G48), .B2(new_n514), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n589), .A2(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G60), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n524), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(new_n511), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n599), .A2(new_n600), .B1(new_n514), .B2(G47), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n598), .A2(KEYINPUT79), .A3(new_n511), .ZN(new_n602));
  AND2_X1   g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n529), .A2(G85), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n570), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(G54), .B2(new_n514), .ZN(new_n610));
  XOR2_X1   g185(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n546), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n529), .A2(G92), .A3(new_n611), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n610), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT81), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n606), .B1(new_n618), .B2(G868), .ZN(G284));
  OAI21_X1  g194(.A(new_n606), .B1(new_n618), .B2(G868), .ZN(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  AND2_X1   g196(.A1(new_n567), .A2(new_n577), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(G297));
  XNOR2_X1  g198(.A(G297), .B(KEYINPUT82), .ZN(G280));
  NOR2_X1   g199(.A1(new_n617), .A2(G559), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(G860), .B2(new_n618), .ZN(G148));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n555), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n625), .B2(new_n627), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n460), .A2(new_n458), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT13), .Z(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n476), .A2(G123), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n478), .A2(G135), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n461), .A2(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n633), .A2(G2100), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n634), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT83), .ZN(G156));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2435), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT84), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT18), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(new_n663), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n668), .A2(KEYINPUT17), .A3(new_n665), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n665), .B1(new_n668), .B2(KEYINPUT17), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n669), .A2(new_n670), .A3(new_n664), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2096), .B(G2100), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n679), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n684));
  OAI221_X1 g259(.A(new_n680), .B1(new_n677), .B2(new_n681), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n684), .B2(new_n683), .ZN(new_n686));
  XOR2_X1   g261(.A(G1981), .B(G1986), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT86), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n689), .B(new_n692), .ZN(G229));
  NAND2_X1  g268(.A1(G168), .A2(G16), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G16), .B2(G21), .ZN(new_n695));
  INV_X1    g270(.A(G1966), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT92), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G5), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G171), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT94), .Z(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(G1961), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(G1961), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n698), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G33), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n458), .A2(G103), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(KEYINPUT25), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT25), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n458), .A2(new_n710), .A3(G103), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n478), .A2(G139), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n712), .B(new_n713), .C1(new_n461), .C2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n707), .B1(new_n716), .B2(new_n706), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT89), .ZN(new_n718));
  INV_X1    g293(.A(G2072), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT91), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT90), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n718), .A2(new_n723), .A3(new_n719), .ZN(new_n724));
  INV_X1    g299(.A(G2084), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n470), .A2(G29), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT24), .ZN(new_n727));
  INV_X1    g302(.A(G34), .ZN(new_n728));
  AOI21_X1  g303(.A(G29), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n727), .B2(new_n728), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n725), .B1(new_n726), .B2(new_n730), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n726), .A2(new_n725), .A3(new_n730), .ZN(new_n732));
  OR2_X1    g307(.A1(G29), .A2(G32), .ZN(new_n733));
  AOI22_X1  g308(.A1(G129), .A2(new_n476), .B1(new_n478), .B2(G141), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n458), .A2(G105), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT26), .Z(new_n737));
  NAND3_X1  g312(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n733), .B1(new_n738), .B2(new_n706), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT27), .B(G1996), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n731), .B(new_n732), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n739), .A2(new_n741), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT31), .B(G11), .Z(new_n744));
  NOR2_X1   g319(.A1(new_n639), .A2(new_n706), .ZN(new_n745));
  INV_X1    g320(.A(G28), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT30), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n744), .B(new_n745), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n724), .A2(new_n742), .A3(new_n743), .A4(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n723), .B1(new_n718), .B2(new_n719), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G27), .A2(G29), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G164), .B2(G29), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT95), .B(G2078), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n695), .A2(new_n696), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT93), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n722), .A2(new_n752), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(KEYINPUT96), .B1(new_n705), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT92), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n697), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n703), .A2(new_n704), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT96), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n720), .B(KEYINPUT91), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(new_n756), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n752), .A2(new_n759), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n765), .A2(new_n766), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G4), .A2(G16), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n618), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1348), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n706), .A2(G35), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G162), .B2(new_n706), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n776), .A2(KEYINPUT29), .ZN(new_n777));
  INV_X1    g352(.A(G2090), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(KEYINPUT29), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n699), .A2(G19), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n556), .B2(new_n699), .ZN(new_n783));
  OAI22_X1  g358(.A1(new_n780), .A2(new_n781), .B1(new_n783), .B2(G1341), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n781), .B2(new_n780), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n699), .A2(G20), .ZN(new_n786));
  OAI211_X1 g361(.A(KEYINPUT23), .B(new_n786), .C1(new_n622), .C2(new_n699), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(KEYINPUT23), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT98), .B(G1956), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n706), .A2(G26), .ZN(new_n792));
  INV_X1    g367(.A(G140), .ZN(new_n793));
  OR3_X1    g368(.A1(new_n462), .A2(KEYINPUT88), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(KEYINPUT88), .B1(new_n462), .B2(new_n793), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n476), .A2(G128), .ZN(new_n796));
  OR2_X1    g371(.A1(G104), .A2(G2105), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n797), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n794), .A2(new_n795), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n792), .B1(new_n799), .B2(G29), .ZN(new_n800));
  MUX2_X1   g375(.A(new_n792), .B(new_n800), .S(KEYINPUT28), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2067), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n778), .B1(new_n777), .B2(new_n779), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G1341), .B2(new_n783), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n785), .A2(new_n791), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n789), .A2(new_n790), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AND4_X1   g382(.A1(new_n761), .A2(new_n770), .A3(new_n774), .A4(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT99), .ZN(new_n809));
  INV_X1    g384(.A(G290), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n699), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n699), .B2(G24), .ZN(new_n812));
  INV_X1    g387(.A(G1986), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n706), .A2(G25), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n476), .A2(G119), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n478), .A2(G131), .ZN(new_n817));
  OR2_X1    g392(.A1(G95), .A2(G2105), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n818), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n815), .B1(new_n821), .B2(new_n706), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n812), .A2(new_n813), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n814), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  MUX2_X1   g401(.A(G23), .B(G288), .S(G16), .Z(new_n827));
  XOR2_X1   g402(.A(KEYINPUT33), .B(G1976), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT87), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n827), .B(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n699), .A2(G22), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G303), .B2(G16), .ZN(new_n832));
  INV_X1    g407(.A(G1971), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n699), .A2(G6), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G305), .B2(G16), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT32), .B(G1981), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n832), .A2(new_n833), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n834), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n830), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT34), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n830), .A2(new_n840), .A3(KEYINPUT34), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n826), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI211_X1 g422(.A(KEYINPUT36), .B(new_n826), .C1(new_n843), .C2(new_n844), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n808), .B(new_n809), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n761), .A2(new_n770), .A3(new_n774), .A4(new_n807), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT99), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n852), .ZN(G311));
  OAI21_X1  g428(.A(new_n808), .B1(new_n847), .B2(new_n848), .ZN(G150));
  NAND2_X1  g429(.A1(new_n618), .A2(G559), .ZN(new_n855));
  XOR2_X1   g430(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(new_n504), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT100), .B(G93), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n529), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n514), .A2(G55), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n861), .A2(KEYINPUT101), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT101), .B1(new_n861), .B2(new_n862), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n859), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n556), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n555), .B(new_n859), .C1(new_n863), .C2(new_n864), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(G860), .B1(new_n857), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n869), .B2(new_n857), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n865), .A2(G860), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT102), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT103), .ZN(G145));
  XNOR2_X1  g451(.A(new_n470), .B(new_n639), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n482), .ZN(new_n878));
  AOI22_X1  g453(.A1(G130), .A2(new_n476), .B1(new_n478), .B2(G142), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n881));
  INV_X1    g456(.A(G118), .ZN(new_n882));
  AOI22_X1  g457(.A1(new_n880), .A2(new_n881), .B1(new_n882), .B2(G2105), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n881), .B2(new_n880), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n632), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n820), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT105), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n799), .B(new_n738), .ZN(new_n890));
  INV_X1    g465(.A(new_n494), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n488), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n890), .B(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n893), .A2(new_n716), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n716), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n889), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n888), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n878), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n889), .A2(new_n896), .ZN(new_n900));
  INV_X1    g475(.A(new_n878), .ZN(new_n901));
  INV_X1    g476(.A(new_n887), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n900), .B(new_n901), .C1(new_n896), .C2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n899), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT40), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n905), .B(KEYINPUT106), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n911), .ZN(G395));
  NOR2_X1   g487(.A1(G288), .A2(G290), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n586), .A2(new_n587), .B1(new_n604), .B2(new_n603), .ZN(new_n914));
  OAI21_X1  g489(.A(G166), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n810), .A2(new_n587), .A3(new_n586), .ZN(new_n916));
  NAND2_X1  g491(.A1(G288), .A2(G290), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n917), .A3(G303), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(G305), .ZN(new_n920));
  INV_X1    g495(.A(G305), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n915), .A2(new_n921), .A3(new_n918), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT42), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n924));
  INV_X1    g499(.A(new_n922), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n921), .B1(new_n915), .B2(new_n918), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n920), .A2(KEYINPUT109), .A3(new_n922), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n923), .B1(new_n929), .B2(KEYINPUT42), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n869), .B(new_n625), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n622), .A2(new_n616), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n610), .A2(new_n614), .A3(new_n615), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(G299), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT41), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT108), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(G299), .B(new_n616), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT41), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n938), .A2(KEYINPUT41), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT107), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(new_n938), .B2(KEYINPUT41), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n941), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n931), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n938), .B2(new_n931), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n930), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n930), .A2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(G868), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n865), .A2(new_n627), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(G295));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n952), .ZN(G331));
  XNOR2_X1  g529(.A(G286), .B(G301), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n868), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n866), .A2(new_n867), .A3(new_n955), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n935), .A2(new_n936), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n959), .B(new_n960), .C1(new_n961), .C2(new_n942), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n866), .A2(new_n867), .A3(new_n955), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n955), .B1(new_n866), .B2(new_n867), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n942), .A2(new_n961), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT110), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n963), .A2(new_n964), .A3(new_n938), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT111), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n959), .B2(new_n938), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n962), .A2(new_n967), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n927), .A2(new_n928), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n968), .B1(new_n946), .B2(new_n959), .ZN(new_n975));
  AOI21_X1  g550(.A(G37), .B1(new_n975), .B2(new_n929), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n974), .A2(new_n976), .A3(KEYINPUT43), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n975), .A2(new_n929), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT43), .B1(new_n978), .B2(new_n976), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT44), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n974), .A2(new_n976), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n978), .B2(new_n976), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n980), .A2(new_n985), .ZN(G397));
  XNOR2_X1  g561(.A(new_n799), .B(G2067), .ZN(new_n987));
  AOI21_X1  g562(.A(G1384), .B1(new_n488), .B2(new_n891), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(KEYINPUT45), .ZN(new_n989));
  INV_X1    g564(.A(G40), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n464), .A2(new_n468), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n987), .A2(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n994), .A2(KEYINPUT113), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(KEYINPUT113), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n738), .B(G1996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n993), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n820), .B(new_n823), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT114), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n993), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(G290), .A2(G1986), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT112), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n813), .B2(new_n810), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1004), .B1(new_n993), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n1009));
  INV_X1    g584(.A(G1384), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n892), .A2(KEYINPUT45), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n991), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n499), .A2(new_n1010), .A3(new_n501), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G2078), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n465), .A2(new_n469), .A3(G40), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n988), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1961), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1017), .A2(new_n1018), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OR2_X1    g600(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n989), .A2(new_n1020), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1018), .A2(G2078), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(G301), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1011), .A3(new_n1028), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(G171), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1009), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT123), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n696), .A2(new_n1039), .B1(new_n1040), .B2(new_n725), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1038), .B1(new_n1041), .B2(G168), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G286), .A2(G8), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1039), .A2(new_n696), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(G2084), .B2(new_n1023), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1042), .A2(new_n1043), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(KEYINPUT51), .B(new_n1044), .C1(new_n1041), .C2(new_n1038), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1030), .A2(G301), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1009), .B1(new_n1033), .B2(G171), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1048), .A2(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n991), .A2(new_n988), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1055), .B1(new_n1056), .B2(G8), .ZN(new_n1057));
  AOI211_X1 g632(.A(KEYINPUT115), .B(new_n1038), .C1(new_n991), .C2(new_n988), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n586), .A2(G1976), .A3(new_n587), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1054), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT52), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n589), .A2(new_n594), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n589), .B2(new_n594), .ZN(new_n1067));
  INV_X1    g642(.A(G1981), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n593), .A2(KEYINPUT116), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n1066), .A2(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1067), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1069), .A2(new_n1068), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1072), .A3(new_n1065), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1073), .A3(new_n1059), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1061), .A2(new_n1063), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(G303), .A2(G8), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1076), .B(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1040), .A2(new_n778), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1015), .A2(G1971), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1038), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1075), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1078), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n499), .A2(new_n1021), .A3(new_n1010), .A4(new_n501), .ZN(new_n1084));
  INV_X1    g659(.A(new_n988), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1020), .B1(new_n1085), .B2(KEYINPUT50), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1015), .A2(G1971), .B1(new_n1087), .B2(G2090), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1088), .A2(KEYINPUT118), .ZN(new_n1089));
  OAI21_X1  g664(.A(G8), .B1(new_n1088), .B2(KEYINPUT118), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1083), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1082), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(KEYINPUT123), .B(new_n1009), .C1(new_n1031), .C2(new_n1034), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1037), .A2(new_n1052), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n567), .A2(new_n577), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n567), .B2(new_n577), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n1101), .B(new_n1012), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1956), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1097), .B(new_n1099), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1012), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n1100), .ZN(new_n1107));
  INV_X1    g682(.A(G1956), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1087), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1097), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1107), .B(new_n1109), .C1(new_n1110), .C2(new_n1098), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1104), .A2(KEYINPUT61), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT61), .B1(new_n1104), .B2(new_n1111), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  NAND2_X1  g690(.A1(new_n1056), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G1996), .ZN(new_n1117));
  AND4_X1   g692(.A1(KEYINPUT120), .A2(new_n1105), .A3(new_n1117), .A4(new_n1106), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT120), .B1(new_n1015), .B2(new_n1117), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1116), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT121), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1105), .A2(new_n1117), .A3(new_n1106), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1015), .A2(KEYINPUT120), .A3(new_n1117), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1126), .A2(new_n1127), .A3(new_n1116), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n555), .B1(new_n1121), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1114), .B1(new_n1129), .B2(KEYINPUT59), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n1131));
  AOI211_X1 g706(.A(new_n1131), .B(new_n555), .C1(new_n1121), .C2(new_n1128), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1095), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1127), .B1(new_n1126), .B2(new_n1116), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1116), .ZN(new_n1135));
  AOI211_X1 g710(.A(KEYINPUT121), .B(new_n1135), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n556), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n1131), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1129), .A2(KEYINPUT59), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1138), .A2(new_n1139), .A3(KEYINPUT122), .A4(new_n1114), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1056), .A2(G2067), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n1023), .B2(new_n773), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT60), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(new_n933), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(KEYINPUT60), .B2(new_n1142), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1133), .A2(new_n1140), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1104), .B1(new_n616), .B2(new_n1142), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1111), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1094), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT117), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1075), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1061), .A2(new_n1063), .A3(KEYINPUT117), .A4(new_n1074), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI211_X1 g730(.A(G1976), .B(G288), .C1(new_n1070), .C2(new_n1073), .ZN(new_n1156));
  NOR2_X1   g731(.A1(G305), .A2(G1981), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1059), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1047), .A2(G8), .A3(G168), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1082), .A2(new_n1091), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT63), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1151), .A2(new_n1163), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(new_n1160), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1165), .A2(new_n1167), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1159), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1043), .B(G8), .C1(new_n1047), .C2(G286), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1047), .A2(new_n1045), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1171), .A2(new_n1172), .A3(new_n1049), .A4(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1174), .A2(new_n1091), .A3(new_n1082), .A4(new_n1031), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1172), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1170), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1082), .A2(new_n1091), .A3(new_n1031), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1171), .A2(new_n1049), .A3(new_n1173), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(KEYINPUT62), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1178), .A2(KEYINPUT124), .A3(new_n1180), .A4(new_n1174), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1169), .A2(new_n1177), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1008), .B1(new_n1149), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n993), .A2(new_n1117), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT46), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n993), .B1(new_n987), .B2(new_n738), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1185), .B1(new_n1186), .B2(KEYINPUT125), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(KEYINPUT125), .B2(new_n1186), .ZN(new_n1188));
  XOR2_X1   g763(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1189));
  XNOR2_X1  g764(.A(new_n1188), .B(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1006), .A2(new_n992), .ZN(new_n1191));
  OR2_X1    g766(.A1(new_n1191), .A2(KEYINPUT48), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1192), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1193), .B1(KEYINPUT48), .B2(new_n1191), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n821), .A2(new_n823), .ZN(new_n1195));
  OAI22_X1  g770(.A1(new_n999), .A2(new_n1195), .B1(G2067), .B2(new_n799), .ZN(new_n1196));
  AOI211_X1 g771(.A(new_n1190), .B(new_n1194), .C1(new_n993), .C2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1183), .A2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g773(.A1(new_n983), .A2(new_n984), .ZN(new_n1200));
  INV_X1    g774(.A(G319), .ZN(new_n1201));
  NOR3_X1   g775(.A1(G229), .A2(new_n1201), .A3(G227), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n1202), .A2(new_n659), .ZN(new_n1203));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n1204));
  XNOR2_X1  g778(.A(new_n1203), .B(new_n1204), .ZN(new_n1205));
  AND2_X1   g779(.A1(new_n905), .A2(new_n906), .ZN(new_n1206));
  NOR2_X1   g780(.A1(new_n905), .A2(new_n906), .ZN(new_n1207));
  OAI21_X1  g781(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g782(.A1(new_n1200), .A2(new_n1208), .ZN(G308));
  OAI211_X1 g783(.A(new_n907), .B(new_n1205), .C1(new_n984), .C2(new_n983), .ZN(G225));
endmodule


