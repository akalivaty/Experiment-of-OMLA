//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT88), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(KEYINPUT88), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(G1gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n203), .A2(new_n208), .A3(new_n204), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT89), .ZN(new_n211));
  AOI21_X1  g010(.A(G8gat), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n207), .B(new_n209), .C1(new_n211), .C2(G8gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  AND2_X1   g016(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G29gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT15), .ZN(new_n224));
  INV_X1    g023(.A(G43gat), .ZN(new_n225));
  INV_X1    g024(.A(G50gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G43gat), .A2(G50gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n224), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT87), .B(G50gat), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n224), .B(new_n228), .C1(new_n231), .C2(G43gat), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n232), .A2(new_n223), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n230), .B1(new_n233), .B2(new_n229), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n234), .A2(KEYINPUT17), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(KEYINPUT17), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n215), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(new_n237), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n242), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n237), .B(KEYINPUT13), .Z(new_n245));
  NOR2_X1   g044(.A1(new_n216), .A2(new_n235), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n215), .A2(new_n234), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n243), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(G197gat), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT11), .B(G169gat), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n253), .B(KEYINPUT12), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n254), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n243), .A2(new_n244), .A3(new_n248), .A4(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G197gat), .B(G204gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT22), .ZN(new_n260));
  INV_X1    g059(.A(G211gat), .ZN(new_n261));
  INV_X1    g060(.A(G218gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G211gat), .B(G218gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n259), .A3(new_n263), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n271));
  INV_X1    g070(.A(KEYINPUT27), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(G183gat), .ZN(new_n273));
  INV_X1    g072(.A(G183gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(KEYINPUT27), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT65), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(KEYINPUT27), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT65), .ZN(new_n278));
  AOI21_X1  g077(.A(G190gat), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n271), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT27), .B(G183gat), .ZN(new_n281));
  INV_X1    g080(.A(G190gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(KEYINPUT28), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n270), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n282), .B1(new_n273), .B2(KEYINPUT65), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n272), .A2(G183gat), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n278), .B1(new_n277), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n286), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(KEYINPUT67), .A3(new_n283), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(G169gat), .B2(G176gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n294), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n285), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n294), .A2(KEYINPUT23), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(KEYINPUT23), .ZN(new_n299));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT24), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n302), .B1(new_n274), .B2(new_n282), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT64), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n274), .A2(new_n282), .ZN(new_n305));
  NAND3_X1  g104(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n303), .A2(KEYINPUT64), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n301), .B(KEYINPUT25), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT25), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT72), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(KEYINPUT73), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n297), .A2(new_n320), .A3(new_n314), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT29), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n316), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n269), .B(new_n318), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G8gat), .B(G36gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(G64gat), .B(G92gat), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n325), .B(new_n326), .Z(new_n327));
  INV_X1    g126(.A(new_n269), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n316), .B1(new_n319), .B2(new_n321), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n317), .B1(new_n315), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n328), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n324), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT74), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT30), .ZN(new_n335));
  INV_X1    g134(.A(G113gat), .ZN(new_n336));
  INV_X1    g135(.A(G120gat), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT1), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G113gat), .A2(G120gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(G127gat), .B(G134gat), .Z(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n344));
  OAI21_X1  g143(.A(G120gat), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G127gat), .B(G134gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n338), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT69), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n342), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n345), .A2(KEYINPUT69), .A3(new_n346), .A4(new_n338), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G155gat), .ZN(new_n352));
  INV_X1    g151(.A(G162gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT2), .B1(new_n352), .B2(new_n353), .ZN(new_n357));
  XNOR2_X1  g156(.A(G141gat), .B(G148gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n357), .B1(new_n358), .B2(KEYINPUT75), .ZN(new_n359));
  INV_X1    g158(.A(G148gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G141gat), .ZN(new_n361));
  INV_X1    g160(.A(G141gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G148gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT75), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n356), .B1(new_n359), .B2(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(G148gat), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n361), .ZN(new_n371));
  INV_X1    g170(.A(new_n356), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n372), .A3(new_n357), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n351), .A2(new_n367), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT2), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n377), .B1(G155gat), .B2(G162gat), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n378), .B1(new_n364), .B2(new_n365), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n358), .A2(KEYINPUT75), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n372), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n357), .B1(new_n354), .B2(new_n355), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n382), .B1(new_n361), .B2(new_n370), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT77), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT77), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n367), .A2(new_n385), .A3(new_n373), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n384), .A2(new_n386), .A3(KEYINPUT4), .A4(new_n351), .ZN(new_n387));
  INV_X1    g186(.A(new_n351), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT3), .B1(new_n381), .B2(new_n383), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n367), .A2(new_n390), .A3(new_n373), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n376), .A2(new_n387), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT5), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n367), .A2(new_n373), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(new_n349), .A3(new_n350), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n374), .ZN(new_n398));
  INV_X1    g197(.A(new_n393), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n395), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n392), .A2(new_n395), .A3(new_n393), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n374), .A2(KEYINPUT4), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n384), .A2(new_n386), .A3(new_n375), .A4(new_n351), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n394), .A2(new_n400), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT0), .ZN(new_n407));
  XNOR2_X1  g206(.A(G57gat), .B(G85gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  NOR2_X1   g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT6), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n400), .A2(new_n394), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n401), .A2(new_n404), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n409), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n412), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n411), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n333), .A2(KEYINPUT74), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n324), .A2(new_n332), .ZN(new_n421));
  INV_X1    g220(.A(new_n327), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n335), .A2(new_n418), .A3(new_n420), .A4(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n267), .B2(new_n268), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n384), .A2(new_n386), .B1(new_n426), .B2(new_n390), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n269), .B1(new_n391), .B2(new_n330), .ZN(new_n428));
  INV_X1    g227(.A(G228gat), .ZN(new_n429));
  INV_X1    g228(.A(G233gat), .ZN(new_n430));
  OAI22_X1  g229(.A1(new_n427), .A2(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G22gat), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n391), .A2(new_n433), .A3(new_n330), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n391), .B2(new_n330), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n434), .A2(new_n435), .A3(new_n269), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT79), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n425), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n390), .B1(new_n425), .B2(new_n437), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n396), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n429), .A2(new_n430), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n431), .B(new_n432), .C1(new_n436), .C2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(new_n226), .ZN(new_n447));
  XNOR2_X1  g246(.A(G78gat), .B(G106gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n431), .B1(new_n436), .B2(new_n442), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(G22gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n443), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n452), .A2(KEYINPUT81), .A3(new_n443), .A4(new_n449), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n424), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(G227gat), .A2(G233gat), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT34), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n458), .B2(KEYINPUT70), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n297), .A2(new_n388), .A3(new_n314), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n388), .B1(new_n297), .B2(new_n314), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n458), .B(new_n461), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n315), .A2(new_n351), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n462), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n461), .B1(new_n468), .B2(new_n458), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n458), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(new_n471), .A3(new_n462), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT32), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT33), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  XOR2_X1   g274(.A(G15gat), .B(G43gat), .Z(new_n476));
  XNOR2_X1  g275(.A(G71gat), .B(G99gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n473), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n478), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n472), .B(KEYINPUT32), .C1(new_n474), .C2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(KEYINPUT71), .B(new_n470), .C1(new_n479), .C2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT71), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n466), .B2(new_n469), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n463), .A2(new_n464), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n460), .B1(new_n486), .B2(new_n471), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n487), .A2(KEYINPUT71), .A3(new_n465), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n475), .A3(new_n478), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n485), .A2(new_n488), .A3(new_n481), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n483), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT36), .ZN(new_n492));
  INV_X1    g291(.A(new_n455), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n445), .A2(new_n449), .B1(new_n452), .B2(new_n443), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n420), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n419), .B1(new_n333), .B2(KEYINPUT74), .ZN(new_n497));
  INV_X1    g296(.A(new_n423), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT40), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n393), .B1(new_n404), .B2(new_n392), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT39), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT82), .B1(new_n398), .B2(new_n399), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n397), .A2(new_n374), .A3(new_n505), .A4(new_n393), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(KEYINPUT39), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n503), .B(new_n409), .C1(new_n501), .C2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT83), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n500), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT84), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n415), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n405), .A2(KEYINPUT84), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n514), .A3(new_n416), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n503), .A2(new_n409), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n507), .A2(new_n501), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n509), .B(new_n500), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n511), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n495), .B1(new_n499), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT37), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n324), .A2(new_n521), .A3(new_n332), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n328), .B(new_n318), .C1(new_n322), .C2(new_n323), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n269), .B1(new_n329), .B2(new_n331), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(KEYINPUT37), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT38), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n522), .A2(new_n525), .A3(new_n526), .A4(new_n422), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT6), .B1(new_n405), .B2(new_n409), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n416), .B1(new_n405), .B2(KEYINPUT84), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n415), .A2(new_n512), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n527), .A2(new_n411), .A3(new_n531), .A4(new_n333), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT85), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n297), .A2(new_n320), .A3(new_n314), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n320), .B1(new_n297), .B2(new_n314), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n323), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n315), .A2(new_n330), .ZN(new_n537));
  INV_X1    g336(.A(new_n317), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n269), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n330), .B1(new_n534), .B2(new_n535), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n541), .A2(new_n316), .B1(new_n317), .B2(new_n315), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n540), .B1(new_n542), .B2(new_n269), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n533), .B(new_n422), .C1(new_n543), .C2(new_n521), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n521), .B1(new_n324), .B2(new_n332), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT85), .B1(new_n545), .B2(new_n327), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n546), .A3(new_n522), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n532), .B1(new_n547), .B2(KEYINPUT38), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n457), .B(new_n492), .C1(new_n520), .C2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT86), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n334), .A2(KEYINPUT30), .B1(new_n422), .B2(new_n421), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n551), .A2(new_n491), .A3(new_n495), .A4(new_n420), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT35), .B1(new_n531), .B2(new_n411), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n550), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n456), .B1(new_n483), .B2(new_n490), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n556), .A2(new_n499), .A3(KEYINPUT86), .A4(new_n553), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n491), .A2(new_n495), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT35), .B1(new_n424), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n555), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n258), .B1(new_n549), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G120gat), .B(G148gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(G176gat), .B(G204gat), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n562), .B(new_n563), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G99gat), .B(G106gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G99gat), .ZN(new_n568));
  INV_X1    g367(.A(G106gat), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT8), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n571));
  NAND2_X1  g370(.A1(G85gat), .A2(G92gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(G85gat), .A2(G92gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n570), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  OAI211_X1 g375(.A(G85gat), .B(G92gat), .C1(KEYINPUT96), .C2(KEYINPUT7), .ZN(new_n577));
  AND2_X1   g376(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n567), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n577), .A2(new_n578), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n574), .B1(new_n572), .B2(new_n571), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n581), .A2(new_n582), .A3(new_n566), .A4(new_n570), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT97), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(KEYINPUT97), .B(new_n567), .C1(new_n576), .C2(new_n579), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G64gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(G57gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n588), .A2(G57gat), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT9), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  INV_X1    g392(.A(G71gat), .ZN(new_n594));
  INV_X1    g393(.A(G78gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT90), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT90), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(G71gat), .B2(G78gat), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n592), .A2(new_n593), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(G57gat), .ZN(new_n600));
  OAI211_X1 g399(.A(KEYINPUT91), .B(G64gat), .C1(new_n600), .C2(KEYINPUT92), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT91), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n602), .B1(new_n588), .B2(G57gat), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n601), .B(new_n603), .C1(KEYINPUT92), .C2(new_n589), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT9), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n593), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n599), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n587), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n599), .A2(new_n607), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n585), .A2(new_n611), .A3(new_n586), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT98), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT10), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT99), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n580), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g415(.A(KEYINPUT99), .B(new_n567), .C1(new_n576), .C2(new_n579), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n608), .A2(new_n616), .A3(new_n583), .A4(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n585), .A2(new_n611), .A3(new_n619), .A4(new_n586), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n613), .A2(new_n614), .A3(new_n618), .A4(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND4_X1   g422(.A1(new_n607), .A2(new_n617), .A3(new_n599), .A4(new_n583), .ZN(new_n624));
  AOI22_X1  g423(.A1(KEYINPUT98), .A2(new_n612), .B1(new_n624), .B2(new_n616), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n625), .A2(KEYINPUT100), .A3(new_n614), .A4(new_n620), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n610), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n628), .B1(new_n625), .B2(new_n620), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n565), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n623), .A2(new_n626), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n609), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT101), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n627), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n638), .A3(new_n628), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n631), .A2(new_n565), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n633), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n628), .B1(new_n627), .B2(new_n637), .ZN(new_n642));
  AOI211_X1 g441(.A(KEYINPUT101), .B(new_n610), .C1(new_n623), .C2(new_n626), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n633), .B(new_n640), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n632), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT21), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n215), .B1(new_n647), .B2(new_n611), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n649));
  NAND2_X1  g448(.A1(G231gat), .A2(G233gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n648), .B(new_n651), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n611), .A2(new_n647), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT93), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT94), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT93), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n654), .B(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT94), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G127gat), .B(G155gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT95), .Z(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(G183gat), .B(G211gat), .Z(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n663), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n656), .A2(new_n660), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n664), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n666), .B1(new_n664), .B2(new_n668), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n653), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n671), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(new_n652), .A3(new_n669), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n238), .A2(new_n239), .A3(new_n586), .A4(new_n585), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n235), .A2(new_n587), .ZN(new_n677));
  NAND3_X1  g476(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(G190gat), .B(G218gat), .Z(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n680), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n676), .A2(new_n682), .A3(new_n677), .A4(new_n678), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G134gat), .B(G162gat), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n681), .A2(new_n687), .A3(new_n683), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n646), .A2(new_n675), .A3(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n561), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n418), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G1gat), .ZN(G1324gat));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n335), .A2(new_n420), .A3(new_n423), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT103), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT16), .B(G8gat), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n698), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(G8gat), .ZN(new_n704));
  OR3_X1    g503(.A1(new_n700), .A2(new_n698), .A3(new_n702), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(G1325gat));
  INV_X1    g505(.A(new_n694), .ZN(new_n707));
  OAI21_X1  g506(.A(G15gat), .B1(new_n707), .B2(new_n492), .ZN(new_n708));
  INV_X1    g507(.A(new_n491), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n709), .A2(G15gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n707), .B2(new_n710), .ZN(G1326gat));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n456), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT104), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT43), .B(G22gat), .Z(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1327gat));
  INV_X1    g514(.A(new_n646), .ZN(new_n716));
  AND4_X1   g515(.A1(new_n561), .A2(new_n675), .A3(new_n692), .A4(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n221), .A3(new_n695), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT45), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n549), .A2(new_n560), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n691), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n675), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n646), .A2(new_n724), .A3(new_n258), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT105), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n518), .A2(new_n515), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n510), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n456), .B1(new_n699), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n522), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n422), .B1(new_n543), .B2(new_n521), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n731), .B2(KEYINPUT85), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n526), .B1(new_n732), .B2(new_n544), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n729), .B1(new_n733), .B2(new_n532), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n457), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n424), .A2(KEYINPUT106), .A3(new_n456), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n734), .A2(new_n492), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n691), .B1(new_n738), .B2(new_n560), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n723), .B(new_n726), .C1(new_n739), .C2(KEYINPUT44), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT107), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n492), .B1(new_n520), .B2(new_n548), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n736), .A2(new_n737), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n560), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n692), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n721), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n746), .A2(new_n747), .A3(new_n723), .A4(new_n726), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n741), .A2(new_n748), .A3(new_n695), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n719), .B1(new_n221), .B2(new_n749), .ZN(G1328gat));
  NAND3_X1  g549(.A1(new_n717), .A2(new_n217), .A3(new_n699), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT46), .Z(new_n752));
  AND3_X1   g551(.A1(new_n741), .A2(new_n748), .A3(new_n699), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n217), .B2(new_n753), .ZN(G1329gat));
  OAI21_X1  g553(.A(G43gat), .B1(new_n740), .B2(new_n492), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n717), .A2(new_n225), .A3(new_n491), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(KEYINPUT47), .A3(new_n756), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n717), .A2(new_n225), .A3(new_n491), .ZN(new_n758));
  INV_X1    g557(.A(new_n492), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n741), .A2(new_n748), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n758), .B1(new_n760), .B2(G43gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n757), .B1(new_n761), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g561(.A(new_n231), .B1(new_n740), .B2(new_n495), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n495), .A2(new_n231), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n717), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(KEYINPUT48), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n741), .A2(new_n748), .A3(new_n456), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n767), .A2(new_n768), .A3(new_n231), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n768), .B1(new_n767), .B2(new_n231), .ZN(new_n770));
  INV_X1    g569(.A(new_n765), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n766), .B1(new_n772), .B2(KEYINPUT48), .ZN(G1331gat));
  AND3_X1   g572(.A1(new_n672), .A2(new_n674), .A3(new_n691), .ZN(new_n774));
  AND4_X1   g573(.A1(new_n258), .A2(new_n744), .A3(new_n774), .A4(new_n646), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n695), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n699), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT49), .B(G64gat), .Z(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n778), .B2(new_n780), .ZN(G1333gat));
  NAND3_X1  g580(.A1(new_n775), .A2(new_n594), .A3(new_n491), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n775), .A2(new_n759), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n594), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n784), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g584(.A1(new_n775), .A2(new_n456), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g586(.A1(new_n646), .A2(new_n258), .A3(new_n675), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT109), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n746), .A2(new_n723), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790), .B2(new_n418), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n255), .A2(new_n257), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n745), .A2(new_n792), .A3(new_n724), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT51), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n716), .B1(new_n794), .B2(KEYINPUT110), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(KEYINPUT110), .B2(new_n794), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n418), .A2(G85gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n791), .B1(new_n796), .B2(new_n797), .ZN(G1336gat));
  NOR3_X1   g597(.A1(new_n716), .A2(G92gat), .A3(new_n499), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT111), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n794), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(G92gat), .B1(new_n790), .B2(new_n499), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g603(.A(G99gat), .B1(new_n790), .B2(new_n492), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n491), .A2(new_n568), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n796), .B2(new_n806), .ZN(G1338gat));
  NAND3_X1  g606(.A1(new_n646), .A2(new_n569), .A3(new_n456), .ZN(new_n808));
  XOR2_X1   g607(.A(new_n808), .B(KEYINPUT112), .Z(new_n809));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(G106gat), .B1(new_n790), .B2(new_n495), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT53), .ZN(G1339gat));
  OAI21_X1  g612(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT102), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n644), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n774), .A2(new_n258), .A3(new_n816), .A4(new_n632), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT113), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n246), .A2(new_n247), .A3(new_n245), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n237), .B1(new_n236), .B2(new_n240), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n253), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g622(.A(KEYINPUT115), .B(new_n253), .C1(new_n819), .C2(new_n820), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n257), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n627), .A2(KEYINPUT54), .A3(new_n629), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT114), .B1(new_n826), .B2(new_n564), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n635), .A2(new_n828), .A3(new_n628), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n830), .A3(new_n565), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n828), .B1(new_n627), .B2(new_n629), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n827), .A2(new_n831), .B1(new_n639), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n825), .B(new_n692), .C1(new_n833), .C2(KEYINPUT55), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n642), .B2(new_n643), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n826), .A2(KEYINPUT114), .A3(new_n564), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n830), .B1(new_n829), .B2(new_n565), .ZN(new_n837));
  OAI211_X1 g636(.A(KEYINPUT55), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n816), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n646), .A2(new_n825), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n816), .A3(new_n792), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n833), .A2(KEYINPUT55), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n840), .B1(new_n844), .B2(new_n691), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n818), .B1(new_n845), .B2(new_n724), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n495), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n499), .A2(new_n695), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n709), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n258), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n846), .A2(new_n695), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n552), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n258), .A2(new_n344), .A3(new_n343), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT116), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n851), .B1(new_n854), .B2(new_n856), .ZN(G1340gat));
  NAND3_X1  g656(.A1(new_n853), .A2(new_n337), .A3(new_n646), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n847), .A2(new_n646), .A3(new_n849), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n859), .A2(KEYINPUT117), .A3(G120gat), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT117), .B1(new_n859), .B2(G120gat), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(G1341gat));
  OAI21_X1  g661(.A(G127gat), .B1(new_n850), .B2(new_n675), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n675), .A2(G127gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n854), .B2(new_n864), .ZN(G1342gat));
  OR3_X1    g664(.A1(new_n854), .A2(G134gat), .A3(new_n691), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n867));
  OAI21_X1  g666(.A(G134gat), .B1(new_n850), .B2(new_n691), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(G1343gat));
  NAND2_X1  g669(.A1(new_n852), .A2(KEYINPUT119), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n846), .A2(new_n872), .A3(new_n695), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n759), .A2(new_n495), .A3(new_n699), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n258), .A2(G141gat), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT113), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n817), .B(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n840), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n838), .A2(new_n792), .A3(new_n816), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n881));
  XNOR2_X1  g680(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n880), .A2(new_n883), .B1(new_n646), .B2(new_n825), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n884), .B2(new_n692), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n878), .B1(new_n885), .B2(new_n675), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n495), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n846), .A2(new_n888), .A3(new_n456), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n759), .A2(new_n848), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n887), .A2(new_n792), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n368), .A2(new_n369), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n875), .A2(new_n876), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n894), .B1(new_n891), .B2(new_n892), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n893), .A2(KEYINPUT58), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n891), .A2(new_n892), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n871), .A2(new_n873), .A3(new_n874), .A4(new_n876), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n897), .B(new_n898), .C1(KEYINPUT120), .C2(KEYINPUT58), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n896), .A2(new_n900), .ZN(G1344gat));
  NAND3_X1  g700(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n902), .A2(G148gat), .A3(new_n716), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n716), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(KEYINPUT59), .A3(new_n360), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n883), .A2(new_n792), .A3(new_n816), .A4(new_n838), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n692), .B1(new_n910), .B2(new_n841), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n675), .B1(new_n911), .B2(new_n840), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n817), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n888), .A3(new_n456), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n846), .A2(new_n456), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(new_n888), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n890), .A2(new_n646), .ZN(new_n917));
  OAI21_X1  g716(.A(G148gat), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(KEYINPUT59), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n905), .A2(new_n906), .B1(new_n909), .B2(new_n919), .ZN(G1345gat));
  OAI21_X1  g719(.A(G155gat), .B1(new_n907), .B2(new_n675), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n724), .A2(new_n352), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n902), .B2(new_n922), .ZN(G1346gat));
  NAND3_X1  g722(.A1(new_n875), .A2(new_n353), .A3(new_n692), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(KEYINPUT122), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(KEYINPUT122), .ZN(new_n926));
  OAI21_X1  g725(.A(G162gat), .B1(new_n907), .B2(new_n691), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(G1347gat));
  NAND2_X1  g727(.A1(new_n699), .A2(new_n418), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n709), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n847), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n258), .ZN(new_n932));
  AND4_X1   g731(.A1(new_n418), .A2(new_n846), .A3(new_n699), .A4(new_n556), .ZN(new_n933));
  INV_X1    g732(.A(G169gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(new_n934), .A3(new_n792), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT123), .ZN(G1348gat));
  OAI21_X1  g736(.A(G176gat), .B1(new_n931), .B2(new_n716), .ZN(new_n938));
  INV_X1    g737(.A(G176gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n933), .A2(new_n939), .A3(new_n646), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT124), .Z(G1349gat));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n943), .A2(KEYINPUT60), .ZN(new_n944));
  OAI21_X1  g743(.A(G183gat), .B1(new_n931), .B2(new_n675), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n933), .A2(new_n281), .A3(new_n724), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n943), .A2(KEYINPUT60), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n947), .B(new_n948), .ZN(G1350gat));
  NAND3_X1  g748(.A1(new_n933), .A2(new_n282), .A3(new_n692), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT126), .Z(new_n951));
  NAND3_X1  g750(.A1(new_n847), .A2(new_n692), .A3(new_n930), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(G190gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT61), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n953), .A2(KEYINPUT61), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n951), .A2(new_n954), .A3(new_n955), .ZN(G1351gat));
  NOR2_X1   g755(.A1(new_n759), .A2(new_n929), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n914), .B(new_n957), .C1(new_n915), .C2(new_n888), .ZN(new_n958));
  INV_X1    g757(.A(G197gat), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n958), .A2(new_n959), .A3(new_n258), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n846), .A2(new_n418), .ZN(new_n961));
  NOR4_X1   g760(.A1(new_n961), .A2(new_n495), .A3(new_n499), .A4(new_n759), .ZN(new_n962));
  AOI21_X1  g761(.A(G197gat), .B1(new_n962), .B2(new_n792), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n960), .A2(new_n963), .ZN(G1352gat));
  AOI21_X1  g763(.A(G204gat), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n962), .A2(new_n646), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n966), .B(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(G204gat), .B1(new_n958), .B2(new_n716), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(G1353gat));
  NAND3_X1  g769(.A1(new_n962), .A2(new_n261), .A3(new_n724), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n958), .A2(new_n675), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT63), .B1(new_n972), .B2(G211gat), .ZN(new_n973));
  OAI211_X1 g772(.A(KEYINPUT63), .B(G211gat), .C1(new_n958), .C2(new_n675), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n971), .B1(new_n973), .B2(new_n975), .ZN(G1354gat));
  OAI21_X1  g775(.A(G218gat), .B1(new_n958), .B2(new_n691), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n962), .A2(new_n262), .A3(new_n692), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(G1355gat));
endmodule


