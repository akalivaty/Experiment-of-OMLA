//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992;
  XOR2_X1   g000(.A(KEYINPUT74), .B(G217), .Z(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G128), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT75), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n195), .B1(new_n192), .B2(new_n194), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT24), .B(G110), .ZN(new_n198));
  OR3_X1    g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n191), .A2(G128), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n192), .B(new_n200), .C1(new_n201), .C2(KEYINPUT23), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G110), .ZN(new_n203));
  INV_X1    g017(.A(G140), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G125), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G140), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT76), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(KEYINPUT76), .A3(G140), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(KEYINPUT16), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n205), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n212), .B1(new_n211), .B2(new_n214), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n199), .B(new_n203), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n217), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n198), .B1(new_n196), .B2(new_n197), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(G110), .B2(new_n202), .ZN(new_n221));
  XNOR2_X1  g035(.A(G125), .B(G140), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n212), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n219), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n218), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G953), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(G221), .A3(G234), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n228), .B(KEYINPUT77), .ZN(new_n229));
  XOR2_X1   g043(.A(KEYINPUT22), .B(G137), .Z(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n225), .B1(new_n218), .B2(new_n224), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI211_X1 g048(.A(new_n225), .B(new_n231), .C1(new_n218), .C2(new_n224), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n188), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(KEYINPUT25), .B(new_n188), .C1(new_n234), .C2(new_n235), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n190), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OR2_X1    g055(.A1(new_n234), .A2(new_n235), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n190), .A2(new_n188), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n243), .B(KEYINPUT79), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n227), .A2(G227), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n248), .B(KEYINPUT81), .ZN(new_n249));
  XNOR2_X1  g063(.A(G110), .B(G140), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n249), .B(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G104), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT3), .B1(new_n252), .B2(G107), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT3), .ZN(new_n254));
  INV_X1    g068(.A(G107), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G104), .ZN(new_n256));
  INV_X1    g070(.A(G101), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(G107), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n253), .A2(new_n256), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n252), .A2(G107), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n255), .A2(G104), .ZN(new_n261));
  OAI21_X1  g075(.A(G101), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G143), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT65), .B1(new_n264), .B2(G146), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n212), .A3(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(G146), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n265), .A2(new_n267), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT1), .B1(new_n264), .B2(G146), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G128), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n263), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT82), .B1(new_n275), .B2(KEYINPUT10), .ZN(new_n276));
  INV_X1    g090(.A(new_n263), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n274), .A2(new_n270), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT82), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT10), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n253), .A2(new_n256), .A3(new_n258), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G101), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT4), .A3(new_n259), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT4), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(new_n287), .A3(G101), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT64), .B1(new_n264), .B2(G146), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT64), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(new_n212), .A3(G143), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n292), .A3(new_n268), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT0), .B(G128), .Z(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(KEYINPUT0), .A2(G128), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(new_n271), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n293), .A2(KEYINPUT68), .A3(new_n273), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT68), .B1(new_n293), .B2(new_n273), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n270), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n263), .A2(new_n281), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n289), .A2(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT11), .ZN(new_n304));
  INV_X1    g118(.A(G134), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n304), .B1(new_n305), .B2(G137), .ZN(new_n306));
  AOI21_X1  g120(.A(G131), .B1(new_n305), .B2(G137), .ZN(new_n307));
  INV_X1    g121(.A(G137), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT11), .A3(G134), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT66), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT66), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n306), .A2(new_n307), .A3(new_n312), .A4(new_n309), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n305), .A2(G137), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n306), .A2(new_n309), .A3(new_n314), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n311), .A2(new_n313), .B1(G131), .B2(new_n315), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n283), .A2(new_n303), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(new_n283), .B2(new_n303), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n251), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n283), .A2(new_n303), .A3(new_n316), .ZN(new_n320));
  INV_X1    g134(.A(new_n251), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT12), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n270), .B(new_n263), .C1(new_n299), .C2(new_n300), .ZN(new_n323));
  AOI211_X1 g137(.A(new_n322), .B(new_n316), .C1(new_n323), .C2(new_n279), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n279), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n311), .A2(new_n313), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n315), .A2(G131), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT12), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n320), .B(new_n321), .C1(new_n324), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n319), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G469), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(new_n188), .ZN(new_n333));
  INV_X1    g147(.A(new_n318), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n321), .A3(new_n320), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n329), .A2(new_n324), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n317), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n335), .B(G469), .C1(new_n337), .C2(new_n321), .ZN(new_n338));
  NAND2_X1  g152(.A1(G469), .A2(G902), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n333), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G113), .B(G122), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(new_n252), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n209), .A2(new_n210), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT87), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(G146), .ZN(new_n346));
  INV_X1    g160(.A(G237), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n227), .A3(G214), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n264), .ZN(new_n349));
  NOR2_X1   g163(.A1(G237), .A2(G953), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(G143), .A3(G214), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(KEYINPUT18), .A2(G131), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n349), .A2(KEYINPUT18), .A3(G131), .A4(new_n351), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(KEYINPUT87), .B(new_n223), .C1(new_n343), .C2(new_n212), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n346), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n348), .A2(new_n264), .ZN(new_n359));
  AOI21_X1  g173(.A(G143), .B1(new_n350), .B2(G214), .ZN(new_n360));
  OAI21_X1  g174(.A(G131), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT17), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT90), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT90), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n352), .A2(new_n364), .A3(KEYINPUT17), .A4(G131), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G131), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n349), .A2(new_n368), .A3(new_n351), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n361), .A2(new_n362), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n219), .A2(new_n215), .A3(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n342), .B(new_n358), .C1(new_n367), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n366), .A2(new_n215), .A3(new_n219), .A4(new_n370), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n342), .B1(new_n374), .B2(new_n358), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n188), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G475), .ZN(new_n377));
  NOR2_X1   g191(.A1(G475), .A2(G902), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n361), .A2(new_n369), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT88), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT88), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n361), .A2(new_n382), .A3(new_n369), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n219), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT89), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n344), .A2(new_n385), .A3(KEYINPUT19), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT19), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n385), .B1(new_n222), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n388), .B1(new_n343), .B2(new_n387), .ZN(new_n389));
  AOI21_X1  g203(.A(G146), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n358), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n342), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI211_X1 g207(.A(KEYINPUT20), .B(new_n379), .C1(new_n393), .C2(new_n372), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n346), .A2(new_n356), .A3(new_n357), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n361), .A2(new_n382), .A3(new_n369), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n382), .B1(new_n361), .B2(new_n369), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n397), .A2(new_n398), .A3(new_n217), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n386), .A2(new_n389), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n212), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n396), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n372), .B1(new_n402), .B2(new_n342), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n395), .B1(new_n403), .B2(new_n378), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n377), .B1(new_n394), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n193), .A2(G143), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n264), .A2(G128), .ZN(new_n407));
  OR3_X1    g221(.A1(new_n406), .A2(new_n407), .A3(G134), .ZN(new_n408));
  OAI21_X1  g222(.A(G134), .B1(new_n406), .B2(new_n407), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G116), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(KEYINPUT14), .A3(G122), .ZN(new_n412));
  XNOR2_X1  g226(.A(G116), .B(G122), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(G107), .B(new_n412), .C1(new_n414), .C2(KEYINPUT14), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n410), .B(new_n415), .C1(G107), .C2(new_n414), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT13), .B1(new_n264), .B2(G128), .ZN(new_n417));
  XOR2_X1   g231(.A(new_n417), .B(KEYINPUT91), .Z(new_n418));
  AOI21_X1  g232(.A(new_n407), .B1(KEYINPUT13), .B2(new_n406), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n305), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n414), .A2(G107), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n413), .A2(new_n255), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n408), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n416), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT9), .B(G234), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT80), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n426), .A2(G953), .A3(new_n187), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n416), .B(new_n427), .C1(new_n420), .C2(new_n423), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT92), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n424), .A2(KEYINPUT92), .A3(new_n428), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n188), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G478), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(KEYINPUT15), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n436), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n432), .A2(new_n188), .A3(new_n433), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n405), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G221), .B1(new_n426), .B2(G902), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n340), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n227), .A2(G952), .ZN(new_n444));
  NAND2_X1  g258(.A1(G234), .A2(G237), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(G902), .A3(G953), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(G898), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G214), .B1(G237), .B2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G210), .B1(G237), .B2(G902), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n206), .B(new_n270), .C1(new_n299), .C2(new_n300), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n297), .A2(G125), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G224), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(G953), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT7), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n457), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n464), .ZN(new_n466));
  AOI211_X1 g280(.A(KEYINPUT85), .B(new_n466), .C1(new_n458), .C2(new_n459), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G122), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT8), .ZN(new_n470));
  INV_X1    g284(.A(G113), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT2), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT2), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G113), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT69), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n411), .B2(G119), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n191), .A2(KEYINPUT69), .A3(G116), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n411), .A2(G119), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n475), .A2(new_n477), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n411), .A2(G119), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT5), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n471), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n483), .B1(new_n484), .B2(new_n482), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n277), .A2(new_n480), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n277), .B1(new_n480), .B2(new_n485), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n470), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n484), .A2(new_n472), .A3(new_n474), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n480), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n286), .A2(new_n491), .A3(new_n288), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n486), .A3(new_n469), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n458), .A2(new_n459), .A3(new_n466), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n489), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n188), .B1(new_n468), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n460), .A2(new_n462), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n458), .A2(new_n459), .A3(new_n463), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n492), .A2(new_n486), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n469), .B(KEYINPUT83), .Z(new_n501));
  AOI22_X1  g315(.A1(new_n493), .A2(KEYINPUT6), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n500), .A2(KEYINPUT6), .A3(new_n501), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT84), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g320(.A(KEYINPUT84), .B(new_n499), .C1(new_n502), .C2(new_n503), .ZN(new_n507));
  AOI211_X1 g321(.A(new_n456), .B(new_n496), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  XOR2_X1   g322(.A(new_n455), .B(KEYINPUT86), .Z(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n506), .A2(new_n507), .ZN(new_n511));
  INV_X1    g325(.A(new_n496), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n454), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n443), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G472), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n188), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT32), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n350), .A2(G210), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT27), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT26), .B(G101), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n491), .B1(new_n298), .B2(new_n328), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n308), .A2(G134), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n368), .B1(new_n525), .B2(new_n314), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n311), .B2(new_n313), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n301), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT28), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n491), .ZN(new_n530));
  INV_X1    g344(.A(new_n526), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n326), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT67), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT67), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n301), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n316), .A2(new_n297), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n530), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n270), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n293), .A2(new_n273), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT68), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n293), .A2(KEYINPUT68), .A3(new_n273), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT70), .B1(new_n545), .B2(new_n532), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT70), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n301), .A2(new_n547), .A3(new_n527), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n546), .A2(new_n524), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT28), .B1(new_n539), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n529), .B1(new_n550), .B2(KEYINPUT72), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n552), .B(KEYINPUT28), .C1(new_n539), .C2(new_n549), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n523), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n546), .A2(KEYINPUT30), .A3(new_n538), .A4(new_n548), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n527), .A2(new_n534), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(new_n545), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n537), .B1(new_n557), .B2(new_n535), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n491), .B(new_n555), .C1(new_n558), .C2(KEYINPUT30), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n546), .A2(new_n524), .A3(new_n548), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT71), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n560), .A2(new_n561), .A3(new_n523), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT31), .ZN(new_n564));
  INV_X1    g378(.A(new_n523), .ZN(new_n565));
  NOR4_X1   g379(.A1(new_n549), .A2(KEYINPUT71), .A3(KEYINPUT31), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n559), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n519), .B1(new_n554), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT73), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT73), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n571), .B(new_n519), .C1(new_n554), .C2(new_n568), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n529), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT28), .ZN(new_n575));
  AOI211_X1 g389(.A(KEYINPUT67), .B(new_n526), .C1(new_n311), .C2(new_n313), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n556), .A2(new_n545), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n491), .B1(new_n577), .B2(new_n537), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n575), .B1(new_n578), .B2(new_n560), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n574), .B1(new_n579), .B2(new_n552), .ZN(new_n580));
  INV_X1    g394(.A(new_n553), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n565), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n563), .A2(KEYINPUT31), .B1(new_n566), .B2(new_n559), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n517), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n523), .A2(KEYINPUT29), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n546), .A2(new_n548), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n546), .A2(new_n538), .A3(new_n548), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n586), .A2(new_n524), .B1(new_n587), .B2(new_n491), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n574), .B(new_n585), .C1(new_n588), .C2(new_n575), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n188), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n550), .A2(KEYINPUT72), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n591), .A2(new_n523), .A3(new_n553), .A4(new_n574), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n559), .A2(new_n560), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT29), .B1(new_n593), .B2(new_n565), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n590), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  OAI22_X1  g409(.A1(new_n584), .A2(KEYINPUT32), .B1(new_n595), .B2(new_n516), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n247), .B(new_n515), .C1(new_n573), .C2(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT93), .B(G101), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G3));
  OAI21_X1  g413(.A(new_n188), .B1(new_n554), .B2(new_n568), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G472), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n584), .B1(new_n601), .B2(KEYINPUT94), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT94), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n603), .A3(G472), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n340), .A2(new_n442), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n246), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n602), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n432), .A2(new_n608), .A3(new_n433), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT33), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n609), .A2(G478), .A3(new_n188), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n434), .A2(new_n435), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n405), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT96), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n451), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n493), .A2(KEYINPUT6), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n500), .A2(new_n501), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n500), .A2(KEYINPUT6), .A3(new_n501), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT84), .B1(new_n622), .B2(new_n499), .ZN(new_n623));
  INV_X1    g437(.A(new_n507), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n512), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(KEYINPUT95), .A3(new_n456), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT95), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n496), .B1(new_n506), .B2(new_n507), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n627), .B1(new_n628), .B2(new_n455), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n455), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n626), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n616), .A2(new_n452), .A3(new_n617), .A4(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n607), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT34), .B(G104), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  INV_X1    g449(.A(new_n404), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n403), .A2(new_n395), .A3(new_n378), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n636), .A2(KEYINPUT97), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n394), .A2(new_n639), .B1(G475), .B2(new_n376), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n440), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n631), .A2(new_n643), .A3(new_n452), .A4(new_n617), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n607), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT35), .B(G107), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  NAND2_X1  g461(.A1(new_n218), .A2(new_n224), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n231), .A2(KEYINPUT36), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n650), .A2(new_n244), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n238), .A2(new_n239), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(new_n652), .B2(new_n189), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n443), .A2(new_n514), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n602), .A2(new_n654), .A3(new_n604), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  OAI211_X1 g471(.A(new_n516), .B(new_n188), .C1(new_n554), .C2(new_n568), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n518), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n592), .A2(new_n594), .ZN(new_n660));
  INV_X1    g474(.A(new_n590), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(G472), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n659), .A2(new_n570), .A3(new_n663), .A4(new_n572), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n340), .A2(new_n442), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT98), .B(G900), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n449), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n446), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n641), .A2(new_n642), .A3(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n670), .A2(KEYINPUT99), .A3(new_n631), .A4(new_n452), .ZN(new_n671));
  INV_X1    g485(.A(new_n653), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n664), .A2(new_n665), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n631), .A2(new_n452), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(KEYINPUT99), .B1(new_n675), .B2(new_n670), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n193), .ZN(G30));
  XNOR2_X1  g492(.A(new_n668), .B(KEYINPUT39), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n665), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT40), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n508), .A2(new_n513), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n636), .A2(new_n637), .B1(G475), .B2(new_n376), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n687), .A2(new_n642), .A3(new_n453), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n683), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n573), .ZN(new_n690));
  INV_X1    g504(.A(new_n587), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n560), .B1(new_n691), .B2(new_n530), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n188), .B1(new_n692), .B2(new_n523), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n565), .B1(new_n559), .B2(new_n560), .ZN(new_n694));
  OAI21_X1  g508(.A(G472), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n695), .B(KEYINPUT101), .Z(new_n696));
  NAND3_X1  g510(.A1(new_n690), .A2(new_n659), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n653), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n681), .A2(new_n682), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n689), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n264), .ZN(G45));
  NOR2_X1   g515(.A1(new_n614), .A2(new_n669), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n674), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n664), .A2(new_n704), .A3(new_n665), .A4(new_n672), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT103), .B(G146), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G48));
  AOI21_X1  g521(.A(new_n332), .B1(new_n331), .B2(new_n188), .ZN(new_n708));
  AOI211_X1 g522(.A(G469), .B(G902), .C1(new_n319), .C2(new_n330), .ZN(new_n709));
  INV_X1    g523(.A(new_n442), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n247), .B(new_n711), .C1(new_n573), .C2(new_n596), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n632), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT105), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT104), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n713), .B(new_n716), .ZN(G15));
  INV_X1    g531(.A(new_n596), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n246), .B1(new_n690), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n644), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(KEYINPUT106), .A3(new_n720), .A4(new_n711), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n712), .B2(new_n644), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  AND3_X1   g539(.A1(new_n631), .A2(new_n711), .A3(new_n452), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n405), .A2(new_n451), .A3(new_n440), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n664), .A2(new_n672), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  NAND3_X1  g543(.A1(new_n241), .A2(KEYINPUT108), .A3(new_n245), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n731));
  INV_X1    g545(.A(new_n245), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n731), .B1(new_n240), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n574), .B1(new_n588), .B2(new_n575), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n565), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n517), .B1(new_n583), .B2(new_n736), .ZN(new_n737));
  XOR2_X1   g551(.A(KEYINPUT107), .B(G472), .Z(new_n738));
  AOI21_X1  g552(.A(new_n737), .B1(new_n600), .B2(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n687), .A2(new_n642), .A3(new_n451), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n726), .A2(new_n734), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT109), .B(G122), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G24));
  NAND2_X1  g557(.A1(new_n739), .A2(new_n672), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n702), .A3(new_n726), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  NAND2_X1  g561(.A1(new_n625), .A2(new_n509), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n630), .A3(new_n452), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n748), .A2(KEYINPUT110), .A3(new_n630), .A4(new_n452), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n751), .A2(new_n665), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n753), .A2(new_n664), .A3(new_n247), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n703), .A2(KEYINPUT42), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n659), .A2(new_n663), .A3(new_n569), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n753), .A2(new_n702), .A3(new_n756), .A4(new_n734), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n754), .A2(new_n755), .B1(new_n757), .B2(KEYINPUT42), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G131), .ZN(G33));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n719), .A2(new_n760), .A3(new_n670), .A4(new_n753), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n753), .A2(new_n664), .A3(new_n247), .A4(new_n670), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT111), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NAND2_X1  g579(.A1(new_n602), .A2(new_n604), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT112), .ZN(new_n768));
  XOR2_X1   g582(.A(KEYINPUT112), .B(KEYINPUT43), .Z(new_n769));
  NAND2_X1  g583(.A1(new_n687), .A2(new_n613), .ZN(new_n770));
  MUX2_X1   g584(.A(new_n768), .B(new_n769), .S(new_n770), .Z(new_n771));
  NAND3_X1  g585(.A1(new_n766), .A2(new_n672), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n751), .A2(new_n752), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n772), .A2(new_n773), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n335), .B1(new_n337), .B2(new_n321), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n332), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n780), .B2(new_n779), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT46), .B1(new_n782), .B2(new_n339), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n709), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(KEYINPUT46), .A3(new_n339), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n710), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n786), .A2(new_n679), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n775), .A2(new_n777), .A3(new_n778), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  XNOR2_X1  g603(.A(new_n786), .B(KEYINPUT47), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n664), .A2(new_n776), .A3(new_n247), .A4(new_n703), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  AND3_X1   g607(.A1(new_n777), .A2(new_n447), .A3(new_n711), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n771), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n756), .A2(new_n734), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XOR2_X1   g611(.A(KEYINPUT122), .B(KEYINPUT48), .Z(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n771), .A2(new_n447), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n734), .A2(new_n739), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n726), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n690), .A2(new_n659), .A3(new_n696), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n794), .A2(new_n804), .A3(new_n247), .ZN(new_n805));
  INV_X1    g619(.A(new_n616), .ZN(new_n806));
  OAI221_X1 g620(.A(new_n444), .B1(new_n802), .B2(new_n803), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n799), .A2(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n805), .A2(new_n405), .A3(new_n613), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n795), .A2(new_n744), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n802), .A2(new_n776), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n708), .A2(new_n709), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n710), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n812), .B1(new_n790), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n817));
  INV_X1    g631(.A(new_n686), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n453), .A3(new_n711), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n802), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n802), .A2(new_n819), .ZN(new_n821));
  INV_X1    g635(.A(new_n817), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n811), .B(new_n816), .C1(new_n820), .C2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n808), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT121), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n824), .A2(new_n829), .A3(new_n825), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n826), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n437), .A2(KEYINPUT115), .A3(new_n439), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT115), .B1(new_n437), .B2(new_n439), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n514), .A2(new_n405), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n602), .A2(new_n604), .A3(new_n606), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n837), .A2(new_n838), .A3(new_n655), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n838), .B1(new_n837), .B2(new_n655), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n741), .B(new_n597), .C1(new_n712), .C2(new_n632), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n614), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n405), .A2(new_n613), .A3(KEYINPUT114), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n514), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n602), .A2(new_n847), .A3(new_n604), .A4(new_n606), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n728), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n841), .A2(new_n724), .A3(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n835), .A2(new_n638), .A3(new_n640), .A4(new_n668), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n776), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(new_n664), .A3(new_n665), .A4(new_n672), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n745), .A2(new_n702), .A3(new_n753), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n764), .A2(new_n758), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n674), .A2(new_n687), .A3(new_n642), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n605), .A2(new_n669), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n697), .A2(new_n860), .A3(new_n653), .A4(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n746), .B(new_n705), .C1(new_n673), .C2(new_n676), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n859), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n677), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n746), .A2(new_n705), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT52), .A4(new_n862), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n867), .A3(new_n862), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n865), .A2(new_n868), .B1(new_n869), .B2(KEYINPUT118), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(KEYINPUT118), .A3(KEYINPUT52), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(KEYINPUT53), .B(new_n858), .C1(new_n870), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n865), .A2(new_n868), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n764), .A2(new_n856), .A3(new_n758), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n850), .A2(new_n724), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .A4(new_n841), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT117), .B1(new_n851), .B2(new_n857), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n875), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g695(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n832), .B(new_n873), .C1(new_n881), .C2(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n841), .A2(new_n724), .A3(new_n850), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n878), .B1(new_n885), .B2(new_n876), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n851), .A2(new_n857), .A3(KEYINPUT117), .ZN(new_n887));
  OAI22_X1  g701(.A1(new_n886), .A2(new_n887), .B1(new_n870), .B2(new_n872), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n888), .A2(new_n889), .B1(new_n881), .B2(new_n883), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n831), .B(new_n884), .C1(new_n832), .C2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(G952), .B2(G953), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n770), .A2(new_n453), .A3(new_n710), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n734), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT113), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n813), .B(KEYINPUT49), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n895), .A2(new_n818), .A3(new_n804), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n892), .A2(new_n897), .ZN(G75));
  XOR2_X1   g712(.A(new_n622), .B(new_n499), .Z(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT55), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n874), .B1(new_n886), .B2(new_n887), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n882), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n188), .B1(new_n902), .B2(new_n873), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(G210), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n881), .A2(new_n883), .ZN(new_n907));
  INV_X1    g721(.A(new_n873), .ZN(new_n908));
  OAI211_X1 g722(.A(G902), .B(new_n509), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(new_n905), .A3(new_n900), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n227), .A2(G952), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n906), .A2(new_n913), .ZN(G51));
  XOR2_X1   g728(.A(new_n339), .B(KEYINPUT57), .Z(new_n915));
  AOI21_X1  g729(.A(new_n832), .B1(new_n902), .B2(new_n873), .ZN(new_n916));
  INV_X1    g730(.A(new_n884), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n331), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n903), .B(new_n781), .C1(new_n780), .C2(new_n779), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n911), .B1(new_n919), .B2(new_n920), .ZN(G54));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n922));
  AND2_X1   g736(.A1(KEYINPUT58), .A2(G475), .ZN(new_n923));
  OAI211_X1 g737(.A(G902), .B(new_n923), .C1(new_n907), .C2(new_n908), .ZN(new_n924));
  INV_X1    g738(.A(new_n403), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n911), .B1(new_n924), .B2(new_n925), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n903), .A2(KEYINPUT123), .A3(new_n403), .A4(new_n923), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(G60));
  NOR2_X1   g743(.A1(new_n916), .A2(new_n917), .ZN(new_n930));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT59), .Z(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n609), .A2(new_n610), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n912), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n884), .B1(new_n890), .B2(new_n832), .ZN(new_n936));
  AOI22_X1  g750(.A1(new_n936), .A2(new_n933), .B1(new_n609), .B2(new_n610), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT60), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n650), .B(new_n941), .C1(new_n907), .C2(new_n908), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n902), .B2(new_n873), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n242), .B(KEYINPUT124), .Z(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n942), .B(new_n912), .C1(new_n943), .C2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n941), .B1(new_n907), .B2(new_n908), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n911), .B1(new_n949), .B2(new_n944), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(KEYINPUT61), .A3(new_n942), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n948), .A2(new_n951), .ZN(G66));
  XNOR2_X1  g766(.A(new_n885), .B(KEYINPUT125), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n227), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n450), .B2(new_n461), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n620), .B(new_n621), .C1(G898), .C2(new_n227), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G69));
  OAI21_X1  g772(.A(new_n555), .B1(new_n558), .B2(KEYINPUT30), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT126), .Z(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(new_n400), .Z(new_n961));
  OR3_X1    g775(.A1(new_n700), .A2(KEYINPUT62), .A3(new_n864), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT62), .B1(new_n700), .B2(new_n864), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n835), .A2(new_n405), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n680), .B(new_n776), .C1(new_n846), .C2(new_n965), .ZN(new_n966));
  AOI22_X1  g780(.A1(new_n790), .A2(new_n791), .B1(new_n719), .B2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n962), .A2(new_n788), .A3(new_n963), .A4(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n961), .B1(new_n968), .B2(new_n227), .ZN(new_n969));
  INV_X1    g783(.A(new_n788), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n787), .A2(new_n734), .A3(new_n756), .A4(new_n860), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n792), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n764), .A2(new_n758), .ZN(new_n973));
  OR4_X1    g787(.A1(new_n970), .A2(new_n972), .A3(new_n973), .A4(new_n864), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n974), .A2(G953), .ZN(new_n975));
  INV_X1    g789(.A(new_n961), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(G900), .B2(G953), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n969), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(G227), .A2(G900), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(G953), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n978), .B(new_n980), .ZN(G72));
  NOR2_X1   g795(.A1(new_n593), .A2(new_n523), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT127), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n974), .A2(new_n953), .ZN(new_n984));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT63), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n983), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n968), .A2(new_n953), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n694), .B1(new_n988), .B2(new_n986), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n987), .A2(new_n989), .A3(new_n912), .ZN(new_n990));
  INV_X1    g804(.A(new_n890), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n982), .A2(new_n694), .A3(new_n986), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(G57));
endmodule


