//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  AOI21_X1  g003(.A(G8gat), .B1(new_n204), .B2(KEYINPUT90), .ZN(new_n205));
  XOR2_X1   g004(.A(G15gat), .B(G22gat), .Z(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n205), .B(new_n208), .C1(KEYINPUT90), .C2(new_n204), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n204), .A3(KEYINPUT89), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n210), .B(G8gat), .C1(KEYINPUT89), .C2(new_n204), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT15), .ZN(new_n214));
  INV_X1    g013(.A(G50gat), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n215), .A2(G43gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n216), .B2(KEYINPUT87), .ZN(new_n217));
  NAND2_X1  g016(.A1(G29gat), .A2(G36gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  INV_X1    g019(.A(G29gat), .ZN(new_n221));
  INV_X1    g020(.A(G36gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT14), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n217), .A2(new_n218), .A3(new_n220), .A4(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G43gat), .B(G50gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n220), .A3(new_n218), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n214), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(new_n224), .B2(new_n225), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n213), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(KEYINPUT88), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n231), .A2(KEYINPUT88), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n230), .B1(new_n234), .B2(new_n212), .ZN(new_n235));
  NAND2_X1  g034(.A1(G229gat), .A2(G233gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(KEYINPUT91), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n212), .B(new_n229), .Z(new_n241));
  XOR2_X1   g040(.A(new_n237), .B(KEYINPUT13), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n235), .A2(KEYINPUT18), .A3(new_n237), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(G169gat), .B(G197gat), .Z(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G141gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n250), .B(KEYINPUT12), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n251), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n240), .A2(new_n253), .A3(new_n243), .A4(new_n244), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT72), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT26), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n258), .A2(G169gat), .A3(G176gat), .ZN(new_n259));
  INV_X1    g058(.A(G169gat), .ZN(new_n260));
  INV_X1    g059(.A(G176gat), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT66), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(KEYINPUT68), .B(new_n257), .C1(new_n259), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT66), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n258), .B1(G169gat), .B2(G176gat), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT26), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n269));
  INV_X1    g068(.A(new_n265), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n269), .B1(new_n270), .B2(KEYINPUT26), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n263), .B(new_n264), .C1(new_n268), .C2(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G190gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT28), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT67), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n281), .B(new_n276), .C1(new_n273), .C2(new_n274), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n278), .A2(KEYINPUT28), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n283), .A2(new_n284), .B1(G183gat), .B2(G190gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n272), .A2(new_n279), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n290), .A2(KEYINPUT65), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n265), .A2(KEYINPUT23), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n294), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n264), .A2(KEYINPUT23), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n293), .B(new_n295), .C1(new_n296), .C2(new_n265), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n287), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n296), .A2(new_n265), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT23), .B1(new_n259), .B2(new_n262), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n290), .A2(new_n291), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT25), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G120gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G113gat), .ZN(new_n306));
  INV_X1    g105(.A(G113gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G120gat), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT1), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G127gat), .A2(G134gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(G127gat), .A2(G134gat), .ZN(new_n312));
  NOR3_X1   g111(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT70), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT70), .ZN(new_n314));
  INV_X1    g113(.A(G127gat), .ZN(new_n315));
  INV_X1    g114(.A(G134gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n314), .B1(new_n317), .B2(new_n310), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n309), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT69), .B1(new_n311), .B2(new_n312), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n317), .A2(new_n321), .A3(new_n310), .ZN(new_n322));
  XNOR2_X1  g121(.A(G113gat), .B(G120gat), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n320), .B(new_n322), .C1(KEYINPUT1), .C2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n304), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n319), .A2(new_n324), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n286), .A2(new_n303), .A3(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n326), .A2(G227gat), .A3(G233gat), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT32), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT33), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G15gat), .B(G43gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(G71gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(G99gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n330), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n329), .B(KEYINPUT32), .C1(new_n331), .C2(new_n335), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n326), .A2(new_n328), .ZN(new_n341));
  NAND2_X1  g140(.A1(G227gat), .A2(G233gat), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT34), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n286), .A2(new_n303), .A3(new_n327), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n327), .B1(new_n286), .B2(new_n303), .ZN(new_n345));
  OAI211_X1 g144(.A(KEYINPUT34), .B(new_n342), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n340), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT34), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(KEYINPUT71), .A3(new_n346), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n256), .B1(new_n339), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n346), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n337), .A2(new_n338), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n338), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n358), .A2(KEYINPUT72), .A3(new_n348), .A4(new_n352), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n354), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT36), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n355), .B1(new_n337), .B2(new_n338), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n356), .A2(new_n362), .A3(KEYINPUT36), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G8gat), .B(G36gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(G64gat), .B(G92gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT73), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n286), .A2(new_n303), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n370), .B1(new_n286), .B2(new_n303), .ZN(new_n372));
  INV_X1    g171(.A(G226gat), .ZN(new_n373));
  INV_X1    g172(.A(G233gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n371), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G197gat), .B(G204gat), .ZN(new_n378));
  AND2_X1   g177(.A1(G211gat), .A2(G218gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n378), .B1(KEYINPUT22), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G211gat), .B(G218gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n375), .A2(KEYINPUT29), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n304), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n377), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n382), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n383), .B1(new_n371), .B2(new_n372), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n286), .A2(new_n303), .A3(new_n375), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n369), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n372), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n286), .A2(new_n303), .A3(new_n370), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n375), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(new_n387), .A3(new_n384), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n388), .A2(new_n389), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n395), .B(new_n368), .C1(new_n396), .C2(new_n387), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n391), .A2(new_n397), .A3(KEYINPUT30), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT30), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n399), .B(new_n369), .C1(new_n386), .C2(new_n390), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n402));
  XNOR2_X1  g201(.A(G57gat), .B(G85gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G1gat), .B(G29gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(KEYINPUT75), .ZN(new_n407));
  INV_X1    g206(.A(G141gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n408), .A2(G148gat), .ZN(new_n409));
  INV_X1    g208(.A(G148gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n410), .A2(G141gat), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n407), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413));
  INV_X1    g212(.A(G155gat), .ZN(new_n414));
  INV_X1    g213(.A(G162gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n413), .B1(new_n416), .B2(KEYINPUT2), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n410), .A2(G141gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n408), .A2(G148gat), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT75), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n412), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT2), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT74), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT74), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT2), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G141gat), .B(G148gat), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n413), .B(new_n416), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT3), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n421), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT76), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n421), .A2(new_n428), .A3(KEYINPUT76), .A4(new_n429), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n325), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n421), .A2(new_n428), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT3), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT75), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT75), .B1(new_n418), .B2(new_n419), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n413), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n418), .A2(new_n419), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT74), .B(KEYINPUT2), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n440), .A2(new_n417), .B1(new_n444), .B2(new_n416), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT77), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n325), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT77), .B1(new_n327), .B2(new_n435), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT4), .ZN(new_n449));
  NAND2_X1  g248(.A1(G225gat), .A2(G233gat), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n447), .B(new_n448), .C1(new_n449), .C2(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n327), .A2(new_n435), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT4), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n437), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n447), .B(new_n448), .C1(new_n445), .C2(new_n325), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n451), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(KEYINPUT5), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n447), .A2(KEYINPUT4), .A3(new_n448), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT79), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n453), .B2(new_n449), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n459), .A2(new_n461), .B1(new_n434), .B2(new_n436), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT5), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n460), .A4(KEYINPUT4), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n462), .A2(new_n463), .A3(new_n450), .A4(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT80), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n465), .A2(new_n466), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n406), .B(new_n458), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n458), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n459), .A2(new_n461), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(new_n437), .A3(new_n464), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n475), .A2(KEYINPUT80), .A3(new_n463), .A4(new_n450), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n465), .A2(new_n466), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(new_n406), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n478), .A2(new_n470), .A3(new_n406), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n401), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT81), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n429), .B1(new_n382), .B2(KEYINPUT29), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n435), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT29), .B1(new_n432), .B2(new_n433), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n486), .B1(new_n387), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(G228gat), .A2(G233gat), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n488), .A2(new_n490), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G22gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT83), .ZN(new_n495));
  INV_X1    g294(.A(G22gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(new_n496), .A3(new_n492), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G78gat), .B(G106gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT31), .B(G50gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n493), .A2(KEYINPUT83), .A3(G22gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n496), .B1(new_n491), .B2(new_n492), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n497), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n501), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n491), .A2(KEYINPUT82), .A3(new_n496), .A4(new_n492), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n458), .B1(new_n467), .B2(new_n468), .ZN(new_n511));
  INV_X1    g310(.A(new_n406), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(new_n470), .A3(new_n469), .ZN(new_n514));
  INV_X1    g313(.A(new_n481), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(KEYINPUT81), .A3(new_n401), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n484), .A2(new_n510), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n510), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT84), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n401), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n398), .A2(KEYINPUT84), .A3(new_n400), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT39), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n474), .A2(KEYINPUT85), .A3(new_n451), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT85), .B1(new_n474), .B2(new_n451), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n526), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n456), .A2(new_n451), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(new_n523), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n524), .A3(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n527), .A2(new_n531), .A3(KEYINPUT40), .A4(new_n406), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n521), .A2(new_n522), .A3(new_n532), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n527), .A2(new_n531), .A3(new_n406), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n513), .B1(new_n534), .B2(KEYINPUT40), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n391), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT37), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(new_n386), .B2(new_n390), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n382), .B1(new_n377), .B2(new_n385), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n388), .A2(new_n387), .A3(new_n389), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(KEYINPUT37), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(new_n542), .A3(new_n368), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT38), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n395), .B(KEYINPUT37), .C1(new_n396), .C2(new_n387), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n539), .A2(new_n546), .A3(KEYINPUT38), .A4(new_n368), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n537), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n548), .A2(new_n514), .A3(new_n515), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n519), .B1(new_n536), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n365), .B1(new_n518), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n356), .A2(new_n362), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n510), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT35), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n521), .A2(new_n522), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n554), .A2(new_n516), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n510), .A2(new_n360), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n484), .A2(new_n517), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n558), .B1(new_n560), .B2(KEYINPUT35), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n255), .B1(new_n551), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT92), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G127gat), .B(G155gat), .Z(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT20), .ZN(new_n566));
  XOR2_X1   g365(.A(G183gat), .B(G211gat), .Z(new_n567));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n566), .B(new_n569), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT21), .ZN(new_n572));
  XNOR2_X1  g371(.A(G57gat), .B(G64gat), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G71gat), .B(G78gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  OAI21_X1  g376(.A(new_n212), .B1(new_n572), .B2(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n578), .A2(KEYINPUT94), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(KEYINPUT94), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT93), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT93), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n579), .A2(new_n583), .A3(new_n580), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n584), .A3(KEYINPUT19), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT19), .B1(new_n582), .B2(new_n584), .ZN(new_n587));
  INV_X1    g386(.A(new_n577), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n588), .A2(KEYINPUT21), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n582), .A2(new_n584), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT19), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n591), .B1(new_n594), .B2(new_n585), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n571), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n589), .B1(new_n586), .B2(new_n587), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n594), .A2(new_n591), .A3(new_n585), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n598), .A3(new_n570), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G99gat), .B(G106gat), .Z(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n601), .A2(KEYINPUT95), .B1(KEYINPUT8), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT7), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n603), .B(new_n605), .C1(G85gat), .C2(G92gat), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n601), .A2(KEYINPUT95), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n234), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n608), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n229), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G190gat), .B(G218gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G134gat), .B(G162gat), .Z(new_n617));
  AOI21_X1  g416(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n616), .B(new_n619), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n564), .A2(new_n600), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n612), .B(new_n577), .ZN(new_n624));
  XOR2_X1   g423(.A(KEYINPUT96), .B(KEYINPUT10), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n612), .A2(KEYINPUT10), .A3(new_n588), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n624), .A2(new_n622), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(G176gat), .B(G204gat), .Z(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n630), .A2(KEYINPUT97), .A3(new_n633), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT97), .B1(new_n630), .B2(new_n633), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n621), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n516), .B(KEYINPUT98), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n207), .ZN(G1324gat));
  INV_X1    g443(.A(new_n556), .ZN(new_n645));
  INV_X1    g444(.A(G8gat), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n203), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n621), .A2(new_n639), .A3(new_n645), .A4(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n203), .A2(new_n646), .ZN(new_n650));
  OR3_X1    g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(G8gat), .B1(new_n640), .B2(new_n556), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n649), .B1(new_n648), .B2(new_n650), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(G1325gat));
  INV_X1    g453(.A(new_n640), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n656), .B1(new_n361), .B2(new_n364), .ZN(new_n657));
  AOI211_X1 g456(.A(KEYINPUT99), .B(new_n363), .C1(new_n360), .C2(KEYINPUT36), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n655), .A2(G15gat), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(G15gat), .B1(new_n655), .B2(new_n552), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(G1326gat));
  NOR2_X1   g461(.A1(new_n640), .A2(new_n519), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT43), .B(G22gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  INV_X1    g464(.A(new_n620), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n600), .A2(new_n638), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n564), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(new_n221), .A3(new_n641), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n669), .A2(KEYINPUT45), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(KEYINPUT45), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n659), .B1(new_n518), .B2(new_n550), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n666), .B1(new_n561), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI211_X1 g474(.A(KEYINPUT44), .B(new_n666), .C1(new_n551), .C2(new_n561), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n675), .A2(new_n255), .A3(new_n667), .A4(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n677), .A2(new_n642), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT100), .ZN(new_n679));
  OAI22_X1  g478(.A1(new_n670), .A2(new_n671), .B1(new_n221), .B2(new_n679), .ZN(G1328gat));
  NAND3_X1  g479(.A1(new_n668), .A2(new_n222), .A3(new_n645), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT46), .ZN(new_n682));
  OAI21_X1  g481(.A(G36gat), .B1(new_n677), .B2(new_n556), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n668), .A2(new_n222), .A3(new_n645), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n681), .A2(KEYINPUT101), .A3(KEYINPUT46), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n682), .B(new_n683), .C1(new_n687), .C2(new_n688), .ZN(G1329gat));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n553), .A2(G43gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n668), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n659), .ZN(new_n693));
  OAI21_X1  g492(.A(G43gat), .B1(new_n677), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n690), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1330gat));
  NAND3_X1  g496(.A1(new_n668), .A2(new_n215), .A3(new_n510), .ZN(new_n698));
  OAI21_X1  g497(.A(G50gat), .B1(new_n677), .B2(new_n519), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT48), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1331gat));
  INV_X1    g501(.A(new_n561), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n518), .A2(new_n550), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n693), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n639), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n600), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n707), .A2(new_n255), .A3(new_n666), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n641), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n710), .A2(new_n645), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT103), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1333gat));
  OAI21_X1  g516(.A(G71gat), .B1(new_n709), .B2(new_n693), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n552), .B(KEYINPUT104), .ZN(new_n719));
  INV_X1    g518(.A(G71gat), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n718), .B1(new_n709), .B2(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g522(.A1(new_n710), .A2(new_n510), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g524(.A1(new_n600), .A2(new_n639), .A3(new_n255), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n675), .A2(new_n676), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(G85gat), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n727), .A2(new_n728), .A3(new_n642), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n600), .A2(new_n255), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n666), .B(new_n730), .C1(new_n561), .C2(new_n672), .ZN(new_n731));
  NOR2_X1   g530(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n639), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n731), .A2(KEYINPUT105), .A3(KEYINPUT51), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n641), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n729), .B1(new_n738), .B2(new_n728), .ZN(G1336gat));
  NOR2_X1   g538(.A1(new_n556), .A2(G92gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742));
  OAI21_X1  g541(.A(G92gat), .B1(new_n727), .B2(new_n556), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n703), .A2(new_n705), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(KEYINPUT51), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n747), .A2(new_n666), .A3(new_n730), .A4(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n749), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n731), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n752), .A3(new_n638), .ZN(new_n753));
  INV_X1    g552(.A(new_n740), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n743), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT52), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n741), .A2(KEYINPUT107), .A3(new_n742), .A4(new_n743), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n746), .A2(new_n756), .A3(new_n757), .ZN(G1337gat));
  INV_X1    g557(.A(G99gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n737), .A2(new_n759), .A3(new_n552), .ZN(new_n760));
  OAI21_X1  g559(.A(G99gat), .B1(new_n727), .B2(new_n693), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(G1338gat));
  AOI21_X1  g561(.A(new_n620), .B1(new_n703), .B2(new_n705), .ZN(new_n763));
  INV_X1    g562(.A(new_n732), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n763), .A2(new_n730), .A3(new_n734), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n519), .A2(G106gat), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n765), .A2(new_n736), .A3(new_n638), .A4(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n735), .A2(KEYINPUT109), .A3(new_n736), .A4(new_n766), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n675), .A2(new_n510), .A3(new_n676), .A4(new_n726), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G106gat), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n769), .A2(new_n770), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n772), .A2(new_n775), .A3(G106gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n772), .B2(G106gat), .ZN(new_n777));
  AND4_X1   g576(.A1(new_n638), .A2(new_n750), .A3(new_n752), .A4(new_n766), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n774), .B1(new_n779), .B2(new_n771), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT110), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n774), .B(new_n782), .C1(new_n779), .C2(new_n771), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1339gat));
  INV_X1    g583(.A(new_n628), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n626), .A2(new_n623), .A3(new_n627), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(KEYINPUT54), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n633), .B1(new_n628), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n629), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n785), .A2(new_n791), .A3(new_n633), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT97), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n790), .A2(KEYINPUT55), .B1(new_n794), .B2(new_n635), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n235), .A2(new_n237), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n241), .A2(new_n242), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n250), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n254), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n787), .A2(new_n789), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n666), .A2(new_n795), .A3(new_n799), .A4(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n795), .A2(new_n255), .A3(new_n802), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n638), .A2(new_n799), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n620), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n805), .B1(new_n804), .B2(new_n806), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n803), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n707), .ZN(new_n811));
  INV_X1    g610(.A(new_n255), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n600), .A2(new_n639), .A3(new_n812), .A4(new_n620), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT111), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n642), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(new_n556), .A3(new_n554), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(new_n307), .A3(new_n812), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(new_n556), .A3(new_n559), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n819), .A2(new_n812), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n818), .B1(new_n307), .B2(new_n820), .ZN(G1340gat));
  OAI21_X1  g620(.A(G120gat), .B1(new_n817), .B2(new_n639), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n638), .A2(new_n305), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n819), .B2(new_n823), .ZN(G1341gat));
  OAI21_X1  g623(.A(G127gat), .B1(new_n817), .B2(new_n707), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n600), .A2(new_n315), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n819), .B2(new_n826), .ZN(G1342gat));
  OR2_X1    g626(.A1(new_n817), .A2(new_n620), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n828), .A2(new_n829), .A3(G134gat), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n828), .B2(G134gat), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n819), .A2(new_n620), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n832), .A2(KEYINPUT56), .A3(new_n316), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT56), .B1(new_n832), .B2(new_n316), .ZN(new_n834));
  OAI22_X1  g633(.A1(new_n830), .A2(new_n831), .B1(new_n833), .B2(new_n834), .ZN(G1343gat));
  NAND2_X1  g634(.A1(new_n693), .A2(new_n510), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n693), .A2(KEYINPUT117), .A3(new_n510), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n816), .A2(KEYINPUT118), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n794), .A2(new_n635), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n789), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n802), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n806), .B1(new_n844), .B2(new_n812), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT112), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n620), .A3(new_n807), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n600), .B1(new_n847), .B2(new_n803), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n641), .B(new_n839), .C1(new_n848), .C2(new_n814), .ZN(new_n849));
  INV_X1    g648(.A(new_n838), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n841), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n840), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n852), .A2(new_n408), .A3(new_n556), .A4(new_n255), .ZN(new_n853));
  XNOR2_X1  g652(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n252), .A2(new_n254), .B1(new_n800), .B2(new_n854), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n795), .A2(new_n855), .B1(new_n638), .B2(new_n799), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(KEYINPUT115), .A3(new_n620), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n856), .B2(new_n666), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n860), .A3(new_n803), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n814), .B1(new_n861), .B2(new_n707), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT57), .B1(new_n862), .B2(new_n519), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n864), .B(new_n510), .C1(new_n848), .C2(new_n814), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n642), .A2(new_n645), .A3(new_n659), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n863), .A2(new_n255), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT58), .B1(new_n867), .B2(G141gat), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n867), .A2(KEYINPUT116), .A3(G141gat), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n816), .A2(new_n838), .A3(new_n839), .ZN(new_n871));
  NOR4_X1   g670(.A1(new_n871), .A2(G141gat), .A3(new_n645), .A4(new_n812), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT116), .B1(new_n867), .B2(G141gat), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n869), .B1(new_n874), .B2(new_n875), .ZN(G1344gat));
  AND2_X1   g675(.A1(new_n852), .A2(new_n556), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n410), .A3(new_n638), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n638), .A3(new_n865), .A4(new_n866), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n880), .A3(G148gat), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n881), .B(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n519), .B1(new_n811), .B2(new_n815), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n803), .B1(new_n856), .B2(new_n666), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n886), .A2(new_n707), .B1(new_n708), .B2(new_n639), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n864), .B1(new_n887), .B2(new_n519), .ZN(new_n888));
  OAI211_X1 g687(.A(KEYINPUT57), .B(new_n510), .C1(new_n848), .C2(new_n814), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n885), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n638), .A3(new_n866), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n880), .B1(new_n893), .B2(G148gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n878), .B1(new_n883), .B2(new_n894), .ZN(G1345gat));
  NAND3_X1  g694(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n896), .A2(new_n414), .A3(new_n707), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n840), .A2(new_n851), .A3(new_n556), .A4(new_n600), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n898), .B(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n897), .B1(new_n900), .B2(new_n414), .ZN(G1346gat));
  NAND3_X1  g700(.A1(new_n877), .A2(new_n415), .A3(new_n666), .ZN(new_n902));
  OAI21_X1  g701(.A(G162gat), .B1(new_n896), .B2(new_n620), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1347gat));
  NAND2_X1  g703(.A1(new_n811), .A2(new_n815), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n641), .A2(new_n556), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n559), .A3(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n260), .A3(new_n255), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n906), .A2(new_n719), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n510), .B1(new_n910), .B2(KEYINPUT122), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n905), .B(new_n911), .C1(KEYINPUT122), .C2(new_n910), .ZN(new_n912));
  OAI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n812), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n909), .A2(new_n913), .ZN(G1348gat));
  AOI21_X1  g713(.A(G176gat), .B1(new_n908), .B2(new_n638), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n912), .A2(new_n261), .A3(new_n639), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(G1349gat));
  NAND3_X1  g716(.A1(new_n908), .A2(new_n275), .A3(new_n600), .ZN(new_n918));
  OAI21_X1  g717(.A(G183gat), .B1(new_n912), .B2(new_n707), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n921));
  AOI22_X1  g720(.A1(new_n918), .A2(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(G1350gat));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n276), .A3(new_n666), .ZN(new_n925));
  OAI21_X1  g724(.A(G190gat), .B1(new_n912), .B2(new_n620), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT124), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n929), .B(G190gat), .C1(new_n912), .C2(new_n620), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n928), .B1(new_n927), .B2(new_n930), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n925), .B1(new_n931), .B2(new_n932), .ZN(G1351gat));
  XOR2_X1   g732(.A(KEYINPUT125), .B(G197gat), .Z(new_n934));
  NOR3_X1   g733(.A1(new_n659), .A2(new_n641), .A3(new_n556), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT126), .Z(new_n936));
  NAND2_X1  g735(.A1(new_n892), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n937), .B2(new_n812), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n884), .A2(new_n935), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n812), .A2(new_n934), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(G1352gat));
  OR3_X1    g740(.A1(new_n939), .A2(G204gat), .A3(new_n639), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n942), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n892), .A2(new_n638), .A3(new_n936), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G204gat), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n942), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(G1353gat));
  OR3_X1    g749(.A1(new_n939), .A2(G211gat), .A3(new_n707), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n892), .A2(new_n600), .A3(new_n936), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n952), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(G1354gat));
  OAI21_X1  g754(.A(G218gat), .B1(new_n937), .B2(new_n620), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n620), .A2(G218gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n939), .B2(new_n957), .ZN(G1355gat));
endmodule


