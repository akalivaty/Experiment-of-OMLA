

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U551 ( .A1(n536), .A2(G2104), .ZN(n881) );
  NOR2_X1 U552 ( .A1(G2084), .A2(n724), .ZN(n712) );
  NOR2_X1 U553 ( .A1(G1966), .A2(n798), .ZN(n739) );
  NOR2_X1 U554 ( .A1(n713), .A2(n739), .ZN(n714) );
  INV_X1 U555 ( .A(KEYINPUT31), .ZN(n720) );
  XNOR2_X1 U556 ( .A(n721), .B(n720), .ZN(n722) );
  INV_X1 U557 ( .A(KEYINPUT96), .ZN(n679) );
  INV_X1 U558 ( .A(KEYINPUT89), .ZN(n677) );
  XNOR2_X1 U559 ( .A(n678), .B(n677), .ZN(n761) );
  NOR2_X1 U560 ( .A1(G651), .A2(n615), .ZN(n630) );
  XNOR2_X1 U561 ( .A(G543), .B(KEYINPUT0), .ZN(n517) );
  XNOR2_X1 U562 ( .A(n517), .B(KEYINPUT65), .ZN(n615) );
  NAND2_X1 U563 ( .A1(n630), .A2(G51), .ZN(n521) );
  INV_X1 U564 ( .A(G651), .ZN(n524) );
  NOR2_X1 U565 ( .A1(G543), .A2(n524), .ZN(n518) );
  XOR2_X1 U566 ( .A(KEYINPUT66), .B(n518), .Z(n519) );
  XNOR2_X1 U567 ( .A(KEYINPUT1), .B(n519), .ZN(n632) );
  NAND2_X1 U568 ( .A1(G63), .A2(n632), .ZN(n520) );
  NAND2_X1 U569 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U570 ( .A(KEYINPUT6), .B(n522), .ZN(n529) );
  NOR2_X1 U571 ( .A1(G651), .A2(G543), .ZN(n636) );
  NAND2_X1 U572 ( .A1(n636), .A2(G89), .ZN(n523) );
  XNOR2_X1 U573 ( .A(n523), .B(KEYINPUT4), .ZN(n526) );
  NOR2_X1 U574 ( .A1(n615), .A2(n524), .ZN(n637) );
  NAND2_X1 U575 ( .A1(G76), .A2(n637), .ZN(n525) );
  NAND2_X1 U576 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U577 ( .A(n527), .B(KEYINPUT5), .Z(n528) );
  NOR2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U579 ( .A(KEYINPUT7), .B(n530), .Z(n531) );
  XNOR2_X1 U580 ( .A(KEYINPUT74), .B(n531), .ZN(G168) );
  XOR2_X1 U581 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  INV_X1 U582 ( .A(G2105), .ZN(n536) );
  AND2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n874) );
  NAND2_X1 U584 ( .A1(n874), .A2(G113), .ZN(n534) );
  NAND2_X1 U585 ( .A1(G101), .A2(n881), .ZN(n532) );
  XOR2_X1 U586 ( .A(KEYINPUT23), .B(n532), .Z(n533) );
  NAND2_X1 U587 ( .A1(n534), .A2(n533), .ZN(n540) );
  NOR2_X1 U588 ( .A1(G2104), .A2(G2105), .ZN(n535) );
  XOR2_X2 U589 ( .A(KEYINPUT17), .B(n535), .Z(n882) );
  NAND2_X1 U590 ( .A1(G137), .A2(n882), .ZN(n538) );
  NOR2_X1 U591 ( .A1(G2104), .A2(n536), .ZN(n875) );
  NAND2_X1 U592 ( .A1(G125), .A2(n875), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U594 ( .A1(n540), .A2(n539), .ZN(G160) );
  NAND2_X1 U595 ( .A1(n630), .A2(G52), .ZN(n542) );
  NAND2_X1 U596 ( .A1(G64), .A2(n632), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n547) );
  NAND2_X1 U598 ( .A1(G90), .A2(n636), .ZN(n544) );
  NAND2_X1 U599 ( .A1(G77), .A2(n637), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U601 ( .A(KEYINPUT9), .B(n545), .Z(n546) );
  NOR2_X1 U602 ( .A1(n547), .A2(n546), .ZN(G171) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U604 ( .A(G57), .ZN(G237) );
  INV_X1 U605 ( .A(G132), .ZN(G219) );
  INV_X1 U606 ( .A(G82), .ZN(G220) );
  NAND2_X1 U607 ( .A1(G7), .A2(G661), .ZN(n548) );
  XNOR2_X1 U608 ( .A(n548), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U609 ( .A(G223), .ZN(n829) );
  NAND2_X1 U610 ( .A1(n829), .A2(G567), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT11), .B(n549), .Z(G234) );
  NAND2_X1 U612 ( .A1(n632), .A2(G56), .ZN(n551) );
  XNOR2_X1 U613 ( .A(KEYINPUT14), .B(KEYINPUT71), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(n557) );
  NAND2_X1 U615 ( .A1(n636), .A2(G81), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n552), .B(KEYINPUT12), .ZN(n554) );
  NAND2_X1 U617 ( .A1(G68), .A2(n637), .ZN(n553) );
  NAND2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U619 ( .A(KEYINPUT13), .B(n555), .Z(n556) );
  NOR2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n630), .A2(G43), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n977) );
  INV_X1 U623 ( .A(G860), .ZN(n581) );
  NOR2_X1 U624 ( .A1(n977), .A2(n581), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT72), .B(n560), .Z(G153) );
  INV_X1 U626 ( .A(G171), .ZN(G301) );
  NAND2_X1 U627 ( .A1(G868), .A2(G301), .ZN(n570) );
  NAND2_X1 U628 ( .A1(G92), .A2(n636), .ZN(n562) );
  NAND2_X1 U629 ( .A1(G66), .A2(n632), .ZN(n561) );
  NAND2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n567) );
  NAND2_X1 U631 ( .A1(G79), .A2(n637), .ZN(n564) );
  NAND2_X1 U632 ( .A1(G54), .A2(n630), .ZN(n563) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U634 ( .A(KEYINPUT73), .B(n565), .Z(n566) );
  NOR2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U636 ( .A(KEYINPUT15), .B(n568), .ZN(n987) );
  INV_X1 U637 ( .A(G868), .ZN(n653) );
  NAND2_X1 U638 ( .A1(n987), .A2(n653), .ZN(n569) );
  NAND2_X1 U639 ( .A1(n570), .A2(n569), .ZN(G284) );
  NAND2_X1 U640 ( .A1(G65), .A2(n632), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G91), .A2(n636), .ZN(n572) );
  NAND2_X1 U642 ( .A1(G78), .A2(n637), .ZN(n571) );
  NAND2_X1 U643 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U644 ( .A1(G53), .A2(n630), .ZN(n573) );
  XNOR2_X1 U645 ( .A(KEYINPUT69), .B(n573), .ZN(n574) );
  NOR2_X1 U646 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U647 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U648 ( .A(n578), .B(KEYINPUT70), .ZN(G299) );
  NAND2_X1 U649 ( .A1(G868), .A2(G286), .ZN(n580) );
  NAND2_X1 U650 ( .A1(G299), .A2(n653), .ZN(n579) );
  NAND2_X1 U651 ( .A1(n580), .A2(n579), .ZN(G297) );
  NAND2_X1 U652 ( .A1(n581), .A2(G559), .ZN(n582) );
  INV_X1 U653 ( .A(n987), .ZN(n899) );
  NAND2_X1 U654 ( .A1(n582), .A2(n899), .ZN(n583) );
  XNOR2_X1 U655 ( .A(n583), .B(KEYINPUT16), .ZN(n584) );
  XOR2_X1 U656 ( .A(KEYINPUT75), .B(n584), .Z(G148) );
  NAND2_X1 U657 ( .A1(n899), .A2(G868), .ZN(n585) );
  NOR2_X1 U658 ( .A1(G559), .A2(n585), .ZN(n586) );
  XOR2_X1 U659 ( .A(KEYINPUT77), .B(n586), .Z(n589) );
  NOR2_X1 U660 ( .A1(G868), .A2(n977), .ZN(n587) );
  XNOR2_X1 U661 ( .A(KEYINPUT76), .B(n587), .ZN(n588) );
  NOR2_X1 U662 ( .A1(n589), .A2(n588), .ZN(G282) );
  NAND2_X1 U663 ( .A1(G99), .A2(n881), .ZN(n591) );
  NAND2_X1 U664 ( .A1(G111), .A2(n874), .ZN(n590) );
  NAND2_X1 U665 ( .A1(n591), .A2(n590), .ZN(n597) );
  NAND2_X1 U666 ( .A1(G123), .A2(n875), .ZN(n592) );
  XNOR2_X1 U667 ( .A(n592), .B(KEYINPUT18), .ZN(n595) );
  NAND2_X1 U668 ( .A1(G135), .A2(n882), .ZN(n593) );
  XNOR2_X1 U669 ( .A(n593), .B(KEYINPUT78), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n960) );
  XNOR2_X1 U672 ( .A(n960), .B(G2096), .ZN(n599) );
  INV_X1 U673 ( .A(G2100), .ZN(n598) );
  NAND2_X1 U674 ( .A1(n599), .A2(n598), .ZN(G156) );
  NAND2_X1 U675 ( .A1(G93), .A2(n636), .ZN(n601) );
  NAND2_X1 U676 ( .A1(G80), .A2(n637), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U678 ( .A1(G67), .A2(n632), .ZN(n602) );
  XNOR2_X1 U679 ( .A(KEYINPUT79), .B(n602), .ZN(n603) );
  NOR2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n630), .A2(G55), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n652) );
  NAND2_X1 U683 ( .A1(G559), .A2(n899), .ZN(n607) );
  XNOR2_X1 U684 ( .A(n607), .B(n977), .ZN(n650) );
  NOR2_X1 U685 ( .A1(G860), .A2(n650), .ZN(n608) );
  XOR2_X1 U686 ( .A(n652), .B(n608), .Z(G145) );
  NAND2_X1 U687 ( .A1(G88), .A2(n636), .ZN(n610) );
  NAND2_X1 U688 ( .A1(G75), .A2(n637), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n630), .A2(G50), .ZN(n612) );
  NAND2_X1 U691 ( .A1(G62), .A2(n632), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U693 ( .A1(n614), .A2(n613), .ZN(G166) );
  NAND2_X1 U694 ( .A1(G87), .A2(n615), .ZN(n617) );
  NAND2_X1 U695 ( .A1(G74), .A2(G651), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U697 ( .A1(n632), .A2(n618), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n630), .A2(G49), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(G288) );
  XOR2_X1 U700 ( .A(KEYINPUT80), .B(KEYINPUT2), .Z(n622) );
  NAND2_X1 U701 ( .A1(G73), .A2(n637), .ZN(n621) );
  XNOR2_X1 U702 ( .A(n622), .B(n621), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G86), .A2(n636), .ZN(n624) );
  NAND2_X1 U704 ( .A1(G61), .A2(n632), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U707 ( .A(KEYINPUT81), .B(n627), .Z(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(G48), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(G305) );
  NAND2_X1 U710 ( .A1(n630), .A2(G47), .ZN(n631) );
  XOR2_X1 U711 ( .A(KEYINPUT67), .B(n631), .Z(n634) );
  NAND2_X1 U712 ( .A1(G60), .A2(n632), .ZN(n633) );
  NAND2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U714 ( .A(KEYINPUT68), .B(n635), .Z(n641) );
  NAND2_X1 U715 ( .A1(G85), .A2(n636), .ZN(n639) );
  NAND2_X1 U716 ( .A1(G72), .A2(n637), .ZN(n638) );
  AND2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(G290) );
  XOR2_X1 U719 ( .A(KEYINPUT19), .B(KEYINPUT83), .Z(n642) );
  XNOR2_X1 U720 ( .A(G288), .B(n642), .ZN(n643) );
  XOR2_X1 U721 ( .A(n643), .B(KEYINPUT84), .Z(n645) );
  XNOR2_X1 U722 ( .A(G299), .B(KEYINPUT82), .ZN(n644) );
  XNOR2_X1 U723 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U724 ( .A(G166), .B(n646), .ZN(n647) );
  XNOR2_X1 U725 ( .A(n647), .B(n652), .ZN(n649) );
  XOR2_X1 U726 ( .A(G305), .B(G290), .Z(n648) );
  XNOR2_X1 U727 ( .A(n649), .B(n648), .ZN(n898) );
  XNOR2_X1 U728 ( .A(n650), .B(n898), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n651), .A2(G868), .ZN(n655) );
  NAND2_X1 U730 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n655), .A2(n654), .ZN(G295) );
  NAND2_X1 U732 ( .A1(G2078), .A2(G2084), .ZN(n656) );
  XNOR2_X1 U733 ( .A(n656), .B(KEYINPUT85), .ZN(n657) );
  XNOR2_X1 U734 ( .A(n657), .B(KEYINPUT20), .ZN(n658) );
  NAND2_X1 U735 ( .A1(n658), .A2(G2090), .ZN(n659) );
  XNOR2_X1 U736 ( .A(KEYINPUT21), .B(n659), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n660), .A2(G2072), .ZN(n661) );
  XNOR2_X1 U738 ( .A(KEYINPUT86), .B(n661), .ZN(G158) );
  XNOR2_X1 U739 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U740 ( .A1(G220), .A2(G219), .ZN(n662) );
  XOR2_X1 U741 ( .A(KEYINPUT22), .B(n662), .Z(n663) );
  NOR2_X1 U742 ( .A1(G218), .A2(n663), .ZN(n664) );
  NAND2_X1 U743 ( .A1(G96), .A2(n664), .ZN(n833) );
  NAND2_X1 U744 ( .A1(n833), .A2(G2106), .ZN(n668) );
  NAND2_X1 U745 ( .A1(G69), .A2(G120), .ZN(n665) );
  NOR2_X1 U746 ( .A1(G237), .A2(n665), .ZN(n666) );
  NAND2_X1 U747 ( .A1(G108), .A2(n666), .ZN(n834) );
  NAND2_X1 U748 ( .A1(n834), .A2(G567), .ZN(n667) );
  NAND2_X1 U749 ( .A1(n668), .A2(n667), .ZN(n835) );
  NAND2_X1 U750 ( .A1(G483), .A2(G661), .ZN(n669) );
  NOR2_X1 U751 ( .A1(n835), .A2(n669), .ZN(n832) );
  NAND2_X1 U752 ( .A1(n832), .A2(G36), .ZN(G176) );
  NAND2_X1 U753 ( .A1(G102), .A2(n881), .ZN(n671) );
  NAND2_X1 U754 ( .A1(G138), .A2(n882), .ZN(n670) );
  NAND2_X1 U755 ( .A1(n671), .A2(n670), .ZN(n675) );
  NAND2_X1 U756 ( .A1(G114), .A2(n874), .ZN(n673) );
  NAND2_X1 U757 ( .A1(G126), .A2(n875), .ZN(n672) );
  NAND2_X1 U758 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U759 ( .A1(n675), .A2(n674), .ZN(G164) );
  XNOR2_X1 U760 ( .A(KEYINPUT87), .B(G166), .ZN(G303) );
  NOR2_X1 U761 ( .A1(G1976), .A2(G288), .ZN(n746) );
  NOR2_X1 U762 ( .A1(G1971), .A2(G303), .ZN(n676) );
  NOR2_X1 U763 ( .A1(n746), .A2(n676), .ZN(n993) );
  XNOR2_X1 U764 ( .A(KEYINPUT106), .B(n993), .ZN(n744) );
  NAND2_X1 U765 ( .A1(G160), .A2(G40), .ZN(n678) );
  XNOR2_X1 U766 ( .A(n761), .B(n679), .ZN(n680) );
  NOR2_X1 U767 ( .A1(G164), .A2(G1384), .ZN(n762) );
  NAND2_X1 U768 ( .A1(n680), .A2(n762), .ZN(n724) );
  NAND2_X1 U769 ( .A1(n724), .A2(G1961), .ZN(n682) );
  INV_X1 U770 ( .A(n724), .ZN(n694) );
  XOR2_X1 U771 ( .A(KEYINPUT25), .B(G2078), .Z(n1002) );
  NAND2_X1 U772 ( .A1(n694), .A2(n1002), .ZN(n681) );
  NAND2_X1 U773 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U774 ( .A(n683), .B(KEYINPUT98), .Z(n716) );
  NAND2_X1 U775 ( .A1(n716), .A2(G171), .ZN(n711) );
  NAND2_X1 U776 ( .A1(n694), .A2(G2072), .ZN(n684) );
  XNOR2_X1 U777 ( .A(n684), .B(KEYINPUT27), .ZN(n686) );
  AND2_X1 U778 ( .A1(G1956), .A2(n724), .ZN(n685) );
  NOR2_X1 U779 ( .A1(n686), .A2(n685), .ZN(n701) );
  INV_X1 U780 ( .A(G299), .ZN(n974) );
  NOR2_X1 U781 ( .A1(n701), .A2(n974), .ZN(n687) );
  XOR2_X1 U782 ( .A(n687), .B(KEYINPUT28), .Z(n707) );
  XOR2_X1 U783 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n689) );
  NAND2_X1 U784 ( .A1(G1996), .A2(n694), .ZN(n688) );
  XNOR2_X1 U785 ( .A(n689), .B(n688), .ZN(n692) );
  NAND2_X1 U786 ( .A1(G1341), .A2(n724), .ZN(n690) );
  XNOR2_X1 U787 ( .A(KEYINPUT99), .B(n690), .ZN(n691) );
  NOR2_X1 U788 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U789 ( .A(n693), .B(KEYINPUT100), .ZN(n699) );
  NAND2_X1 U790 ( .A1(G1348), .A2(n724), .ZN(n696) );
  NAND2_X1 U791 ( .A1(n694), .A2(G2067), .ZN(n695) );
  NAND2_X1 U792 ( .A1(n696), .A2(n695), .ZN(n700) );
  AND2_X1 U793 ( .A1(n700), .A2(n987), .ZN(n697) );
  NOR2_X1 U794 ( .A1(n697), .A2(n977), .ZN(n698) );
  NAND2_X1 U795 ( .A1(n699), .A2(n698), .ZN(n705) );
  NOR2_X1 U796 ( .A1(n987), .A2(n700), .ZN(n703) );
  AND2_X1 U797 ( .A1(n701), .A2(n974), .ZN(n702) );
  NOR2_X1 U798 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U799 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n707), .A2(n706), .ZN(n709) );
  XNOR2_X1 U801 ( .A(KEYINPUT101), .B(KEYINPUT29), .ZN(n708) );
  XNOR2_X1 U802 ( .A(n709), .B(n708), .ZN(n710) );
  NAND2_X1 U803 ( .A1(n711), .A2(n710), .ZN(n723) );
  XNOR2_X1 U804 ( .A(n712), .B(KEYINPUT97), .ZN(n735) );
  NAND2_X1 U805 ( .A1(G8), .A2(n735), .ZN(n713) );
  NAND2_X1 U806 ( .A1(G8), .A2(n724), .ZN(n798) );
  XOR2_X1 U807 ( .A(n714), .B(KEYINPUT30), .Z(n715) );
  OR2_X1 U808 ( .A1(G168), .A2(n715), .ZN(n719) );
  OR2_X1 U809 ( .A1(n716), .A2(G171), .ZN(n717) );
  XNOR2_X1 U810 ( .A(KEYINPUT102), .B(n717), .ZN(n718) );
  AND2_X1 U811 ( .A1(n719), .A2(n718), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n723), .A2(n722), .ZN(n737) );
  NAND2_X1 U813 ( .A1(n737), .A2(G286), .ZN(n731) );
  NOR2_X1 U814 ( .A1(G2090), .A2(n724), .ZN(n725) );
  XOR2_X1 U815 ( .A(KEYINPUT103), .B(n725), .Z(n727) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n798), .ZN(n726) );
  NOR2_X1 U817 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U818 ( .A1(n728), .A2(G303), .ZN(n729) );
  XNOR2_X1 U819 ( .A(n729), .B(KEYINPUT104), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U821 ( .A(KEYINPUT105), .B(n732), .Z(n733) );
  NAND2_X1 U822 ( .A1(G8), .A2(n733), .ZN(n734) );
  XNOR2_X1 U823 ( .A(n734), .B(KEYINPUT32), .ZN(n743) );
  INV_X1 U824 ( .A(n735), .ZN(n736) );
  NAND2_X1 U825 ( .A1(G8), .A2(n736), .ZN(n741) );
  INV_X1 U826 ( .A(n737), .ZN(n738) );
  NOR2_X1 U827 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U828 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U829 ( .A1(n743), .A2(n742), .ZN(n797) );
  AND2_X1 U830 ( .A1(n744), .A2(n797), .ZN(n786) );
  NAND2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n990) );
  INV_X1 U832 ( .A(n798), .ZN(n745) );
  NAND2_X1 U833 ( .A1(n990), .A2(n745), .ZN(n784) );
  NAND2_X1 U834 ( .A1(n746), .A2(KEYINPUT33), .ZN(n747) );
  NOR2_X1 U835 ( .A1(n747), .A2(n798), .ZN(n782) );
  XNOR2_X1 U836 ( .A(G1981), .B(KEYINPUT107), .ZN(n748) );
  XNOR2_X1 U837 ( .A(n748), .B(G305), .ZN(n980) );
  XNOR2_X1 U838 ( .A(G2067), .B(KEYINPUT37), .ZN(n749) );
  XOR2_X1 U839 ( .A(n749), .B(KEYINPUT90), .Z(n813) );
  XNOR2_X1 U840 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n760) );
  NAND2_X1 U841 ( .A1(G104), .A2(n881), .ZN(n751) );
  NAND2_X1 U842 ( .A1(G140), .A2(n882), .ZN(n750) );
  NAND2_X1 U843 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U844 ( .A(KEYINPUT34), .B(n752), .ZN(n757) );
  NAND2_X1 U845 ( .A1(G116), .A2(n874), .ZN(n754) );
  NAND2_X1 U846 ( .A1(G128), .A2(n875), .ZN(n753) );
  NAND2_X1 U847 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U848 ( .A(n755), .B(KEYINPUT35), .Z(n756) );
  NOR2_X1 U849 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U850 ( .A(KEYINPUT36), .B(n758), .Z(n759) );
  XOR2_X1 U851 ( .A(n760), .B(n759), .Z(n894) );
  AND2_X1 U852 ( .A1(n813), .A2(n894), .ZN(n959) );
  NOR2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n824) );
  AND2_X1 U854 ( .A1(n959), .A2(n824), .ZN(n820) );
  XNOR2_X1 U855 ( .A(KEYINPUT94), .B(n824), .ZN(n779) );
  NAND2_X1 U856 ( .A1(G95), .A2(n881), .ZN(n764) );
  NAND2_X1 U857 ( .A1(G107), .A2(n874), .ZN(n763) );
  NAND2_X1 U858 ( .A1(n764), .A2(n763), .ZN(n768) );
  NAND2_X1 U859 ( .A1(G131), .A2(n882), .ZN(n766) );
  NAND2_X1 U860 ( .A1(G119), .A2(n875), .ZN(n765) );
  NAND2_X1 U861 ( .A1(n766), .A2(n765), .ZN(n767) );
  OR2_X1 U862 ( .A1(n768), .A2(n767), .ZN(n887) );
  NAND2_X1 U863 ( .A1(G1991), .A2(n887), .ZN(n778) );
  NAND2_X1 U864 ( .A1(G105), .A2(n881), .ZN(n769) );
  XNOR2_X1 U865 ( .A(n769), .B(KEYINPUT38), .ZN(n776) );
  NAND2_X1 U866 ( .A1(G141), .A2(n882), .ZN(n771) );
  NAND2_X1 U867 ( .A1(G117), .A2(n874), .ZN(n770) );
  NAND2_X1 U868 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U869 ( .A1(G129), .A2(n875), .ZN(n772) );
  XNOR2_X1 U870 ( .A(KEYINPUT93), .B(n772), .ZN(n773) );
  NOR2_X1 U871 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U872 ( .A1(n776), .A2(n775), .ZN(n890) );
  NAND2_X1 U873 ( .A1(G1996), .A2(n890), .ZN(n777) );
  NAND2_X1 U874 ( .A1(n778), .A2(n777), .ZN(n967) );
  NAND2_X1 U875 ( .A1(n779), .A2(n967), .ZN(n780) );
  XNOR2_X1 U876 ( .A(KEYINPUT95), .B(n780), .ZN(n816) );
  NOR2_X1 U877 ( .A1(n820), .A2(n816), .ZN(n803) );
  NAND2_X1 U878 ( .A1(n980), .A2(n803), .ZN(n781) );
  NOR2_X1 U879 ( .A1(n782), .A2(n781), .ZN(n787) );
  INV_X1 U880 ( .A(n787), .ZN(n783) );
  OR2_X1 U881 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U882 ( .A1(n786), .A2(n785), .ZN(n789) );
  AND2_X1 U883 ( .A1(n787), .A2(KEYINPUT33), .ZN(n788) );
  NOR2_X1 U884 ( .A1(n789), .A2(n788), .ZN(n805) );
  NOR2_X1 U885 ( .A1(G2090), .A2(G303), .ZN(n790) );
  NAND2_X1 U886 ( .A1(G8), .A2(n790), .ZN(n791) );
  XNOR2_X1 U887 ( .A(n791), .B(KEYINPUT108), .ZN(n795) );
  NOR2_X1 U888 ( .A1(G1981), .A2(G305), .ZN(n792) );
  XOR2_X1 U889 ( .A(n792), .B(KEYINPUT24), .Z(n793) );
  NOR2_X1 U890 ( .A1(n798), .A2(n793), .ZN(n799) );
  INV_X1 U891 ( .A(n799), .ZN(n794) );
  AND2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n801) );
  OR2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n800) );
  AND2_X1 U895 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n805), .A2(n804), .ZN(n810) );
  XNOR2_X1 U898 ( .A(KEYINPUT88), .B(G1986), .ZN(n806) );
  XNOR2_X1 U899 ( .A(n806), .B(G290), .ZN(n984) );
  NAND2_X1 U900 ( .A1(n824), .A2(n984), .ZN(n807) );
  NAND2_X1 U901 ( .A1(n810), .A2(n807), .ZN(n809) );
  INV_X1 U902 ( .A(KEYINPUT109), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n812) );
  NAND2_X1 U904 ( .A1(n810), .A2(KEYINPUT109), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n827) );
  NAND2_X1 U906 ( .A1(n984), .A2(KEYINPUT109), .ZN(n823) );
  NOR2_X1 U907 ( .A1(n813), .A2(n894), .ZN(n963) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n890), .ZN(n954) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n814) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n887), .ZN(n961) );
  NOR2_X1 U911 ( .A1(n814), .A2(n961), .ZN(n815) );
  NOR2_X1 U912 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U913 ( .A1(n954), .A2(n817), .ZN(n818) );
  XOR2_X1 U914 ( .A(KEYINPUT39), .B(n818), .Z(n819) );
  NOR2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U916 ( .A1(n963), .A2(n821), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U920 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n829), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U923 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  INV_X1 U929 ( .A(G69), .ZN(G235) );
  NOR2_X1 U930 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  INV_X1 U932 ( .A(n835), .ZN(G319) );
  XNOR2_X1 U933 ( .A(G1996), .B(KEYINPUT41), .ZN(n845) );
  XOR2_X1 U934 ( .A(G1991), .B(G1971), .Z(n837) );
  XNOR2_X1 U935 ( .A(G1956), .B(G1961), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U937 ( .A(G1986), .B(G1976), .Z(n839) );
  XNOR2_X1 U938 ( .A(G1966), .B(G1981), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U940 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U941 ( .A(KEYINPUT114), .B(G2474), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(G229) );
  XOR2_X1 U944 ( .A(G2100), .B(G2096), .Z(n847) );
  XNOR2_X1 U945 ( .A(KEYINPUT42), .B(G2678), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT43), .B(G2090), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U950 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U951 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(G227) );
  NAND2_X1 U953 ( .A1(G124), .A2(n875), .ZN(n854) );
  XOR2_X1 U954 ( .A(KEYINPUT115), .B(n854), .Z(n855) );
  XNOR2_X1 U955 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U956 ( .A1(G112), .A2(n874), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U958 ( .A1(G100), .A2(n881), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G136), .A2(n882), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U961 ( .A1(n861), .A2(n860), .ZN(G162) );
  XOR2_X1 U962 ( .A(KEYINPUT117), .B(KEYINPUT46), .Z(n872) );
  NAND2_X1 U963 ( .A1(G118), .A2(n874), .ZN(n863) );
  NAND2_X1 U964 ( .A1(G130), .A2(n875), .ZN(n862) );
  NAND2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n869) );
  NAND2_X1 U966 ( .A1(G106), .A2(n881), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G142), .A2(n882), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U969 ( .A(KEYINPUT45), .B(n866), .Z(n867) );
  XNOR2_X1 U970 ( .A(KEYINPUT116), .B(n867), .ZN(n868) );
  NOR2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U972 ( .A(KEYINPUT48), .B(n870), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n960), .B(n873), .ZN(n889) );
  XNOR2_X1 U975 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n880) );
  NAND2_X1 U976 ( .A1(G115), .A2(n874), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G127), .A2(n875), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n878), .B(KEYINPUT47), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n886) );
  NAND2_X1 U981 ( .A1(G103), .A2(n881), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G139), .A2(n882), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n885) );
  NOR2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n947) );
  XNOR2_X1 U985 ( .A(n887), .B(n947), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n896) );
  XNOR2_X1 U987 ( .A(n890), .B(G162), .ZN(n892) );
  XNOR2_X1 U988 ( .A(G160), .B(G164), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U990 ( .A(n894), .B(n893), .Z(n895) );
  XNOR2_X1 U991 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U992 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U993 ( .A(G171), .B(n898), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n977), .B(n899), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U996 ( .A(n902), .B(G286), .Z(n903) );
  NOR2_X1 U997 ( .A1(G37), .A2(n903), .ZN(G397) );
  XOR2_X1 U998 ( .A(KEYINPUT112), .B(G2454), .Z(n905) );
  XNOR2_X1 U999 ( .A(G1348), .B(G1341), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n915) );
  XOR2_X1 U1001 ( .A(KEYINPUT113), .B(KEYINPUT110), .Z(n907) );
  XNOR2_X1 U1002 ( .A(G2427), .B(G2451), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U1004 ( .A(G2430), .B(G2443), .Z(n909) );
  XNOR2_X1 U1005 ( .A(G2438), .B(G2435), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1007 ( .A(n911), .B(n910), .Z(n913) );
  XNOR2_X1 U1008 ( .A(KEYINPUT111), .B(G2446), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n915), .B(n914), .ZN(n916) );
  NAND2_X1 U1011 ( .A1(n916), .A2(G14), .ZN(n922) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n922), .ZN(n919) );
  NOR2_X1 U1013 ( .A1(G229), .A2(G227), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G108), .ZN(G238) );
  INV_X1 U1020 ( .A(n922), .ZN(G401) );
  XNOR2_X1 U1021 ( .A(G1966), .B(G21), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(G5), .B(G1961), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n937) );
  XNOR2_X1 U1024 ( .A(KEYINPUT60), .B(KEYINPUT127), .ZN(n935) );
  XNOR2_X1 U1025 ( .A(KEYINPUT125), .B(G1956), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(n925), .B(G20), .ZN(n933) );
  XOR2_X1 U1027 ( .A(G1981), .B(G6), .Z(n928) );
  XOR2_X1 U1028 ( .A(G19), .B(KEYINPUT126), .Z(n926) );
  XNOR2_X1 U1029 ( .A(G1341), .B(n926), .ZN(n927) );
  NAND2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n931) );
  XOR2_X1 U1031 ( .A(KEYINPUT59), .B(G1348), .Z(n929) );
  XNOR2_X1 U1032 ( .A(G4), .B(n929), .ZN(n930) );
  NOR2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1035 ( .A(n935), .B(n934), .ZN(n936) );
  NAND2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(G1971), .B(G22), .ZN(n939) );
  XNOR2_X1 U1038 ( .A(G23), .B(G1976), .ZN(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n941) );
  XOR2_X1 U1040 ( .A(G1986), .B(G24), .Z(n940) );
  NAND2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(KEYINPUT58), .B(n942), .ZN(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1044 ( .A(KEYINPUT61), .B(n945), .Z(n946) );
  NOR2_X1 U1045 ( .A1(G16), .A2(n946), .ZN(n1025) );
  XNOR2_X1 U1046 ( .A(KEYINPUT55), .B(KEYINPUT123), .ZN(n1016) );
  XOR2_X1 U1047 ( .A(G2072), .B(n947), .Z(n948) );
  XNOR2_X1 U1048 ( .A(KEYINPUT120), .B(n948), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(G2078), .B(G164), .ZN(n949) );
  XNOR2_X1 U1050 ( .A(KEYINPUT121), .B(n949), .ZN(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(KEYINPUT50), .B(n952), .ZN(n957) );
  XOR2_X1 U1053 ( .A(G2090), .B(G162), .Z(n953) );
  NOR2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1055 ( .A(KEYINPUT51), .B(n955), .Z(n956) );
  NAND2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n969) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n965) );
  XOR2_X1 U1059 ( .A(G2084), .B(G160), .Z(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(KEYINPUT52), .B(n970), .ZN(n971) );
  XOR2_X1 U1065 ( .A(KEYINPUT122), .B(n971), .Z(n972) );
  NAND2_X1 U1066 ( .A1(n1016), .A2(n972), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n973), .A2(G29), .ZN(n1023) );
  XOR2_X1 U1068 ( .A(KEYINPUT56), .B(G16), .Z(n998) );
  XNOR2_X1 U1069 ( .A(G171), .B(G1961), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n974), .B(G1956), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(G1341), .B(n977), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G168), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1076 ( .A(KEYINPUT57), .B(n982), .Z(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n996) );
  XNOR2_X1 U1079 ( .A(G1348), .B(KEYINPUT124), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(n988), .B(n987), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(G1971), .A2(G303), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n1021) );
  XNOR2_X1 U1087 ( .A(G2090), .B(G35), .ZN(n1011) );
  XOR2_X1 U1088 ( .A(G1991), .B(G25), .Z(n999) );
  NAND2_X1 U1089 ( .A1(n999), .A2(G28), .ZN(n1008) );
  XNOR2_X1 U1090 ( .A(G1996), .B(G32), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(G33), .B(G2072), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(G2067), .B(G26), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G27), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(KEYINPUT53), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XOR2_X1 U1100 ( .A(G2084), .B(G34), .Z(n1012) );
  XNOR2_X1 U1101 ( .A(KEYINPUT54), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(n1016), .B(n1015), .ZN(n1018) );
  INV_X1 U1104 ( .A(G29), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(G11), .A2(n1019), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1110 ( .A(n1026), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

