//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971;
  XNOR2_X1  g000(.A(G64gat), .B(G92gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT78), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G8gat), .ZN(new_n204));
  INV_X1    g003(.A(G36gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT76), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT22), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G197gat), .B(G204gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND3_X1   g011(.A1(new_n211), .A2(KEYINPUT22), .A3(new_n207), .ZN(new_n213));
  OR3_X1    g012(.A1(new_n212), .A2(G218gat), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(G218gat), .B1(new_n212), .B2(new_n213), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT77), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n214), .A2(KEYINPUT77), .A3(new_n215), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  INV_X1    g023(.A(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n223), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT65), .ZN(new_n231));
  NOR2_X1   g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n232), .B1(KEYINPUT23), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n234), .B1(KEYINPUT23), .B2(new_n232), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n223), .A2(new_n228), .A3(new_n236), .A4(new_n229), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n231), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n234), .A2(new_n221), .ZN(new_n239));
  INV_X1    g038(.A(new_n222), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(new_n227), .A3(new_n226), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n232), .B(KEYINPUT66), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n239), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n232), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT66), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n247), .A2(KEYINPUT66), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT23), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n251), .A2(new_n239), .A3(KEYINPUT67), .A4(new_n241), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n221), .A2(new_n238), .B1(new_n246), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n224), .A2(new_n225), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n243), .A2(KEYINPUT26), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT26), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n233), .B1(new_n232), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n255), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT27), .B(G183gat), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT28), .B1(new_n260), .B2(new_n225), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT69), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n260), .B(KEYINPUT70), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(KEYINPUT28), .A3(new_n225), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n259), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G226gat), .ZN(new_n266));
  INV_X1    g065(.A(G233gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n253), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n265), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n238), .A2(new_n221), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n246), .A2(new_n252), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT68), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT68), .B1(new_n272), .B2(new_n273), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n268), .A2(KEYINPUT29), .ZN(new_n277));
  AOI211_X1 g076(.A(new_n220), .B(new_n270), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n271), .B(new_n268), .C1(new_n274), .C2(new_n275), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n277), .B1(new_n253), .B2(new_n265), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n216), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n206), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n281), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n276), .A2(new_n277), .ZN(new_n284));
  INV_X1    g083(.A(new_n220), .ZN(new_n285));
  INV_X1    g084(.A(new_n270), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n206), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n282), .A2(new_n289), .A3(KEYINPUT30), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n283), .A2(new_n287), .A3(new_n291), .A4(new_n288), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G227gat), .A2(G233gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G120gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G113gat), .ZN(new_n298));
  INV_X1    g097(.A(G113gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G120gat), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT1), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G127gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G134gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n301), .A2(new_n302), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n302), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(G134gat), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n272), .A2(new_n273), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT68), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n253), .A2(KEYINPUT68), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n310), .B1(new_n315), .B2(new_n271), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n310), .B(new_n271), .C1(new_n274), .C2(new_n275), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n296), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(KEYINPUT71), .A2(KEYINPUT33), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(KEYINPUT71), .A2(KEYINPUT33), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n319), .A2(KEYINPUT32), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT72), .B(G71gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(G99gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(G15gat), .B(G43gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n327), .B(new_n328), .Z(new_n329));
  AND3_X1   g128(.A1(new_n324), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n325), .B1(new_n324), .B2(new_n329), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT75), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n324), .A2(new_n329), .ZN(new_n333));
  INV_X1    g132(.A(new_n325), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n324), .A2(new_n325), .A3(new_n329), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT34), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n276), .A2(new_n309), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(new_n295), .A3(new_n317), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n341), .A2(new_n342), .A3(new_n339), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n341), .A4(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n346), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT74), .B1(new_n348), .B2(new_n343), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n338), .A3(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n330), .A2(new_n331), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n352), .A2(new_n336), .A3(new_n347), .A4(new_n349), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT36), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G78gat), .B(G106gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n357), .B(G22gat), .Z(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G148gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G141gat), .ZN(new_n361));
  INV_X1    g160(.A(G141gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G148gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT79), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT2), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n366), .B1(G155gat), .B2(G162gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n361), .A2(new_n363), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n365), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(G155gat), .B(G162gat), .Z(new_n372));
  XOR2_X1   g171(.A(KEYINPUT80), .B(G141gat), .Z(new_n373));
  OAI21_X1  g172(.A(new_n361), .B1(new_n373), .B2(new_n360), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n372), .A2(new_n367), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n371), .A2(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n285), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n377), .B1(new_n216), .B2(KEYINPUT29), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n371), .A2(new_n372), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n374), .A2(new_n375), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n381), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT87), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT31), .B(G50gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n380), .A2(new_n216), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n387), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n394), .B(KEYINPUT86), .Z(new_n395));
  AND3_X1   g194(.A1(new_n390), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n392), .B1(new_n390), .B2(new_n395), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n359), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n390), .A2(new_n395), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n391), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n390), .A2(new_n392), .A3(new_n395), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n358), .A3(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n351), .A2(new_n353), .A3(KEYINPUT36), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n356), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n354), .A2(new_n403), .A3(KEYINPUT35), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n294), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n305), .A2(new_n376), .A3(new_n409), .A4(new_n308), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n410), .A2(KEYINPUT83), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(KEYINPUT83), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n305), .A2(new_n376), .A3(new_n308), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT4), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  XOR2_X1   g214(.A(KEYINPUT81), .B(KEYINPUT5), .Z(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n385), .A2(KEYINPUT3), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(new_n309), .A3(new_n378), .ZN(new_n419));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n415), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n414), .A2(new_n410), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(new_n420), .A3(new_n419), .ZN(new_n424));
  INV_X1    g223(.A(new_n420), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n310), .A2(new_n376), .ZN(new_n426));
  INV_X1    g225(.A(new_n413), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n428), .A3(new_n416), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n417), .B1(new_n421), .B2(new_n423), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT82), .B1(new_n432), .B2(new_n428), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n422), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT0), .B(G57gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(G85gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(G1gat), .B(G29gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n422), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n429), .A2(new_n430), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n432), .A2(KEYINPUT82), .A3(new_n428), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT6), .B1(new_n444), .B2(new_n438), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n440), .B1(new_n446), .B2(KEYINPUT84), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(KEYINPUT84), .B2(new_n446), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n434), .A2(KEYINPUT6), .A3(new_n439), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT85), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n444), .A2(new_n438), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(KEYINPUT85), .A3(KEYINPUT6), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n408), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n420), .B1(new_n415), .B2(new_n419), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n426), .A2(new_n427), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n459), .B(KEYINPUT39), .C1(new_n425), .C2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT39), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n439), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT40), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n466), .A2(new_n452), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n465), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n290), .A2(KEYINPUT88), .A3(new_n292), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT88), .B1(new_n290), .B2(new_n292), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n467), .B(new_n468), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT37), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(new_n278), .B2(new_n281), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n283), .A2(KEYINPUT37), .A3(new_n287), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n206), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT89), .B1(new_n477), .B2(KEYINPUT38), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT89), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT38), .ZN(new_n480));
  AOI211_X1 g279(.A(new_n479), .B(new_n480), .C1(new_n476), .C2(new_n206), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n289), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n445), .A2(new_n440), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n279), .A2(new_n216), .A3(new_n280), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n270), .B1(new_n276), .B2(new_n277), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n484), .B(KEYINPUT37), .C1(new_n485), .C2(new_n285), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n474), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n487), .A2(new_n480), .A3(new_n206), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n453), .A2(new_n451), .A3(new_n483), .A4(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n472), .B1(new_n482), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n356), .A2(new_n490), .A3(new_n403), .A4(new_n405), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n451), .A2(new_n453), .A3(new_n483), .ZN(new_n492));
  INV_X1    g291(.A(new_n471), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n492), .A2(new_n469), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n354), .A2(new_n494), .A3(new_n403), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT35), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n457), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(G57gat), .B(G64gat), .Z(new_n501));
  OR2_X1    g300(.A1(G71gat), .A2(G78gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(G71gat), .A2(G78gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT9), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n501), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G57gat), .B(G64gat), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n503), .B(new_n502), .C1(new_n508), .C2(new_n505), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT21), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n512), .B(new_n513), .Z(new_n514));
  XNOR2_X1  g313(.A(G127gat), .B(G155gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(new_n207), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT93), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n519), .A2(G1gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT91), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT16), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n519), .B1(new_n523), .B2(G1gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n525), .A3(G8gat), .ZN(new_n526));
  INV_X1    g325(.A(G8gat), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n520), .B(new_n524), .C1(new_n521), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n510), .A2(new_n511), .ZN(new_n530));
  OR3_X1    g329(.A1(new_n529), .A2(G183gat), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(G183gat), .B1(new_n529), .B2(new_n530), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n518), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(new_n518), .A3(new_n532), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n534), .A2(G231gat), .A3(G233gat), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G231gat), .A2(G233gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n535), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n537), .B1(new_n538), .B2(new_n533), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n517), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n536), .A2(new_n539), .A3(new_n517), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n514), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n542), .ZN(new_n544));
  INV_X1    g343(.A(new_n514), .ZN(new_n545));
  NOR3_X1   g344(.A1(new_n544), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT41), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT97), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT14), .ZN(new_n552));
  INV_X1    g351(.A(G29gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n553), .A3(new_n205), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n554), .A2(new_n555), .B1(G29gat), .B2(G36gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(G43gat), .B(G50gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n556), .B1(KEYINPUT15), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(KEYINPUT15), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n561));
  NOR2_X1   g360(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n562));
  INV_X1    g361(.A(G85gat), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  OAI22_X1  g363(.A1(new_n561), .A2(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT95), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT7), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(G85gat), .A2(G92gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT8), .A2(new_n572), .B1(new_n563), .B2(new_n564), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n565), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n577), .A3(new_n572), .ZN(new_n578));
  AND2_X1   g377(.A1(G99gat), .A2(G106gat), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT96), .B1(new_n579), .B2(new_n575), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n574), .A2(new_n581), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n560), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n548), .A2(new_n549), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n551), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI221_X1 g386(.A(KEYINPUT97), .B1(new_n549), .B2(new_n548), .C1(new_n560), .C2(new_n584), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n558), .B(new_n559), .Z(new_n590));
  AOI21_X1  g389(.A(KEYINPUT17), .B1(new_n590), .B2(KEYINPUT90), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT90), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n560), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n584), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n550), .B1(new_n589), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n589), .A2(new_n595), .A3(new_n550), .ZN(new_n598));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT94), .B(KEYINPUT98), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n597), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n598), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n601), .B1(new_n604), .B2(new_n596), .ZN(new_n605));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n606), .B1(new_n603), .B2(new_n605), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n547), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G148gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT102), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n297), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n507), .A2(new_n509), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(new_n582), .B2(new_n583), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n565), .A2(new_n571), .A3(new_n573), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n578), .A2(new_n580), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n574), .A2(new_n581), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n510), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(KEYINPUT99), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n625), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n629), .A3(new_n620), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n619), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  AOI211_X1 g433(.A(KEYINPUT101), .B(new_n632), .C1(new_n627), .C2(new_n630), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n628), .A2(KEYINPUT10), .A3(new_n620), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n618), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n631), .A2(new_n617), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n616), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n631), .A2(new_n633), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT101), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n631), .A2(new_n619), .A3(new_n633), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n637), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n617), .ZN(new_n645));
  INV_X1    g444(.A(new_n639), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n646), .A3(new_n615), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n640), .A2(KEYINPUT103), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n649), .B(new_n616), .C1(new_n638), .C2(new_n639), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n529), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(new_n591), .B2(new_n594), .ZN(new_n654));
  NAND2_X1  g453(.A1(G229gat), .A2(G233gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n590), .A2(new_n529), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT18), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OR3_X1    g458(.A1(new_n590), .A2(new_n529), .A3(KEYINPUT92), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT92), .B1(new_n590), .B2(new_n529), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(new_n656), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n655), .B(KEYINPUT13), .Z(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n654), .A2(KEYINPUT18), .A3(new_n655), .A4(new_n656), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n659), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT11), .B(G169gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G197gat), .ZN(new_n668));
  XOR2_X1   g467(.A(G113gat), .B(G141gat), .Z(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT12), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n659), .A2(new_n671), .A3(new_n664), .A4(new_n665), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n652), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n500), .A2(new_n611), .A3(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n456), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT104), .B(G1gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1324gat));
  INV_X1    g480(.A(new_n678), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n470), .A2(new_n471), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT16), .B(G8gat), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n682), .A2(KEYINPUT42), .A3(new_n684), .A4(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n500), .A2(new_n611), .A3(new_n684), .A4(new_n677), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(G8gat), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n688), .B2(new_n685), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n687), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n687), .A2(KEYINPUT105), .A3(new_n691), .A4(new_n689), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(G1325gat));
  INV_X1    g495(.A(new_n354), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n678), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n356), .A2(new_n405), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n356), .A2(KEYINPUT106), .A3(new_n405), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G15gat), .ZN(new_n705));
  OAI22_X1  g504(.A1(new_n698), .A2(G15gat), .B1(new_n678), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT107), .ZN(G1326gat));
  NOR2_X1   g506(.A1(new_n678), .A2(new_n403), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT43), .B(G22gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  AND2_X1   g509(.A1(new_n677), .A2(new_n547), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n500), .A2(new_n610), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n553), .A3(new_n455), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n498), .B1(new_n408), .B2(new_n456), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n717), .B2(new_n609), .ZN(new_n718));
  AOI211_X1 g517(.A(new_n455), .B(new_n294), .C1(new_n406), .C2(new_n407), .ZN(new_n719));
  OAI211_X1 g518(.A(KEYINPUT44), .B(new_n610), .C1(new_n719), .C2(new_n498), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n547), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n722), .A2(new_n652), .A3(new_n676), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n721), .A2(new_n455), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G29gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n715), .A2(new_n725), .ZN(G1328gat));
  NAND4_X1  g525(.A1(new_n718), .A2(new_n684), .A3(new_n720), .A4(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G36gat), .ZN(new_n728));
  NAND2_X1  g527(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n712), .A2(new_n205), .A3(new_n684), .A4(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n717), .A2(new_n609), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n731), .A2(new_n205), .A3(new_n684), .A4(new_n711), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n728), .A2(new_n730), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT110), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n728), .A2(new_n730), .A3(new_n734), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1329gat));
  NOR2_X1   g538(.A1(new_n697), .A2(G43gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n712), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n718), .A2(new_n704), .A3(new_n720), .A4(new_n723), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n742), .A2(KEYINPUT111), .B1(G43gat), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n718), .A2(new_n699), .A3(new_n720), .A4(new_n723), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n745), .A2(KEYINPUT47), .A3(G43gat), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n741), .B1(new_n747), .B2(KEYINPUT47), .ZN(new_n748));
  OAI22_X1  g547(.A1(new_n744), .A2(KEYINPUT47), .B1(new_n746), .B2(new_n748), .ZN(G1330gat));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT48), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n500), .A2(new_n610), .A3(new_n404), .A4(new_n711), .ZN(new_n752));
  INV_X1    g551(.A(G50gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n718), .A2(new_n404), .A3(new_n720), .A4(new_n723), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n751), .B(new_n754), .C1(new_n755), .C2(new_n753), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n750), .A2(KEYINPUT48), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1331gat));
  NAND3_X1  g557(.A1(new_n611), .A2(new_n676), .A3(new_n652), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n717), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n455), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G57gat), .ZN(G1332gat));
  INV_X1    g561(.A(new_n760), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n683), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  AND2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n764), .B2(new_n765), .ZN(G1333gat));
  INV_X1    g567(.A(G71gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n763), .B2(new_n697), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n717), .A2(new_n769), .A3(new_n759), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n771), .A2(KEYINPUT113), .A3(new_n704), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT113), .B1(new_n771), .B2(new_n704), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT50), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n776), .B(new_n770), .C1(new_n772), .C2(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1334gat));
  NAND2_X1  g577(.A1(new_n760), .A2(new_n404), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n722), .A2(new_n675), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n652), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT114), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n721), .A2(G85gat), .A3(new_n783), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n610), .B(new_n781), .C1(new_n719), .C2(new_n498), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT51), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n500), .A2(new_n787), .A3(new_n610), .A4(new_n781), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n786), .A2(new_n788), .A3(new_n455), .A4(new_n652), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n784), .A2(new_n455), .B1(new_n563), .B2(new_n789), .ZN(G1336gat));
  NAND4_X1  g589(.A1(new_n718), .A2(new_n684), .A3(new_n720), .A4(new_n783), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G92gat), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n683), .A2(G92gat), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n786), .A2(new_n788), .A3(new_n652), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n792), .A2(KEYINPUT115), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT52), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n792), .A2(KEYINPUT115), .A3(new_n794), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(G1337gat));
  NAND3_X1  g598(.A1(new_n721), .A2(new_n704), .A3(new_n783), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G99gat), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n697), .A2(G99gat), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n788), .A3(new_n652), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(G1338gat));
  NAND4_X1  g603(.A1(new_n718), .A2(new_n404), .A3(new_n720), .A4(new_n783), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G106gat), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n786), .A2(new_n788), .A3(new_n404), .A4(new_n652), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(G106gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT53), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n806), .B(new_n810), .C1(new_n807), .C2(G106gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1339gat));
  NAND3_X1  g611(.A1(new_n611), .A2(new_n676), .A3(new_n651), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n642), .A2(new_n618), .A3(new_n637), .A4(new_n643), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT54), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n638), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n644), .A2(new_n818), .A3(new_n617), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n616), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n814), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n645), .A2(KEYINPUT54), .A3(new_n815), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n822), .A2(KEYINPUT55), .A3(new_n616), .A4(new_n819), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n662), .A2(new_n663), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n655), .B1(new_n654), .B2(new_n656), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n670), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n674), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n821), .A2(new_n823), .A3(new_n647), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n609), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n648), .A2(new_n650), .A3(new_n827), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT116), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n648), .A2(new_n827), .A3(new_n832), .A4(new_n650), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n821), .A2(new_n823), .A3(new_n675), .A4(new_n647), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n829), .B1(new_n835), .B2(new_n609), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n813), .B1(new_n836), .B2(new_n722), .ZN(new_n837));
  AND4_X1   g636(.A1(new_n455), .A2(new_n837), .A3(new_n403), .A4(new_n354), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n683), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n839), .A2(new_n676), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(new_n299), .ZN(G1340gat));
  NOR2_X1   g640(.A1(new_n839), .A2(new_n651), .ZN(new_n842));
  XNOR2_X1  g641(.A(KEYINPUT117), .B(G120gat), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n842), .B(new_n843), .ZN(G1341gat));
  NOR2_X1   g643(.A1(new_n839), .A2(new_n547), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(new_n302), .ZN(G1342gat));
  NAND2_X1  g645(.A1(new_n683), .A2(new_n610), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT118), .Z(new_n848));
  NAND3_X1  g647(.A1(new_n838), .A2(new_n304), .A3(new_n848), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n849), .A2(KEYINPUT56), .ZN(new_n850));
  OAI21_X1  g649(.A(G134gat), .B1(new_n839), .B2(new_n609), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(KEYINPUT56), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(G1343gat));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n404), .ZN(new_n854));
  NOR4_X1   g653(.A1(new_n704), .A2(new_n456), .A3(new_n684), .A4(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n362), .A3(new_n675), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n834), .A2(new_n833), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n610), .B1(new_n860), .B2(new_n831), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n547), .B1(new_n861), .B2(new_n829), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n403), .B1(new_n862), .B2(new_n813), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n859), .B1(new_n863), .B2(KEYINPUT57), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n834), .A2(new_n830), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n609), .ZN(new_n866));
  INV_X1    g665(.A(new_n829), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n722), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR4_X1   g667(.A1(new_n547), .A2(new_n610), .A3(new_n652), .A4(new_n675), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n404), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n854), .A2(KEYINPUT119), .A3(new_n871), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n864), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n356), .A2(new_n455), .A3(new_n683), .A4(new_n405), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n675), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT58), .B1(new_n878), .B2(new_n373), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n855), .A2(KEYINPUT121), .A3(new_n362), .A4(new_n675), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n858), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n856), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n875), .A2(KEYINPUT120), .A3(new_n877), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT120), .B1(new_n875), .B2(new_n877), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n675), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n882), .B1(new_n885), .B2(new_n373), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n881), .B1(new_n886), .B2(new_n887), .ZN(G1344gat));
  NAND2_X1  g687(.A1(new_n855), .A2(new_n652), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(KEYINPUT59), .A3(new_n360), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n870), .A2(KEYINPUT57), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n854), .A2(KEYINPUT57), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n895), .A2(KEYINPUT59), .A3(new_n652), .A4(new_n877), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT119), .B1(new_n854), .B2(new_n871), .ZN(new_n898));
  AOI211_X1 g697(.A(new_n859), .B(KEYINPUT57), .C1(new_n837), .C2(new_n404), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n898), .A2(new_n899), .A3(new_n872), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n897), .B1(new_n900), .B2(new_n876), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n875), .A2(KEYINPUT120), .A3(new_n877), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n651), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n896), .B1(new_n903), .B2(KEYINPUT59), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n891), .B1(new_n904), .B2(G148gat), .ZN(G1345gat));
  AOI21_X1  g704(.A(G155gat), .B1(new_n855), .B2(new_n722), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n901), .A2(new_n902), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n722), .A2(G155gat), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT122), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n906), .B1(new_n907), .B2(new_n909), .ZN(G1346gat));
  NOR3_X1   g709(.A1(new_n704), .A2(new_n456), .A3(new_n854), .ZN(new_n911));
  INV_X1    g710(.A(G162gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n912), .A3(new_n848), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n609), .B1(new_n901), .B2(new_n902), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n912), .ZN(G1347gat));
  AOI21_X1  g714(.A(new_n455), .B1(new_n862), .B2(new_n813), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n697), .A2(new_n404), .A3(new_n683), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(G169gat), .B1(new_n918), .B2(new_n676), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n917), .A2(KEYINPUT123), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n917), .A2(KEYINPUT123), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n916), .A3(new_n921), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(G169gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n923), .B2(new_n676), .ZN(G1348gat));
  INV_X1    g723(.A(G176gat), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n918), .A2(new_n925), .A3(new_n651), .ZN(new_n926));
  INV_X1    g725(.A(new_n922), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n652), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n928), .B2(new_n925), .ZN(G1349gat));
  NAND3_X1  g728(.A1(new_n927), .A2(new_n722), .A3(new_n263), .ZN(new_n930));
  OAI21_X1  g729(.A(G183gat), .B1(new_n918), .B2(new_n547), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g732(.A1(new_n927), .A2(new_n225), .A3(new_n610), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n916), .A2(new_n610), .A3(new_n917), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n935), .A2(new_n936), .A3(G190gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n935), .B2(G190gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(G1351gat));
  NAND3_X1  g738(.A1(new_n703), .A2(new_n456), .A3(new_n684), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n894), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n676), .ZN(new_n943));
  INV_X1    g742(.A(new_n940), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(KEYINPUT124), .A3(new_n863), .ZN(new_n945));
  INV_X1    g744(.A(G197gat), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n947), .B1(new_n940), .B2(new_n854), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n943), .B1(new_n676), .B2(new_n949), .ZN(G1352gat));
  NOR4_X1   g749(.A1(new_n940), .A2(G204gat), .A3(new_n651), .A4(new_n854), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT62), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n895), .A2(new_n944), .A3(new_n652), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G204gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1353gat));
  NAND2_X1  g754(.A1(new_n941), .A2(new_n722), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G211gat), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n957), .A2(new_n958), .A3(KEYINPUT63), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(KEYINPUT63), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n958), .A2(KEYINPUT63), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n956), .A2(G211gat), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n945), .A2(new_n207), .A3(new_n722), .A4(new_n948), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(KEYINPUT125), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(KEYINPUT125), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n959), .B(new_n962), .C1(new_n964), .C2(new_n965), .ZN(G1354gat));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n609), .B1(new_n942), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n208), .B1(new_n941), .B2(KEYINPUT127), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n945), .A2(new_n610), .A3(new_n948), .ZN(new_n970));
  INV_X1    g769(.A(G218gat), .ZN(new_n971));
  AOI22_X1  g770(.A1(new_n968), .A2(new_n969), .B1(new_n970), .B2(new_n971), .ZN(G1355gat));
endmodule


