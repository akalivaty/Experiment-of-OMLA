//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G235), .A3(G237), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT68), .Z(G261));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n452), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(G2106), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT69), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n465), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n461), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n472), .B1(G2104), .B2(new_n461), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NOR3_X1   g049(.A1(new_n474), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n475));
  OAI21_X1  g050(.A(G101), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n461), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n471), .A2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n466), .A2(new_n467), .ZN(new_n482));
  OR3_X1    g057(.A1(new_n482), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n478), .A2(KEYINPUT71), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  XOR2_X1   g063(.A(new_n488), .B(KEYINPUT72), .Z(new_n489));
  INV_X1    g064(.A(G112), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n474), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n482), .A2(new_n461), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n489), .A2(new_n491), .B1(new_n492), .B2(G124), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n487), .A2(new_n493), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n465), .A2(new_n468), .A3(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n495), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(KEYINPUT74), .C1(new_n467), .C2(new_n466), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT74), .B1(new_n477), .B2(new_n498), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G2105), .ZN(new_n505));
  OAI211_X1 g080(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n477), .A2(KEYINPUT73), .A3(G126), .A4(G2105), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n502), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G62), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(KEYINPUT75), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT75), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n514), .A2(new_n517), .A3(G62), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n513), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n514), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n520), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n519), .A2(new_n527), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n524), .B2(new_n531), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT5), .B(G543), .Z(new_n533));
  NAND2_X1  g108(.A1(new_n523), .A2(G89), .ZN(new_n534));
  NAND2_X1  g109(.A1(G63), .A2(G651), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n532), .A2(new_n536), .ZN(G168));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n538), .A2(new_n524), .B1(new_n525), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n513), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n513), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n521), .A2(new_n522), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n533), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n547), .A2(G81), .B1(new_n549), .B2(G43), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT76), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT76), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n545), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n533), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(new_n547), .B2(G91), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n524), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n549), .A2(new_n569), .A3(G53), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(KEYINPUT78), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(KEYINPUT78), .B1(new_n568), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n566), .B1(new_n572), .B2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  INV_X1    g150(.A(G168), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND2_X1  g152(.A1(new_n547), .A2(G87), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n549), .A2(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  INV_X1    g156(.A(G48), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n582), .A2(new_n524), .B1(new_n525), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n513), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n533), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n513), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n592), .B2(new_n591), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n547), .A2(G85), .B1(new_n549), .B2(G47), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n525), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n547), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n600), .A2(new_n601), .B1(G54), .B2(new_n549), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  INV_X1    g178(.A(G79), .ZN(new_n604));
  OAI22_X1  g179(.A1(new_n533), .A2(new_n603), .B1(new_n604), .B2(new_n548), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT80), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n607));
  OAI221_X1 g182(.A(new_n607), .B1(new_n604), .B2(new_n548), .C1(new_n533), .C2(new_n603), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n606), .A2(G651), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n597), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n597), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G299), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT81), .ZN(G148));
  INV_X1    g195(.A(KEYINPUT82), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n610), .B2(G559), .ZN(new_n622));
  NAND4_X1  g197(.A1(new_n602), .A2(KEYINPUT82), .A3(new_n618), .A4(new_n609), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n492), .A2(G123), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT83), .Z(new_n629));
  OR2_X1    g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n630), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(G135), .B2(new_n486), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2096), .ZN(new_n634));
  AND2_X1   g209(.A1(new_n465), .A2(new_n468), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n473), .A2(new_n475), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  INV_X1    g214(.A(G2100), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n634), .A2(new_n641), .A3(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT85), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(KEYINPUT14), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G1341), .B(G1348), .Z(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G14), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n654), .A2(new_n657), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XNOR2_X1  g237(.A(G2084), .B(G2090), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT86), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT88), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n665), .B(KEYINPUT17), .Z(new_n671));
  INV_X1    g246(.A(new_n666), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n669), .B(new_n670), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n663), .A2(new_n666), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n663), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n665), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n673), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2096), .B(G2100), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G227));
  XOR2_X1   g258(.A(G1971), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(new_n688), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT20), .Z(new_n692));
  AOI211_X1 g267(.A(new_n690), .B(new_n692), .C1(new_n685), .C2(new_n689), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT90), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n693), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT89), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n697), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  NOR2_X1   g278(.A1(G6), .A2(G16), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n587), .B2(G16), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT32), .ZN(new_n706));
  INV_X1    g281(.A(G1981), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G16), .A2(G23), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT91), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(G288), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT33), .ZN(new_n713));
  INV_X1    g288(.A(G1976), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(G16), .A2(G22), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G166), .B2(G16), .ZN(new_n717));
  INV_X1    g292(.A(G1971), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n708), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(KEYINPUT34), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT34), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n708), .A2(new_n722), .A3(new_n715), .A4(new_n719), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G25), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n486), .A2(G131), .ZN(new_n726));
  OAI21_X1  g301(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n727));
  INV_X1    g302(.A(G107), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(G2105), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n492), .B2(G119), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n725), .B1(new_n732), .B2(new_n724), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT35), .B(G1991), .Z(new_n734));
  XOR2_X1   g309(.A(new_n733), .B(new_n734), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n711), .A2(G24), .ZN(new_n736));
  INV_X1    g311(.A(G290), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(new_n711), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(G1986), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n738), .A2(G1986), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n735), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n721), .A2(new_n723), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT36), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n724), .A2(G32), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n636), .A2(G105), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT26), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n492), .A2(G129), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n486), .B2(G141), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n744), .B1(new_n750), .B2(new_n724), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT27), .B(G1996), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n751), .B(new_n752), .Z(new_n753));
  NAND2_X1  g328(.A1(G162), .A2(G29), .ZN(new_n754));
  OR2_X1    g329(.A1(G29), .A2(G35), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT29), .B(G2090), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n753), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G168), .A2(new_n711), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n711), .B2(G21), .ZN(new_n761));
  INV_X1    g336(.A(G1966), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n633), .A2(G29), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT31), .B(G11), .Z(new_n765));
  INV_X1    g340(.A(G28), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n766), .A2(KEYINPUT30), .ZN(new_n767));
  AOI21_X1  g342(.A(G29), .B1(new_n766), .B2(KEYINPUT30), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n761), .A2(new_n762), .ZN(new_n770));
  AND4_X1   g345(.A1(new_n763), .A2(new_n764), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n711), .A2(G5), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G171), .B2(new_n711), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1961), .ZN(new_n774));
  INV_X1    g349(.A(new_n756), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n757), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n759), .A2(new_n771), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n711), .A2(G19), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n556), .B2(new_n711), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1341), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n724), .A2(G27), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT95), .Z(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n511), .B2(G29), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G2078), .Z(new_n784));
  NOR3_X1   g359(.A1(new_n777), .A2(new_n780), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT25), .Z(new_n787));
  INV_X1    g362(.A(G139), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n485), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n635), .A2(G127), .ZN(new_n790));
  NAND2_X1  g365(.A1(G115), .A2(G2104), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n461), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(KEYINPUT92), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n795), .A2(G29), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G29), .B2(G33), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(G2072), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n711), .A2(G20), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT23), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n615), .B2(new_n711), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT96), .B(G1956), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(KEYINPUT24), .A2(G34), .ZN(new_n807));
  NOR2_X1   g382(.A1(KEYINPUT24), .A2(G34), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n724), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT93), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G160), .B2(G29), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(G2084), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT94), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n711), .A2(G4), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n611), .B2(new_n711), .ZN(new_n815));
  INV_X1    g390(.A(G1348), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n724), .A2(G26), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT28), .Z(new_n819));
  NAND3_X1  g394(.A1(new_n483), .A2(G140), .A3(new_n484), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n821));
  INV_X1    g396(.A(G116), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(G2105), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n492), .B2(G128), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n819), .B1(new_n825), .B2(G29), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G2067), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n811), .A2(G2084), .ZN(new_n828));
  AND4_X1   g403(.A1(new_n813), .A2(new_n817), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n785), .A2(new_n806), .A3(new_n829), .ZN(new_n830));
  AND3_X1   g405(.A1(new_n743), .A2(KEYINPUT97), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(KEYINPUT97), .B1(new_n743), .B2(new_n830), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(G311));
  NAND2_X1  g408(.A1(new_n743), .A2(new_n830), .ZN(G150));
  INV_X1    g409(.A(G55), .ZN(new_n835));
  INV_X1    g410(.A(G93), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n835), .A2(new_n524), .B1(new_n525), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(new_n513), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n555), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n551), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT38), .Z(new_n846));
  NOR2_X1   g421(.A1(new_n610), .A2(new_n618), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n849));
  AOI21_X1  g424(.A(G860), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n849), .B2(new_n848), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n841), .A2(G860), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT37), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(G145));
  NAND2_X1  g429(.A1(new_n492), .A2(G130), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n461), .A2(G118), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  INV_X1    g432(.A(G142), .ZN(new_n858));
  OAI221_X1 g433(.A(new_n855), .B1(new_n856), .B2(new_n857), .C1(new_n485), .C2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n638), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n795), .A2(KEYINPUT99), .A3(new_n797), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n820), .A2(KEYINPUT98), .A3(new_n824), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT98), .B1(new_n820), .B2(new_n824), .ZN(new_n865));
  OAI21_X1  g440(.A(G164), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n865), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(new_n511), .A3(new_n863), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n866), .A2(new_n868), .A3(new_n750), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n750), .B1(new_n866), .B2(new_n868), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n862), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n866), .A2(new_n868), .ZN(new_n872));
  INV_X1    g447(.A(new_n750), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n866), .A2(new_n868), .A3(new_n750), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n794), .B1(KEYINPUT92), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n871), .A2(new_n878), .A3(new_n731), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n731), .B1(new_n871), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n861), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n871), .A2(new_n878), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n732), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n871), .A2(new_n878), .A3(new_n731), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n860), .A3(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(G162), .B(G160), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n633), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n881), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n887), .B1(new_n881), .B2(new_n885), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT100), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n881), .A2(new_n885), .ZN(new_n893));
  INV_X1    g468(.A(new_n887), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n895), .A2(new_n896), .A3(new_n889), .A4(new_n888), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n892), .A2(KEYINPUT40), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT40), .B1(new_n892), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(G395));
  NAND2_X1  g475(.A1(new_n845), .A2(new_n624), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n842), .A2(new_n844), .A3(new_n622), .A4(new_n623), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n573), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n571), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n611), .A2(new_n905), .A3(new_n566), .ZN(new_n906));
  NAND2_X1  g481(.A1(G299), .A2(new_n610), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n903), .A2(KEYINPUT101), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT41), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n912), .A2(new_n901), .A3(new_n902), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT101), .B1(new_n903), .B2(new_n909), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT42), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G288), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n737), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(G290), .A2(G288), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT102), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n923), .A3(new_n920), .ZN(new_n924));
  XNOR2_X1  g499(.A(G166), .B(new_n587), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n925), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n927), .A2(new_n921), .A3(KEYINPUT102), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n903), .A2(new_n909), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n932), .A2(new_n933), .A3(new_n914), .A4(new_n910), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n917), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n929), .B1(new_n917), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g511(.A(G868), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n840), .A2(G868), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n937), .B2(new_n939), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(G295));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n939), .ZN(G331));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n926), .A2(new_n928), .ZN(new_n945));
  NAND2_X1  g520(.A1(G286), .A2(G171), .ZN(new_n946));
  NAND2_X1  g521(.A1(G301), .A2(G168), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n842), .A2(new_n844), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n946), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n840), .B1(new_n552), .B2(new_n554), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n949), .B1(new_n950), .B2(new_n843), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n912), .A2(new_n913), .A3(new_n948), .A4(new_n951), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n842), .A2(new_n844), .B1(new_n946), .B2(new_n947), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n949), .A2(new_n950), .A3(new_n843), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n909), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT104), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT41), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT41), .B1(new_n906), .B2(new_n907), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n953), .A2(new_n954), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n945), .B1(new_n956), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n952), .A2(KEYINPUT104), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n908), .B1(new_n948), .B2(new_n951), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n965), .B1(new_n960), .B2(new_n961), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n929), .B(new_n964), .C1(new_n966), .C2(KEYINPUT104), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n963), .A2(new_n967), .A3(new_n889), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n929), .A2(new_n966), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(G37), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n967), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n944), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI211_X1 g551(.A(KEYINPUT105), .B(KEYINPUT44), .C1(new_n969), .C2(new_n973), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n972), .B1(new_n971), .B2(new_n967), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n963), .A2(new_n967), .A3(new_n972), .A4(new_n889), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT44), .ZN(new_n980));
  OAI22_X1  g555(.A1(new_n976), .A2(new_n977), .B1(new_n978), .B2(new_n980), .ZN(G397));
  XNOR2_X1  g556(.A(new_n731), .B(new_n734), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT107), .Z(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n511), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  INV_X1    g561(.A(G40), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n471), .A2(new_n987), .A3(new_n480), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n983), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n750), .B(G1996), .ZN(new_n992));
  INV_X1    g567(.A(G2067), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n825), .B(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n989), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT106), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n991), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(G290), .B(G1986), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n990), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT122), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n985), .A2(new_n986), .ZN(new_n1001));
  AOI21_X1  g576(.A(G1384), .B1(new_n502), .B2(new_n510), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT45), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n988), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1000), .B1(new_n1004), .B2(G2078), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT53), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1000), .B(new_n1007), .C1(new_n1004), .C2(G2078), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n988), .B1(new_n1002), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n511), .A2(new_n1009), .A3(new_n984), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1002), .A2(KEYINPUT108), .A3(new_n1009), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1015), .A2(G1961), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1006), .A2(new_n1008), .A3(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G301), .A2(KEYINPUT123), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(G171), .ZN(new_n1019));
  OAI221_X1 g594(.A(KEYINPUT54), .B1(new_n1017), .B2(new_n1018), .C1(new_n1019), .C2(KEYINPUT123), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1019), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1017), .A2(G171), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n482), .A2(G2105), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n636), .A2(G101), .B1(new_n1027), .B2(G137), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n469), .A2(new_n470), .ZN(new_n1029));
  OAI211_X1 g604(.A(G40), .B(new_n1028), .C1(new_n1029), .C2(new_n461), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1002), .A2(KEYINPUT45), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n988), .B1(new_n1002), .B2(KEYINPUT45), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n1032), .A2(G2084), .B1(G1966), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT111), .B(G8), .Z(new_n1038));
  NOR2_X1   g613(.A1(G168), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1025), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1038), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1036), .A2(G286), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1036), .A2(new_n1042), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1039), .A2(KEYINPUT51), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1041), .A2(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1038), .B1(new_n988), .B2(new_n1002), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n714), .B2(G288), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n918), .A2(G1976), .ZN(new_n1049));
  OR3_X1    g624(.A1(new_n1048), .A2(KEYINPUT52), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(KEYINPUT52), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G305), .A2(G1981), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n587), .A2(new_n707), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT49), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1052), .A2(KEYINPUT49), .A3(new_n1053), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1047), .A3(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1050), .A2(new_n1051), .A3(new_n1058), .ZN(new_n1059));
  OAI22_X1  g634(.A1(new_n1032), .A2(G2090), .B1(G1971), .B2(new_n1035), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1061));
  NAND3_X1  g636(.A1(G303), .A2(G8), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1061), .ZN(new_n1063));
  INV_X1    g638(.A(G8), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(G166), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1066), .A2(KEYINPUT110), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(KEYINPUT110), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1060), .A2(new_n1067), .A3(G8), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1066), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1011), .A2(KEYINPUT112), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT112), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1002), .A2(new_n1072), .A3(new_n1009), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1010), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G2090), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1074), .A2(new_n1075), .B1(new_n1004), .B2(new_n718), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1070), .B1(new_n1076), .B2(new_n1038), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1059), .A2(new_n1069), .A3(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1020), .A2(new_n1024), .A3(new_n1046), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n988), .A2(new_n1002), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(G2067), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(KEYINPUT60), .B(new_n1082), .C1(new_n1015), .C2(G1348), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n611), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT120), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1081), .B1(new_n1032), .B2(new_n816), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1086), .A2(new_n1087), .A3(KEYINPUT60), .A4(new_n610), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT119), .B1(new_n1083), .B2(new_n611), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1083), .A2(new_n1090), .A3(new_n611), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1085), .A2(new_n1088), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1086), .A2(KEYINPUT60), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT121), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT56), .B(G2072), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1001), .A2(new_n988), .A3(new_n1003), .A4(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1074), .B2(G1956), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n568), .A2(new_n570), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1099), .A2(new_n1100), .A3(new_n566), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1002), .A2(new_n1072), .A3(new_n1009), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1072), .B1(new_n1002), .B2(new_n1009), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1031), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G1956), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1107), .A2(new_n1108), .B1(new_n1035), .B2(new_n1096), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT113), .B1(new_n1109), .B2(new_n1102), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1102), .B(new_n1097), .C1(new_n1074), .C2(G1956), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT113), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1104), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(KEYINPUT118), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1119), .A2(KEYINPUT113), .A3(new_n1097), .A4(new_n1102), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1118), .A2(new_n1120), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1117), .B1(new_n1121), .B2(KEYINPUT61), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT115), .B(KEYINPUT58), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(G1341), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1080), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1004), .B2(G1996), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n555), .B1(KEYINPUT116), .B2(KEYINPUT59), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT117), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT117), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1127), .A2(new_n1131), .A3(new_n1128), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(KEYINPUT116), .A2(KEYINPUT59), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1130), .B(new_n1132), .C1(KEYINPUT116), .C2(KEYINPUT59), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT114), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1102), .B1(new_n1098), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1137), .B2(new_n1098), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1115), .B1(new_n1109), .B2(new_n1102), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1135), .A2(new_n1136), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1092), .A2(new_n1142), .A3(new_n1093), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1095), .A2(new_n1123), .A3(new_n1141), .A4(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1139), .B1(new_n610), .B2(new_n1086), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1079), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1058), .A2(new_n714), .A3(new_n918), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1053), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1047), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1059), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(new_n1069), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1044), .A2(G286), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1153), .A2(new_n1077), .A3(new_n1069), .A4(new_n1059), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT63), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1044), .A2(new_n1155), .A3(G286), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1060), .A2(G8), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1070), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1157), .A2(new_n1069), .A3(new_n1059), .A4(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1152), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1046), .A2(KEYINPUT62), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1078), .A2(new_n1022), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1046), .A2(KEYINPUT62), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1161), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n999), .B1(new_n1147), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n989), .A2(G1996), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT46), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n989), .B1(new_n994), .B2(new_n750), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(KEYINPUT124), .B(KEYINPUT47), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1171), .B(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n825), .A2(G2067), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n732), .A2(new_n734), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1174), .B1(new_n996), .B2(new_n1175), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n989), .A2(G1986), .A3(G290), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT48), .ZN(new_n1178));
  OAI221_X1 g753(.A(new_n1173), .B1(new_n1176), .B2(new_n989), .C1(new_n997), .C2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT125), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1179), .B(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1167), .A2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g757(.A1(new_n661), .A2(new_n682), .A3(G319), .ZN(new_n1184));
  INV_X1    g758(.A(KEYINPUT126), .ZN(new_n1185));
  XNOR2_X1  g759(.A(new_n1184), .B(new_n1185), .ZN(new_n1186));
  NAND2_X1  g760(.A1(new_n1186), .A2(new_n702), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n1187), .A2(KEYINPUT127), .ZN(new_n1188));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n1189));
  NAND3_X1  g763(.A1(new_n1186), .A2(new_n702), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n892), .A2(new_n897), .ZN(new_n1192));
  AND3_X1   g766(.A1(new_n1191), .A2(new_n1192), .A3(new_n974), .ZN(G308));
  NAND3_X1  g767(.A1(new_n1191), .A2(new_n1192), .A3(new_n974), .ZN(G225));
endmodule


