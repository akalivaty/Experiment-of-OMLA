//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n209));
  INV_X1    g0009(.A(G244), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n209), .B1(new_n202), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n208), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT65), .Z(new_n218));
  INV_X1    g0018(.A(KEYINPUT1), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n218), .A2(new_n219), .ZN(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n206), .ZN(new_n225));
  AND2_X1   g0025(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n208), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NOR4_X1   g0029(.A1(new_n220), .A2(new_n221), .A3(new_n226), .A4(new_n229), .ZN(G361));
  XOR2_X1   g0030(.A(G226), .B(G232), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT67), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  INV_X1    g0042(.A(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT68), .B(G50), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(new_n224), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(G222), .A3(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n256), .B(KEYINPUT70), .Z(new_n257));
  AND3_X1   g0057(.A1(new_n254), .A2(G223), .A3(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n258), .B1(G77), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n253), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G274), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n252), .A2(KEYINPUT69), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT69), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G33), .A3(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(new_n272), .A3(new_n251), .ZN(new_n273));
  INV_X1    g0073(.A(new_n268), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G226), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n269), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n265), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT72), .ZN(new_n280));
  INV_X1    g0080(.A(G190), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(KEYINPUT72), .B1(new_n278), .B2(G190), .ZN(new_n283));
  INV_X1    g0083(.A(G200), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT71), .ZN(new_n287));
  AOI21_X1  g0087(.A(KEYINPUT10), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G150), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n206), .A2(G33), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n290), .B1(new_n201), .B2(new_n206), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n224), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n295), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n205), .A2(G20), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(G50), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G13), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G1), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G20), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n296), .B(new_n299), .C1(G50), .C2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT9), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n286), .A2(new_n304), .ZN(new_n305));
  XOR2_X1   g0105(.A(new_n288), .B(new_n305), .Z(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n279), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n278), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n303), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(G58), .B(G68), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n313), .A2(G20), .B1(G159), .B2(new_n289), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT77), .B1(new_n259), .B2(KEYINPUT3), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT77), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(new_n261), .A3(G33), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n317), .A3(new_n260), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT7), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(new_n319), .A3(new_n206), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G68), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n319), .B1(new_n318), .B2(new_n206), .ZN(new_n322));
  OAI211_X1 g0122(.A(KEYINPUT16), .B(new_n314), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT7), .B1(new_n254), .B2(G20), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n263), .A2(new_n319), .A3(new_n206), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(new_n325), .A3(G68), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n314), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT16), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n323), .A2(new_n329), .A3(new_n295), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n291), .B1(new_n205), .B2(G20), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n300), .A2(new_n206), .A3(G1), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(new_n295), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n331), .A2(new_n333), .B1(new_n332), .B2(new_n291), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT78), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT18), .ZN(new_n337));
  NOR2_X1   g0137(.A1(G223), .A2(G1698), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(new_n276), .B2(G1698), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n339), .A2(new_n260), .A3(new_n315), .A4(new_n317), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G87), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n253), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G232), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n269), .B1(new_n275), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G179), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n307), .B2(new_n345), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n336), .A2(new_n337), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n337), .B1(new_n336), .B2(new_n347), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT79), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n276), .A2(G1698), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(G223), .B2(G1698), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n341), .B1(new_n318), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n253), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n224), .B1(KEYINPUT69), .B2(new_n252), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n268), .B1(new_n357), .B2(new_n272), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G232), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n356), .A2(new_n281), .A3(new_n269), .A4(new_n359), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n360), .B(KEYINPUT80), .C1(new_n345), .C2(G200), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT80), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n345), .A2(new_n362), .A3(new_n281), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n361), .A2(new_n330), .A3(new_n335), .A4(new_n363), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT17), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n336), .A2(new_n347), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT18), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT79), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n368), .A3(new_n348), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n351), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n292), .A2(new_n202), .B1(new_n206), .B2(G68), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT73), .B1(new_n289), .B2(G50), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n289), .A2(KEYINPUT73), .A3(G50), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n297), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT11), .ZN(new_n376));
  INV_X1    g0176(.A(G68), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n332), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT12), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n375), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT11), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n297), .A2(new_n302), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n298), .A2(G68), .ZN(new_n384));
  OR3_X1    g0184(.A1(new_n383), .A2(KEYINPUT74), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT74), .B1(new_n383), .B2(new_n384), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n381), .A2(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n358), .A2(G238), .ZN(new_n388));
  INV_X1    g0188(.A(G97), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n259), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(G226), .A2(G1698), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n343), .B2(G1698), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n392), .B2(new_n254), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n388), .B(new_n269), .C1(new_n253), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT13), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n393), .A2(new_n253), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT13), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n396), .A2(new_n397), .A3(new_n269), .A4(new_n388), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n380), .B(new_n387), .C1(new_n399), .C2(new_n281), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n284), .B1(new_n395), .B2(new_n398), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT75), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n399), .B2(new_n309), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n395), .A2(new_n398), .A3(KEYINPUT75), .A4(G179), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n399), .A2(G169), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT14), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT14), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n399), .A2(new_n409), .A3(G169), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n385), .A2(new_n386), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(KEYINPUT11), .B2(new_n375), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n376), .A2(new_n379), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT76), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT76), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n387), .A2(new_n416), .A3(new_n376), .A4(new_n379), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n402), .B1(new_n411), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(G232), .A2(G1698), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n255), .A2(G238), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n254), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n422), .B(new_n355), .C1(G107), .C2(new_n254), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n423), .B(new_n269), .C1(new_n210), .C2(new_n275), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G200), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n297), .A2(G77), .A3(new_n298), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(G77), .B2(new_n302), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G20), .A2(G77), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n206), .A2(new_n259), .ZN(new_n430));
  OAI221_X1 g0230(.A(new_n428), .B1(new_n429), .B2(new_n292), .C1(new_n430), .C2(new_n291), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n427), .B1(new_n431), .B2(new_n295), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n425), .B(new_n432), .C1(new_n281), .C2(new_n424), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n432), .B1(new_n307), .B2(new_n424), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n424), .A2(G179), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n419), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n312), .A2(new_n370), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G33), .A2(G294), .ZN(new_n440));
  INV_X1    g0240(.A(G250), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n255), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(G257), .B2(new_n255), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n440), .B1(new_n318), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n355), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n267), .A2(G1), .ZN(new_n446));
  AND2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n273), .A2(new_n449), .A3(G264), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT5), .B(G41), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n273), .A2(G274), .A3(new_n446), .A4(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n445), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n307), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(G179), .B2(new_n453), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n332), .A2(KEYINPUT25), .A3(new_n211), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT25), .B1(new_n332), .B2(new_n211), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n205), .A2(G33), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n297), .A2(new_n302), .A3(new_n458), .ZN(new_n459));
  OAI22_X1  g0259(.A1(new_n456), .A2(new_n457), .B1(new_n459), .B2(new_n211), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n315), .A2(new_n317), .A3(new_n260), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n461), .A2(KEYINPUT22), .A3(new_n206), .A4(G87), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT24), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT22), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n206), .A2(G87), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n464), .B1(new_n263), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G116), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G20), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT23), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n206), .B2(G107), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n211), .A2(KEYINPUT23), .A3(G20), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n462), .A2(new_n463), .A3(new_n466), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n466), .A2(new_n472), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT22), .A2(G87), .ZN(new_n475));
  NOR3_X1   g0275(.A1(new_n318), .A2(G20), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT24), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n460), .B1(new_n478), .B2(new_n295), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n455), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n445), .A2(new_n281), .A3(new_n450), .A4(new_n452), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT90), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n272), .A2(new_n357), .B1(new_n451), .B2(new_n446), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n444), .A2(new_n355), .B1(new_n483), .B2(G264), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT90), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n484), .A2(new_n485), .A3(new_n281), .A4(new_n452), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n453), .A2(new_n284), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n482), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n479), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT91), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n488), .A2(new_n479), .A3(KEYINPUT91), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n480), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n273), .B(G250), .C1(G1), .C2(new_n267), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n446), .A2(G274), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT85), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n210), .A2(G1698), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(G238), .B2(G1698), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n461), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n497), .B1(new_n501), .B2(new_n467), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n497), .B(new_n467), .C1(new_n318), .C2(new_n499), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n355), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n496), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G200), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n496), .B(G190), .C1(new_n502), .C2(new_n504), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n461), .A2(new_n206), .A3(G68), .ZN(new_n508));
  XOR2_X1   g0308(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n509));
  NOR2_X1   g0309(.A1(new_n292), .A2(new_n389), .ZN(new_n510));
  OR2_X1    g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(G20), .B1(new_n509), .B2(new_n390), .ZN(new_n512));
  NOR3_X1   g0312(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n508), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(new_n295), .B1(new_n332), .B2(new_n429), .ZN(new_n515));
  INV_X1    g0315(.A(G87), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n459), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT88), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n517), .B(new_n518), .ZN(new_n519));
  AND4_X1   g0319(.A1(new_n506), .A2(new_n507), .A3(new_n515), .A4(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n496), .B(new_n309), .C1(new_n502), .C2(new_n504), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n494), .A2(new_n495), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n503), .A2(new_n355), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n467), .B1(new_n318), .B2(new_n499), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT85), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n522), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n521), .B1(new_n526), .B2(G169), .ZN(new_n527));
  INV_X1    g0327(.A(new_n459), .ZN(new_n528));
  INV_X1    g0328(.A(new_n429), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n527), .A2(KEYINPUT86), .B1(new_n515), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT86), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n532), .B(new_n521), .C1(new_n526), .C2(G169), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n520), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n261), .A2(G33), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n536));
  OAI21_X1  g0336(.A(G303), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n212), .A2(G1698), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(G257), .B2(G1698), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n537), .B1(new_n318), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n355), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n273), .A2(new_n449), .A3(G270), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n452), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n333), .A2(G116), .A3(new_n458), .ZN(new_n544));
  INV_X1    g0344(.A(G116), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n332), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n294), .A2(new_n224), .B1(G20), .B2(new_n545), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G283), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n548), .B(new_n206), .C1(G33), .C2(new_n389), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n547), .A2(KEYINPUT20), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT20), .B1(new_n547), .B2(new_n549), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n544), .B(new_n546), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n543), .A2(KEYINPUT21), .A3(G169), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n452), .A2(new_n542), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n552), .A2(new_n555), .A3(G179), .A4(new_n541), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(KEYINPUT89), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT89), .B1(new_n553), .B2(new_n556), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n307), .B1(new_n555), .B2(new_n541), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT21), .B1(new_n560), .B2(new_n552), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n555), .A2(G190), .A3(new_n541), .ZN(new_n562));
  NOR2_X1   g0362(.A1(G257), .A2(G1698), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n212), .B2(G1698), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n564), .A2(new_n260), .A3(new_n315), .A4(new_n317), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n253), .B1(new_n565), .B2(new_n537), .ZN(new_n566));
  OAI21_X1  g0366(.A(G200), .B1(new_n566), .B2(new_n554), .ZN(new_n567));
  INV_X1    g0367(.A(new_n552), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n562), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NOR4_X1   g0369(.A1(new_n558), .A2(new_n559), .A3(new_n561), .A4(new_n569), .ZN(new_n570));
  XOR2_X1   g0370(.A(G97), .B(G107), .Z(new_n571));
  XNOR2_X1  g0371(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n389), .A2(G107), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(G20), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n324), .A2(new_n325), .A3(G107), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n289), .A2(G77), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n295), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT82), .B1(new_n302), .B2(G97), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT82), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n332), .A2(new_n582), .A3(new_n389), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n389), .B2(new_n459), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n483), .A2(G257), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n452), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n255), .A2(G244), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n590), .A2(new_n591), .B1(new_n441), .B2(new_n255), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(new_n254), .B1(G33), .B2(G283), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n210), .A2(G1698), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n315), .A2(new_n317), .A3(new_n260), .A4(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT83), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n593), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n589), .B1(new_n600), .B2(new_n355), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n587), .B1(G190), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT84), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n317), .A2(new_n260), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n604), .A2(KEYINPUT83), .A3(new_n315), .A4(new_n594), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(new_n597), .A3(new_n591), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n253), .B1(new_n606), .B2(new_n593), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n603), .B1(new_n607), .B2(new_n589), .ZN(new_n608));
  INV_X1    g0408(.A(new_n589), .ZN(new_n609));
  INV_X1    g0409(.A(new_n593), .ZN(new_n610));
  INV_X1    g0410(.A(new_n599), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n610), .B1(new_n611), .B2(new_n597), .ZN(new_n612));
  OAI211_X1 g0412(.A(KEYINPUT84), .B(new_n609), .C1(new_n612), .C2(new_n253), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n608), .A2(new_n613), .A3(G200), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n585), .B1(new_n579), .B2(new_n295), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n609), .B1(new_n612), .B2(new_n253), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n616), .B2(new_n307), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n601), .A2(new_n309), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n602), .A2(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n493), .A2(new_n534), .A3(new_n570), .A4(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n439), .A2(new_n620), .ZN(G372));
  INV_X1    g0421(.A(new_n311), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n349), .A2(new_n350), .ZN(new_n623));
  INV_X1    g0423(.A(new_n402), .ZN(new_n624));
  INV_X1    g0424(.A(new_n436), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n418), .A2(new_n411), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n365), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n622), .B1(new_n306), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n515), .A2(new_n519), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n523), .A2(KEYINPUT92), .A3(new_n525), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT92), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n502), .B2(new_n504), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n522), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n630), .B(new_n507), .C1(new_n284), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n515), .A2(new_n530), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n521), .B(new_n636), .C1(new_n634), .C2(G169), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n491), .A2(new_n492), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n639), .A3(new_n619), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n553), .A2(new_n556), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n480), .A2(new_n641), .A3(new_n561), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n618), .B(new_n587), .C1(G169), .C2(new_n601), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n534), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT26), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n638), .A2(new_n649), .A3(new_n646), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n650), .A2(new_n637), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n644), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n629), .B1(new_n439), .B2(new_n653), .ZN(G369));
  NAND2_X1  g0454(.A1(new_n301), .A2(new_n206), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(G213), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n639), .B1(new_n479), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n480), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n559), .ZN(new_n665));
  INV_X1    g0465(.A(new_n561), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n557), .A3(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n667), .A2(new_n661), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n480), .A2(new_n661), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n664), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n669), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n664), .A2(new_n669), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n661), .A2(new_n568), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n641), .B2(new_n561), .ZN(new_n675));
  INV_X1    g0475(.A(new_n569), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n665), .A2(new_n557), .A3(new_n666), .A4(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n675), .B1(new_n677), .B2(new_n674), .ZN(new_n678));
  XOR2_X1   g0478(.A(KEYINPUT93), .B(G330), .Z(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n673), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n672), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n227), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n513), .A2(new_n545), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n686), .A2(new_n687), .A3(new_n205), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n223), .B2(new_n686), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT28), .Z(new_n690));
  INV_X1    g0490(.A(KEYINPUT96), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n660), .A2(KEYINPUT31), .ZN(new_n692));
  INV_X1    g0492(.A(new_n634), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n453), .A2(new_n543), .A3(new_n309), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n601), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n541), .A2(G179), .A3(new_n452), .A4(new_n542), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n445), .A2(new_n450), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n601), .A3(new_n526), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n703), .A2(KEYINPUT94), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n505), .A2(new_n698), .A3(new_n697), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT95), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n705), .A2(new_n706), .A3(KEYINPUT30), .A4(new_n601), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n699), .A2(new_n601), .A3(KEYINPUT30), .A4(new_n526), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT95), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n703), .A2(KEYINPUT94), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n692), .B1(new_n704), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT31), .B1(new_n620), .B2(new_n660), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n709), .A2(new_n707), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n693), .A2(new_n695), .B1(new_n700), .B2(new_n701), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n661), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n711), .B1(new_n712), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n691), .B1(new_n717), .B2(new_n679), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n608), .A2(new_n613), .A3(G200), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n615), .B1(new_n616), .B2(new_n281), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n645), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n677), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(new_n493), .A3(new_n534), .A4(new_n661), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n715), .B1(new_n723), .B2(KEYINPUT31), .ZN(new_n724));
  OAI211_X1 g0524(.A(KEYINPUT96), .B(new_n680), .C1(new_n724), .C2(new_n711), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n718), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n652), .A2(new_n661), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT29), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n667), .A2(new_n480), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n640), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n635), .A2(new_n637), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT26), .B1(new_n733), .B2(new_n645), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n534), .A2(new_n649), .A3(new_n646), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n734), .A2(new_n735), .A3(new_n637), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n660), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT29), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n730), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n727), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n690), .B1(new_n741), .B2(G1), .ZN(G364));
  INV_X1    g0542(.A(new_n681), .ZN(new_n743));
  INV_X1    g0543(.A(new_n686), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n300), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n205), .B1(new_n745), .B2(G45), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n744), .A2(KEYINPUT97), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT97), .ZN(new_n748));
  INV_X1    g0548(.A(new_n746), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n748), .B1(new_n686), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n743), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(new_n680), .B2(new_n678), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G13), .A2(G33), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n755), .B(KEYINPUT98), .Z(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n224), .B1(G20), .B2(new_n307), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n223), .A2(new_n267), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n685), .A2(new_n461), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n760), .B(new_n762), .C1(new_n246), .C2(G45), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n685), .A2(new_n263), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G355), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G116), .B2(new_n227), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n759), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n206), .A2(G190), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n284), .A2(G179), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n211), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n206), .A2(new_n281), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n769), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n263), .B(new_n771), .C1(G87), .C2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT99), .Z(new_n776));
  NOR2_X1   g0576(.A1(G179), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n768), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G159), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT32), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n206), .B1(new_n777), .B2(G190), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n389), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n309), .A2(new_n284), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n772), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G50), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n309), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n772), .A2(new_n787), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n785), .A2(new_n786), .B1(new_n788), .B2(new_n243), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n784), .A2(new_n768), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n787), .A2(new_n768), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n790), .A2(new_n377), .B1(new_n791), .B2(new_n202), .ZN(new_n792));
  NOR4_X1   g0592(.A1(new_n781), .A2(new_n783), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n790), .ZN(new_n794));
  INV_X1    g0594(.A(G317), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(KEYINPUT33), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n795), .A2(KEYINPUT33), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n794), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G322), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n799), .B2(new_n788), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT100), .Z(new_n801));
  INV_X1    g0601(.A(new_n785), .ZN(new_n802));
  INV_X1    g0602(.A(new_n791), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n802), .A2(G326), .B1(new_n803), .B2(G311), .ZN(new_n804));
  INV_X1    g0604(.A(new_n770), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G303), .A2(new_n774), .B1(new_n805), .B2(G283), .ZN(new_n806));
  INV_X1    g0606(.A(new_n782), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G294), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n254), .B1(new_n779), .B2(G329), .ZN(new_n809));
  AND4_X1   g0609(.A1(new_n804), .A2(new_n806), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n776), .A2(new_n793), .B1(new_n801), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n758), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n767), .B(new_n752), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT101), .ZN(new_n814));
  INV_X1    g0614(.A(new_n757), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n678), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n754), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  OAI21_X1  g0618(.A(new_n433), .B1(new_n432), .B2(new_n661), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n436), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n625), .A2(new_n661), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n728), .B(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n824), .A2(new_n726), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n751), .B1(new_n824), .B2(new_n726), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n790), .A2(new_n828), .B1(new_n791), .B2(new_n545), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT102), .Z(new_n830));
  AOI22_X1  g0630(.A1(G303), .A2(new_n802), .B1(new_n774), .B2(G107), .ZN(new_n831));
  INV_X1    g0631(.A(new_n788), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G294), .A2(new_n832), .B1(new_n779), .B2(G311), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n254), .B(new_n783), .C1(G87), .C2(new_n805), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n830), .A2(new_n831), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n778), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n770), .A2(new_n377), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n837), .B(new_n838), .C1(G50), .C2(new_n774), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n318), .B1(G58), .B2(new_n807), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G143), .A2(new_n832), .B1(new_n803), .B2(G159), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  INV_X1    g0642(.A(G150), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n841), .B1(new_n842), .B2(new_n785), .C1(new_n843), .C2(new_n790), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT34), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n839), .B(new_n840), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n835), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n758), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n758), .A2(new_n755), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n751), .B1(new_n202), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n849), .B(new_n851), .C1(new_n823), .C2(new_n756), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n827), .A2(new_n852), .ZN(G384));
  NOR2_X1   g0653(.A1(new_n745), .A2(new_n205), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n438), .A2(new_n730), .A3(new_n738), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n629), .ZN(new_n856));
  INV_X1    g0656(.A(new_n658), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n623), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n418), .B(new_n660), .C1(new_n411), .C2(new_n402), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n415), .A2(new_n417), .A3(new_n660), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n861), .B(new_n402), .C1(new_n411), .C2(new_n418), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n648), .A2(new_n637), .A3(new_n650), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n661), .B(new_n823), .C1(new_n864), .C2(new_n643), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n863), .B1(new_n865), .B2(new_n821), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n314), .B1(new_n321), .B2(new_n322), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n328), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(new_n295), .A3(new_n323), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n658), .B1(new_n869), .B2(new_n334), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n370), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n347), .A2(new_n857), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n334), .B2(new_n869), .ZN(new_n873));
  INV_X1    g0673(.A(new_n364), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n336), .A2(new_n857), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n366), .A2(new_n876), .A3(new_n364), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(KEYINPUT37), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n871), .A2(new_n878), .A3(KEYINPUT38), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n858), .B1(new_n866), .B2(new_n883), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n877), .B(KEYINPUT37), .Z(new_n885));
  AOI21_X1  g0685(.A(new_n876), .B1(new_n365), .B2(new_n623), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n880), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n882), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT39), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n411), .A2(new_n418), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n891), .A2(new_n660), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n890), .B(new_n892), .C1(new_n883), .C2(new_n889), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n884), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n856), .B(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT103), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n713), .A2(new_n714), .ZN(new_n897));
  AND4_X1   g0697(.A1(new_n896), .A2(new_n897), .A3(KEYINPUT31), .A4(new_n660), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n715), .B2(KEYINPUT31), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n712), .A2(new_n716), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n438), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n823), .B1(new_n860), .B2(new_n862), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n900), .B2(new_n901), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(KEYINPUT40), .A3(new_n888), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n871), .A2(new_n878), .A3(KEYINPUT38), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT38), .B1(new_n871), .B2(new_n878), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n861), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n419), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n822), .B1(new_n913), .B2(new_n859), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n898), .A2(new_n899), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(new_n724), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n908), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT104), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(KEYINPUT104), .B(new_n908), .C1(new_n911), .C2(new_n916), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n907), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n903), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n903), .A2(new_n921), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n680), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n854), .B1(new_n895), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n895), .B2(new_n924), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n573), .A2(new_n575), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n927), .A2(KEYINPUT35), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(KEYINPUT35), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n928), .A2(G116), .A3(new_n225), .A4(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT36), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n223), .B(G77), .C1(new_n243), .C2(new_n377), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(G50), .B2(new_n377), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(G1), .A3(new_n300), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n926), .A2(new_n931), .A3(new_n934), .ZN(G367));
  INV_X1    g0735(.A(new_n670), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n619), .B1(new_n615), .B2(new_n661), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n646), .A2(new_n660), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n480), .B1(new_n719), .B2(new_n720), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n660), .B1(new_n942), .B2(new_n645), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n940), .B2(KEYINPUT42), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n630), .A2(new_n661), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n638), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n945), .A2(new_n637), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n941), .A2(new_n944), .B1(KEYINPUT43), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n949), .B(new_n950), .Z(new_n951));
  INV_X1    g0751(.A(new_n939), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n683), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n686), .B(KEYINPUT41), .Z(new_n955));
  AOI21_X1  g0755(.A(new_n668), .B1(new_n664), .B2(new_n669), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n936), .A2(new_n743), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n743), .B1(new_n936), .B2(new_n956), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n741), .A2(KEYINPUT106), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n727), .A2(new_n739), .A3(new_n959), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT106), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n671), .A2(new_n952), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT44), .ZN(new_n965));
  XOR2_X1   g0765(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n966));
  NAND3_X1  g0766(.A1(new_n672), .A2(new_n939), .A3(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n966), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n671), .B2(new_n952), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n682), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT44), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n964), .B(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n973), .A2(new_n683), .A3(new_n967), .A4(new_n969), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n960), .A2(new_n963), .A3(new_n971), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n955), .B1(new_n975), .B2(new_n741), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n954), .B1(new_n976), .B2(new_n749), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n759), .B1(new_n227), .B2(new_n429), .C1(new_n762), .C2(new_n240), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT107), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n751), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n979), .B2(new_n978), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n773), .A2(new_n243), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n254), .B1(new_n788), .B2(new_n843), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(G143), .C2(new_n802), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n770), .A2(new_n202), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G137), .B2(new_n779), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G159), .A2(new_n794), .B1(new_n803), .B2(G50), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n807), .A2(G68), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n984), .A2(new_n986), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n773), .B2(new_n545), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT110), .ZN(new_n992));
  XNOR2_X1  g0792(.A(KEYINPUT108), .B(G311), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n785), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n770), .A2(new_n389), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n994), .A2(new_n995), .A3(new_n461), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G303), .A2(new_n832), .B1(new_n779), .B2(G317), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n773), .A2(new_n545), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n998), .A2(KEYINPUT46), .B1(G107), .B2(new_n807), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G294), .A2(new_n794), .B1(new_n803), .B2(G283), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n996), .A2(new_n997), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n989), .B1(new_n992), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT47), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n981), .B1(new_n1003), .B2(new_n758), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n948), .B2(new_n815), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n977), .A2(new_n1005), .ZN(G387));
  NAND2_X1  g0806(.A1(new_n960), .A2(new_n963), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1007), .B(new_n686), .C1(new_n741), .C2(new_n959), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n764), .A2(new_n687), .B1(new_n211), .B2(new_n685), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n236), .A2(new_n267), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n291), .A2(G50), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT50), .ZN(new_n1012));
  AOI211_X1 g0812(.A(G45), .B(new_n687), .C1(G68), .C2(G77), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n762), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT111), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1009), .B1(new_n1010), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n759), .ZN(new_n1017));
  INV_X1    g0817(.A(G159), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n785), .A2(new_n1018), .B1(new_n790), .B2(new_n291), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G50), .B2(new_n832), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n995), .B1(G68), .B2(new_n803), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G77), .A2(new_n774), .B1(new_n779), .B2(G150), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n782), .A2(new_n429), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1023), .A2(new_n318), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G116), .A2(new_n805), .B1(new_n779), .B2(G326), .ZN(new_n1026));
  INV_X1    g0826(.A(G294), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n773), .A2(new_n1027), .B1(new_n782), .B2(new_n828), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n785), .A2(new_n799), .B1(new_n788), .B2(new_n795), .ZN(new_n1029));
  INV_X1    g0829(.A(G303), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n790), .A2(new_n993), .B1(new_n791), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1028), .B1(new_n1032), .B2(KEYINPUT48), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(KEYINPUT48), .B2(new_n1032), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT49), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n318), .B(new_n1026), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1025), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n758), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1017), .A2(new_n752), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n673), .B2(new_n757), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n959), .B2(new_n749), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1008), .A2(new_n1042), .ZN(G393));
  AND2_X1   g0843(.A1(new_n975), .A2(new_n686), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n971), .A2(new_n974), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1007), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n759), .B1(new_n389), .B2(new_n227), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n249), .B2(new_n761), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n790), .A2(new_n786), .B1(new_n791), .B2(new_n291), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n782), .A2(new_n202), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT112), .Z(new_n1053));
  OAI22_X1  g0853(.A1(new_n785), .A2(new_n843), .B1(new_n788), .B2(new_n1018), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT51), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n773), .A2(new_n377), .B1(new_n770), .B2(new_n516), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n318), .B(new_n1056), .C1(G143), .C2(new_n779), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1053), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G317), .A2(new_n802), .B1(new_n832), .B2(G311), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT52), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n254), .B(new_n771), .C1(G116), .C2(new_n807), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G303), .A2(new_n794), .B1(new_n803), .B2(G294), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G283), .A2(new_n774), .B1(new_n779), .B2(G322), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1058), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n751), .B(new_n1049), .C1(new_n1065), .C2(new_n758), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n939), .B2(new_n815), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1045), .B2(new_n746), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT113), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1047), .A2(new_n1072), .ZN(G390));
  NAND2_X1  g0873(.A1(new_n737), .A2(new_n820), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n821), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n863), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n892), .B1(new_n887), .B2(new_n882), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n890), .B1(new_n883), .B2(new_n889), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n892), .B2(new_n866), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n726), .A2(new_n914), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n905), .A2(G330), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n749), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n751), .B1(new_n291), .B2(new_n850), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n774), .A2(G150), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT53), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G159), .B2(new_n807), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n794), .A2(G137), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n802), .A2(G128), .B1(new_n779), .B2(G125), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT54), .B(G143), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1094), .A2(new_n791), .B1(new_n770), .B2(new_n786), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n263), .B(new_n1095), .C1(G132), .C2(new_n832), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1096), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n254), .B(new_n1051), .C1(G87), .C2(new_n774), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n838), .B1(G116), .B2(new_n832), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n802), .A2(G283), .B1(new_n779), .B2(G294), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n790), .A2(new_n211), .B1(new_n791), .B2(new_n389), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT118), .Z(new_n1103));
  OAI21_X1  g0903(.A(new_n1097), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1104), .A2(KEYINPUT119), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(KEYINPUT119), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n758), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1080), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1088), .B1(new_n1105), .B2(new_n1107), .C1(new_n1108), .C2(new_n756), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1087), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT117), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n822), .B1(new_n718), .B2(new_n725), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1084), .B1(new_n1112), .B2(new_n1076), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n865), .A2(new_n821), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(G330), .B(new_n823), .C1(new_n724), .C2(new_n915), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT114), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1116), .A2(new_n1117), .A3(new_n863), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1117), .B1(new_n1116), .B2(new_n863), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1075), .B1(new_n726), .B2(new_n914), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT115), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1122), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1115), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n438), .A2(G330), .A3(new_n902), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n855), .A2(new_n1126), .A3(new_n629), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT116), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n1084), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n686), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(KEYINPUT116), .B(new_n1086), .C1(new_n1125), .C2(new_n1128), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1111), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT115), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1127), .B1(new_n1139), .B2(new_n1115), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1086), .B1(new_n1140), .B2(KEYINPUT116), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT116), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n1132), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1141), .A2(KEYINPUT117), .A3(new_n686), .A4(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1110), .B1(new_n1135), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(G378));
  XOR2_X1   g0947(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n303), .A2(new_n857), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT55), .Z(new_n1151));
  NAND2_X1  g0951(.A1(new_n312), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n312), .A2(new_n1151), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1149), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1154), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1156), .A2(new_n1148), .A3(new_n1152), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1158), .A2(new_n756), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n790), .A2(new_n836), .B1(new_n791), .B2(new_n842), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT120), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n807), .A2(G150), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n832), .A2(G128), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1094), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G125), .A2(new_n802), .B1(new_n774), .B2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1165), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1168));
  AOI211_X1 g0968(.A(G33), .B(G41), .C1(new_n779), .C2(G124), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n1018), .B2(new_n770), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1167), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G77), .A2(new_n774), .B1(new_n803), .B2(new_n529), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G107), .A2(new_n832), .B1(new_n805), .B2(G58), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n1173), .A3(new_n988), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G97), .A2(new_n794), .B1(new_n779), .B2(G283), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n545), .B2(new_n785), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n318), .A2(new_n266), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1174), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1178), .A2(KEYINPUT58), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(KEYINPUT58), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1177), .B(new_n786), .C1(G33), .C2(G41), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n758), .B1(new_n1171), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n751), .B1(new_n786), .B2(new_n850), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1159), .A2(new_n1185), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n921), .A2(G330), .A3(new_n894), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n894), .B1(new_n921), .B2(G330), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1158), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n921), .A2(G330), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n894), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n921), .A2(G330), .A3(new_n894), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1189), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1186), .B1(new_n1196), .B2(new_n749), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1137), .A2(new_n1138), .B1(new_n1114), .B2(new_n1113), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1128), .B1(new_n1198), .B2(new_n1132), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1196), .A2(new_n1199), .A3(KEYINPUT57), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n686), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1197), .B1(new_n1201), .B2(new_n1202), .ZN(G375));
  OAI21_X1  g1003(.A(KEYINPUT122), .B1(new_n1198), .B2(new_n746), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT122), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1125), .A2(new_n1205), .A3(new_n749), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n863), .A2(new_n755), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n751), .B1(new_n377), .B2(new_n850), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n773), .A2(new_n389), .B1(new_n778), .B2(new_n1030), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT123), .Z(new_n1210));
  AOI22_X1  g1010(.A1(G116), .A2(new_n794), .B1(new_n832), .B2(G283), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n802), .A2(G294), .B1(new_n803), .B2(G107), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n985), .A2(new_n1023), .A3(new_n254), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT124), .Z(new_n1215));
  OAI22_X1  g1015(.A1(new_n842), .A2(new_n788), .B1(new_n773), .B2(new_n1018), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G150), .B2(new_n803), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n794), .A2(new_n1164), .B1(new_n805), .B2(G58), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n802), .A2(G132), .B1(new_n779), .B2(G128), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n318), .B1(G50), .B2(new_n807), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1215), .A2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1222), .A2(KEYINPUT125), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(KEYINPUT125), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n758), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1207), .B(new_n1208), .C1(new_n1223), .C2(new_n1225), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1204), .A2(new_n1206), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1198), .A2(new_n1127), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n955), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(new_n1142), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(G381));
  INV_X1    g1031(.A(G375), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1141), .A2(new_n686), .A3(new_n1144), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1110), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(G393), .A2(G396), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1044), .A2(new_n1046), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1238));
  INV_X1    g1038(.A(G384), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  OR4_X1    g1040(.A1(G387), .A2(new_n1236), .A3(G381), .A4(new_n1240), .ZN(G407));
  OAI211_X1 g1041(.A(G407), .B(G213), .C1(G343), .C2(new_n1236), .ZN(G409));
  INV_X1    g1042(.A(new_n1197), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1196), .A2(new_n1199), .A3(new_n1229), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1234), .B(new_n1233), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1146), .B2(G375), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n659), .A2(G213), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT126), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1239), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1198), .A2(KEYINPUT60), .A3(new_n1127), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT60), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n744), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1251), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1204), .A2(new_n1206), .A3(new_n1226), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1248), .B(new_n1250), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1251), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1227), .A2(new_n1249), .A3(new_n1239), .A4(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1246), .A2(new_n1247), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT62), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n659), .A2(G213), .A3(G2897), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1257), .A2(new_n1259), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT61), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1246), .A2(new_n1270), .A3(new_n1247), .A4(new_n1260), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1262), .A2(new_n1268), .A3(new_n1269), .A4(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT127), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G387), .A2(new_n1238), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(G390), .A2(new_n977), .A3(new_n1005), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n817), .B1(new_n1008), .B2(new_n1042), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1237), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1272), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT61), .B1(new_n1263), .B2(new_n1267), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1261), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1246), .A2(KEYINPUT63), .A3(new_n1247), .A4(new_n1260), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1286), .A2(new_n1283), .A3(new_n1288), .A4(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1285), .A2(new_n1290), .ZN(G405));
  INV_X1    g1091(.A(new_n1260), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1146), .A2(G375), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(G375), .B2(new_n1235), .ZN(new_n1295));
  OR2_X1    g1095(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1296), .A2(new_n1260), .A3(new_n1280), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1293), .A2(new_n1295), .A3(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1295), .B1(new_n1293), .B2(new_n1297), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(G402));
endmodule


