

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803;

  XNOR2_X1 U379 ( .A(G143), .B(G104), .ZN(n450) );
  XNOR2_X1 U380 ( .A(n407), .B(n476), .ZN(n365) );
  XNOR2_X1 U381 ( .A(n473), .B(G128), .ZN(n474) );
  BUF_X4 U382 ( .A(G953), .Z(n798) );
  NAND2_X4 U383 ( .A1(n663), .A2(n798), .ZN(n690) );
  XNOR2_X1 U384 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n505) );
  XNOR2_X1 U385 ( .A(G143), .B(G128), .ZN(n405) );
  XNOR2_X1 U386 ( .A(KEYINPUT16), .B(G122), .ZN(n499) );
  XOR2_X1 U387 ( .A(KEYINPUT105), .B(G122), .Z(n528) );
  INV_X2 U388 ( .A(G953), .ZN(n793) );
  AND2_X1 U389 ( .A1(n565), .A2(n631), .ZN(n357) );
  AND2_X2 U390 ( .A1(n430), .A2(KEYINPUT35), .ZN(n406) );
  XNOR2_X2 U391 ( .A(n435), .B(n561), .ZN(n622) );
  NOR2_X1 U392 ( .A1(n572), .A2(n402), .ZN(n573) );
  INV_X1 U393 ( .A(G119), .ZN(n473) );
  NOR2_X2 U394 ( .A1(G953), .A2(G237), .ZN(n517) );
  XNOR2_X2 U395 ( .A(G137), .B(G140), .ZN(n478) );
  NOR2_X1 U396 ( .A1(n398), .A2(n362), .ZN(n394) );
  XNOR2_X1 U397 ( .A(n641), .B(n363), .ZN(n398) );
  NOR2_X1 U398 ( .A1(n550), .A2(n599), .ZN(n608) );
  XNOR2_X1 U399 ( .A(n424), .B(KEYINPUT32), .ZN(n359) );
  NAND2_X1 U400 ( .A1(n357), .A2(n425), .ZN(n424) );
  INV_X2 U401 ( .A(n737), .ZN(n624) );
  XNOR2_X1 U402 ( .A(n360), .B(n553), .ZN(n589) );
  NAND2_X1 U403 ( .A1(n403), .A2(n751), .ZN(n360) );
  XNOR2_X1 U404 ( .A(n535), .B(n534), .ZN(n592) );
  XOR2_X1 U405 ( .A(KEYINPUT62), .B(n358), .Z(n675) );
  XOR2_X1 U406 ( .A(n367), .B(KEYINPUT59), .Z(n661) );
  XNOR2_X1 U407 ( .A(n532), .B(n531), .ZN(n680) );
  XNOR2_X1 U408 ( .A(n526), .B(n525), .ZN(n532) );
  XNOR2_X1 U409 ( .A(n434), .B(n433), .ZN(n501) );
  XNOR2_X1 U410 ( .A(n462), .B(KEYINPUT3), .ZN(n434) );
  INV_X1 U411 ( .A(G131), .ZN(n452) );
  XNOR2_X2 U412 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n448) );
  XNOR2_X2 U413 ( .A(G122), .B(G113), .ZN(n447) );
  XNOR2_X2 U414 ( .A(G146), .B(G125), .ZN(n503) );
  XNOR2_X2 U415 ( .A(KEYINPUT18), .B(KEYINPUT94), .ZN(n502) );
  XOR2_X1 U416 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n529) );
  XNOR2_X2 U417 ( .A(KEYINPUT69), .B(G101), .ZN(n508) );
  XOR2_X2 U418 ( .A(KEYINPUT4), .B(G131), .Z(n372) );
  BUF_X1 U419 ( .A(n674), .Z(n358) );
  NAND2_X1 U420 ( .A1(n359), .A2(n640), .ZN(n647) );
  XNOR2_X1 U421 ( .A(n359), .B(G119), .ZN(G21) );
  NAND2_X1 U422 ( .A1(n589), .A2(n559), .ZN(n435) );
  XNOR2_X2 U423 ( .A(n404), .B(n514), .ZN(n403) );
  XNOR2_X2 U424 ( .A(n361), .B(n563), .ZN(n425) );
  NAND2_X1 U425 ( .A1(n622), .A2(n371), .ZN(n361) );
  INV_X1 U426 ( .A(KEYINPUT89), .ZN(n362) );
  INV_X1 U427 ( .A(KEYINPUT66), .ZN(n363) );
  INV_X1 U428 ( .A(n454), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n407), .B(n476), .ZN(n791) );
  XNOR2_X1 U430 ( .A(n453), .B(n369), .ZN(n575) );
  AND2_X1 U431 ( .A1(n738), .A2(n425), .ZN(n633) );
  XNOR2_X1 U432 ( .A(n639), .B(n638), .ZN(n400) );
  NOR2_X1 U433 ( .A1(n399), .A2(n396), .ZN(n395) );
  NOR2_X1 U434 ( .A1(n400), .A2(KEYINPUT89), .ZN(n399) );
  NOR2_X1 U435 ( .A1(n674), .A2(G902), .ZN(n453) );
  NAND2_X1 U436 ( .A1(n738), .A2(n425), .ZN(n366) );
  BUF_X1 U437 ( .A(n660), .Z(n367) );
  XNOR2_X1 U438 ( .A(n368), .B(G469), .ZN(n546) );
  NOR2_X1 U439 ( .A1(n693), .A2(G902), .ZN(n368) );
  NOR2_X2 U440 ( .A1(n760), .A2(n374), .ZN(n441) );
  XNOR2_X2 U441 ( .A(n461), .B(n423), .ZN(n789) );
  XNOR2_X1 U442 ( .A(G902), .B(KEYINPUT15), .ZN(n610) );
  NAND2_X1 U443 ( .A1(n413), .A2(n373), .ZN(n655) );
  OR2_X1 U444 ( .A1(n444), .A2(KEYINPUT87), .ZN(n417) );
  XNOR2_X1 U445 ( .A(n477), .B(n370), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n472), .B(n471), .ZN(n524) );
  INV_X1 U447 ( .A(KEYINPUT8), .ZN(n471) );
  XNOR2_X1 U448 ( .A(n451), .B(n450), .ZN(n449) );
  XNOR2_X1 U449 ( .A(n452), .B(G140), .ZN(n451) );
  XNOR2_X1 U450 ( .A(n448), .B(n447), .ZN(n446) );
  INV_X1 U451 ( .A(KEYINPUT10), .ZN(n476) );
  BUF_X1 U452 ( .A(n564), .Z(n738) );
  XNOR2_X1 U453 ( .A(n738), .B(KEYINPUT93), .ZN(n603) );
  INV_X1 U454 ( .A(KEYINPUT48), .ZN(n445) );
  NOR2_X1 U455 ( .A1(n605), .A2(n717), .ZN(n606) );
  NAND2_X1 U456 ( .A1(n397), .A2(n650), .ZN(n396) );
  NAND2_X1 U457 ( .A1(n398), .A2(n362), .ZN(n397) );
  INV_X1 U458 ( .A(KEYINPUT107), .ZN(n456) );
  AND2_X1 U459 ( .A1(n440), .A2(n618), .ZN(n436) );
  NOR2_X1 U460 ( .A1(G237), .A2(G902), .ZN(n466) );
  XNOR2_X1 U461 ( .A(n546), .B(KEYINPUT1), .ZN(n564) );
  XNOR2_X1 U462 ( .A(G137), .B(KEYINPUT5), .ZN(n458) );
  XNOR2_X1 U463 ( .A(G119), .B(G116), .ZN(n433) );
  NOR2_X1 U464 ( .A1(n611), .A2(n610), .ZN(n411) );
  XNOR2_X1 U465 ( .A(n501), .B(n432), .ZN(n781) );
  XNOR2_X1 U466 ( .A(n500), .B(n499), .ZN(n432) );
  NAND2_X1 U467 ( .A1(G237), .A2(G234), .ZN(n493) );
  AND2_X1 U468 ( .A1(n741), .A2(n542), .ZN(n390) );
  XNOR2_X1 U469 ( .A(n475), .B(n386), .ZN(n385) );
  XNOR2_X1 U470 ( .A(G107), .B(G116), .ZN(n527) );
  XNOR2_X1 U471 ( .A(n520), .B(n519), .ZN(n660) );
  XNOR2_X1 U472 ( .A(n791), .B(n518), .ZN(n520) );
  XNOR2_X1 U473 ( .A(n449), .B(n446), .ZN(n519) );
  XNOR2_X1 U474 ( .A(n426), .B(KEYINPUT109), .ZN(n565) );
  NAND2_X1 U475 ( .A1(n603), .A2(n741), .ZN(n426) );
  XNOR2_X1 U476 ( .A(n376), .B(n375), .ZN(n595) );
  INV_X1 U477 ( .A(KEYINPUT79), .ZN(n375) );
  NOR2_X1 U478 ( .A1(n380), .A2(n574), .ZN(n378) );
  NOR2_X1 U479 ( .A1(n547), .A2(n408), .ZN(n548) );
  XOR2_X1 U480 ( .A(n465), .B(G472), .Z(n369) );
  INV_X1 U481 ( .A(n707), .ZN(n389) );
  XOR2_X1 U482 ( .A(G110), .B(KEYINPUT24), .Z(n370) );
  NOR2_X1 U483 ( .A1(n754), .A2(n740), .ZN(n371) );
  INV_X1 U484 ( .A(G902), .ZN(n533) );
  AND2_X1 U485 ( .A1(n417), .A2(n609), .ZN(n373) );
  XNOR2_X1 U486 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n374) );
  INV_X1 U487 ( .A(KEYINPUT35), .ZN(n429) );
  NAND2_X1 U488 ( .A1(n378), .A2(n377), .ZN(n376) );
  XNOR2_X1 U489 ( .A(n379), .B(KEYINPUT30), .ZN(n377) );
  INV_X1 U490 ( .A(n574), .ZN(n626) );
  NOR2_X2 U491 ( .A1(n575), .A2(n552), .ZN(n379) );
  NAND2_X1 U492 ( .A1(n624), .A2(n540), .ZN(n380) );
  XNOR2_X2 U493 ( .A(n382), .B(n381), .ZN(n500) );
  XNOR2_X2 U494 ( .A(G104), .B(KEYINPUT77), .ZN(n381) );
  XNOR2_X2 U495 ( .A(G110), .B(G107), .ZN(n382) );
  INV_X1 U496 ( .A(n479), .ZN(n687) );
  XNOR2_X1 U497 ( .A(n385), .B(n383), .ZN(n479) );
  XNOR2_X1 U498 ( .A(n384), .B(n365), .ZN(n383) );
  XNOR2_X1 U499 ( .A(n474), .B(n478), .ZN(n384) );
  NAND2_X1 U500 ( .A1(n455), .A2(n387), .ZN(n597) );
  NAND2_X1 U501 ( .A1(n388), .A2(KEYINPUT47), .ZN(n387) );
  NAND2_X1 U502 ( .A1(n389), .A2(n454), .ZN(n388) );
  NAND2_X1 U503 ( .A1(n390), .A2(n567), .ZN(n577) );
  NAND2_X1 U504 ( .A1(n391), .A2(n390), .ZN(n543) );
  INV_X1 U505 ( .A(n584), .ZN(n391) );
  XNOR2_X2 U506 ( .A(n392), .B(G143), .ZN(n523) );
  XNOR2_X2 U507 ( .A(G128), .B(G134), .ZN(n392) );
  NAND2_X1 U508 ( .A1(n395), .A2(n393), .ZN(n443) );
  NAND2_X1 U509 ( .A1(n400), .A2(n394), .ZN(n393) );
  INV_X1 U510 ( .A(n754), .ZN(n401) );
  NAND2_X1 U511 ( .A1(n751), .A2(n401), .ZN(n402) );
  INV_X2 U512 ( .A(n403), .ZN(n551) );
  NOR2_X2 U513 ( .A1(n668), .A2(n651), .ZN(n404) );
  XOR2_X2 U514 ( .A(KEYINPUT38), .B(n551), .Z(n572) );
  BUF_X1 U515 ( .A(n546), .Z(n574) );
  XNOR2_X1 U516 ( .A(n580), .B(n579), .ZN(n803) );
  XNOR2_X1 U517 ( .A(n470), .B(n469), .ZN(n410) );
  BUF_X1 U518 ( .A(n523), .Z(n526) );
  XNOR2_X1 U519 ( .A(n464), .B(n463), .ZN(n674) );
  XNOR2_X2 U520 ( .A(G146), .B(G125), .ZN(n407) );
  NOR2_X2 U521 ( .A1(n685), .A2(n803), .ZN(n583) );
  INV_X1 U522 ( .A(n738), .ZN(n408) );
  BUF_X1 U523 ( .A(n685), .Z(n409) );
  BUF_X1 U524 ( .A(n656), .Z(n776) );
  XNOR2_X1 U525 ( .A(n789), .B(n410), .ZN(n693) );
  INV_X1 U526 ( .A(n564), .ZN(n612) );
  NAND2_X1 U527 ( .A1(n642), .A2(KEYINPUT44), .ZN(n422) );
  NAND2_X1 U528 ( .A1(n420), .A2(n421), .ZN(n642) );
  NAND2_X1 U529 ( .A1(n411), .A2(n656), .ZN(n428) );
  XNOR2_X2 U530 ( .A(n443), .B(KEYINPUT45), .ZN(n656) );
  OR2_X2 U531 ( .A1(n715), .A2(n702), .ZN(n629) );
  NAND2_X1 U532 ( .A1(n412), .A2(n414), .ZN(n413) );
  NAND2_X1 U533 ( .A1(n416), .A2(KEYINPUT87), .ZN(n412) );
  NAND2_X1 U534 ( .A1(n419), .A2(n429), .ZN(n421) );
  XNOR2_X1 U535 ( .A(n422), .B(n619), .ZN(n637) );
  NAND2_X1 U536 ( .A1(n441), .A2(n436), .ZN(n430) );
  INV_X1 U537 ( .A(n418), .ZN(n416) );
  XNOR2_X1 U538 ( .A(n442), .B(n445), .ZN(n418) );
  NAND2_X1 U539 ( .A1(n418), .A2(n415), .ZN(n414) );
  NAND2_X1 U540 ( .A1(n444), .A2(KEYINPUT87), .ZN(n415) );
  NAND2_X1 U541 ( .A1(n406), .A2(n431), .ZN(n420) );
  NAND2_X1 U542 ( .A1(n431), .A2(n430), .ZN(n419) );
  INV_X1 U543 ( .A(n478), .ZN(n423) );
  XNOR2_X2 U544 ( .A(n523), .B(n372), .ZN(n461) );
  NAND2_X1 U545 ( .A1(n647), .A2(KEYINPUT44), .ZN(n641) );
  NAND2_X1 U546 ( .A1(n427), .A2(n652), .ZN(n654) );
  XNOR2_X1 U547 ( .A(n428), .B(KEYINPUT86), .ZN(n427) );
  NAND2_X1 U548 ( .A1(n438), .A2(n437), .ZN(n431) );
  AND2_X1 U549 ( .A1(n618), .A2(n374), .ZN(n437) );
  NAND2_X1 U550 ( .A1(n439), .A2(n440), .ZN(n438) );
  INV_X1 U551 ( .A(n760), .ZN(n439) );
  INV_X1 U552 ( .A(n616), .ZN(n440) );
  NAND2_X1 U553 ( .A1(n607), .A2(n606), .ZN(n442) );
  INV_X1 U554 ( .A(n608), .ZN(n444) );
  INV_X1 U555 ( .A(n756), .ZN(n454) );
  NAND2_X1 U556 ( .A1(n628), .A2(n591), .ZN(n455) );
  XNOR2_X1 U557 ( .A(n756), .B(n587), .ZN(n628) );
  XNOR2_X2 U558 ( .A(n586), .B(n456), .ZN(n756) );
  BUF_X2 U559 ( .A(n539), .Z(n741) );
  INV_X1 U560 ( .A(n539), .ZN(n492) );
  XNOR2_X2 U561 ( .A(n701), .B(KEYINPUT106), .ZN(n585) );
  XNOR2_X1 U562 ( .A(n461), .B(n460), .ZN(n464) );
  BUF_X1 U563 ( .A(n686), .Z(n692) );
  NAND2_X1 U564 ( .A1(G234), .A2(n793), .ZN(n472) );
  INV_X1 U565 ( .A(n740), .ZN(n491) );
  XNOR2_X1 U566 ( .A(n781), .B(n511), .ZN(n668) );
  XNOR2_X1 U567 ( .A(n634), .B(KEYINPUT108), .ZN(n684) );
  NAND2_X1 U568 ( .A1(n517), .A2(G210), .ZN(n457) );
  XNOR2_X1 U569 ( .A(n457), .B(KEYINPUT76), .ZN(n459) );
  XNOR2_X1 U570 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X2 U571 ( .A(G113), .B(KEYINPUT70), .ZN(n462) );
  XNOR2_X1 U572 ( .A(n508), .B(G146), .ZN(n469) );
  XNOR2_X1 U573 ( .A(n501), .B(n469), .ZN(n463) );
  INV_X1 U574 ( .A(KEYINPUT102), .ZN(n465) );
  XNOR2_X1 U575 ( .A(KEYINPUT75), .B(n466), .ZN(n512) );
  AND2_X1 U576 ( .A1(n512), .A2(G214), .ZN(n552) );
  NAND2_X1 U577 ( .A1(n793), .A2(G227), .ZN(n467) );
  XNOR2_X1 U578 ( .A(n467), .B(KEYINPUT97), .ZN(n468) );
  XNOR2_X1 U579 ( .A(n500), .B(n468), .ZN(n470) );
  NAND2_X1 U580 ( .A1(n524), .A2(G221), .ZN(n475) );
  XNOR2_X1 U581 ( .A(KEYINPUT98), .B(KEYINPUT23), .ZN(n477) );
  NAND2_X1 U582 ( .A1(n479), .A2(n533), .ZN(n486) );
  NAND2_X1 U583 ( .A1(n610), .A2(G234), .ZN(n480) );
  XNOR2_X1 U584 ( .A(n480), .B(KEYINPUT20), .ZN(n487) );
  NAND2_X1 U585 ( .A1(n487), .A2(G217), .ZN(n484) );
  XNOR2_X1 U586 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n482) );
  INV_X1 U587 ( .A(KEYINPUT25), .ZN(n481) );
  XNOR2_X1 U588 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U589 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U590 ( .A(n486), .B(n485), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n487), .A2(G221), .ZN(n490) );
  INV_X1 U592 ( .A(KEYINPUT101), .ZN(n488) );
  XNOR2_X1 U593 ( .A(n488), .B(KEYINPUT21), .ZN(n489) );
  XNOR2_X1 U594 ( .A(n490), .B(n489), .ZN(n740) );
  NAND2_X1 U595 ( .A1(n492), .A2(n491), .ZN(n737) );
  XNOR2_X1 U596 ( .A(n493), .B(KEYINPUT14), .ZN(n497) );
  AND2_X1 U597 ( .A1(n798), .A2(G902), .ZN(n494) );
  NAND2_X1 U598 ( .A1(n497), .A2(n494), .ZN(n554) );
  XNOR2_X1 U599 ( .A(KEYINPUT111), .B(n554), .ZN(n496) );
  INV_X1 U600 ( .A(G900), .ZN(n495) );
  NAND2_X1 U601 ( .A1(n496), .A2(n495), .ZN(n498) );
  NAND2_X1 U602 ( .A1(G952), .A2(n497), .ZN(n768) );
  OR2_X1 U603 ( .A1(n768), .A2(n798), .ZN(n557) );
  NAND2_X1 U604 ( .A1(n498), .A2(n557), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n503), .B(n502), .ZN(n507) );
  NAND2_X1 U606 ( .A1(n793), .A2(G224), .ZN(n504) );
  XNOR2_X1 U607 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U608 ( .A(n507), .B(n506), .ZN(n510) );
  XNOR2_X1 U609 ( .A(n405), .B(n508), .ZN(n509) );
  XNOR2_X1 U610 ( .A(n510), .B(n509), .ZN(n511) );
  INV_X1 U611 ( .A(n610), .ZN(n651) );
  AND2_X1 U612 ( .A1(n512), .A2(G210), .ZN(n513) );
  XNOR2_X1 U613 ( .A(n513), .B(KEYINPUT95), .ZN(n514) );
  NOR2_X1 U614 ( .A1(n595), .A2(n572), .ZN(n515) );
  XNOR2_X1 U615 ( .A(n515), .B(KEYINPUT39), .ZN(n570) );
  BUF_X1 U616 ( .A(n570), .Z(n516) );
  INV_X1 U617 ( .A(n516), .ZN(n536) );
  NAND2_X1 U618 ( .A1(n517), .A2(G214), .ZN(n518) );
  NAND2_X1 U619 ( .A1(n660), .A2(n533), .ZN(n522) );
  XNOR2_X1 U620 ( .A(KEYINPUT13), .B(G475), .ZN(n521) );
  XNOR2_X2 U621 ( .A(n522), .B(n521), .ZN(n593) );
  XNOR2_X1 U622 ( .A(n593), .B(KEYINPUT104), .ZN(n538) );
  NAND2_X1 U623 ( .A1(n524), .A2(G217), .ZN(n525) );
  XNOR2_X1 U624 ( .A(n528), .B(n527), .ZN(n530) );
  XNOR2_X1 U625 ( .A(n530), .B(n529), .ZN(n531) );
  NAND2_X1 U626 ( .A1(n680), .A2(n533), .ZN(n535) );
  INV_X1 U627 ( .A(G478), .ZN(n534) );
  INV_X1 U628 ( .A(n592), .ZN(n537) );
  AND2_X2 U629 ( .A1(n538), .A2(n537), .ZN(n701) );
  NAND2_X1 U630 ( .A1(n536), .A2(n585), .ZN(n609) );
  XNOR2_X1 U631 ( .A(n609), .B(G134), .ZN(G36) );
  XNOR2_X1 U632 ( .A(KEYINPUT43), .B(KEYINPUT113), .ZN(n549) );
  INV_X1 U633 ( .A(n575), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT6), .ZN(n631) );
  OR2_X1 U635 ( .A1(n538), .A2(n537), .ZN(n584) );
  INV_X1 U636 ( .A(n540), .ZN(n541) );
  NOR2_X1 U637 ( .A1(n740), .A2(n541), .ZN(n542) );
  NOR2_X1 U638 ( .A1(n631), .A2(n543), .ZN(n544) );
  XNOR2_X1 U639 ( .A(n544), .B(KEYINPUT112), .ZN(n545) );
  INV_X1 U640 ( .A(n552), .ZN(n751) );
  AND2_X1 U641 ( .A1(n545), .A2(n751), .ZN(n600) );
  INV_X1 U642 ( .A(n600), .ZN(n547) );
  XOR2_X1 U643 ( .A(n549), .B(n548), .Z(n550) );
  INV_X1 U644 ( .A(n551), .ZN(n599) );
  XOR2_X1 U645 ( .A(G140), .B(n608), .Z(G42) );
  XNOR2_X1 U646 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n553) );
  NOR2_X1 U647 ( .A1(G898), .A2(n554), .ZN(n556) );
  INV_X1 U648 ( .A(KEYINPUT96), .ZN(n555) );
  XNOR2_X1 U649 ( .A(n556), .B(n555), .ZN(n558) );
  NAND2_X1 U650 ( .A1(n558), .A2(n557), .ZN(n559) );
  INV_X1 U651 ( .A(KEYINPUT68), .ZN(n560) );
  XNOR2_X1 U652 ( .A(n560), .B(KEYINPUT0), .ZN(n561) );
  NAND2_X1 U653 ( .A1(n593), .A2(n592), .ZN(n754) );
  XNOR2_X1 U654 ( .A(KEYINPUT72), .B(KEYINPUT22), .ZN(n562) );
  XNOR2_X1 U655 ( .A(n562), .B(KEYINPUT67), .ZN(n563) );
  INV_X1 U656 ( .A(n741), .ZN(n630) );
  INV_X1 U657 ( .A(KEYINPUT110), .ZN(n566) );
  XNOR2_X1 U658 ( .A(n366), .B(n566), .ZN(n569) );
  INV_X1 U659 ( .A(n567), .ZN(n743) );
  AND2_X1 U660 ( .A1(n743), .A2(n741), .ZN(n568) );
  NAND2_X1 U661 ( .A1(n569), .A2(n568), .ZN(n640) );
  XNOR2_X1 U662 ( .A(n640), .B(G110), .ZN(G12) );
  NOR2_X1 U663 ( .A1(n570), .A2(n584), .ZN(n571) );
  XNOR2_X1 U664 ( .A(n571), .B(KEYINPUT40), .ZN(n685) );
  INV_X1 U665 ( .A(n572), .ZN(n752) );
  NAND2_X1 U666 ( .A1(n752), .A2(n751), .ZN(n755) );
  XNOR2_X1 U667 ( .A(KEYINPUT41), .B(n573), .ZN(n769) );
  INV_X1 U668 ( .A(KEYINPUT28), .ZN(n576) );
  XNOR2_X1 U669 ( .A(n577), .B(n576), .ZN(n578) );
  NAND2_X1 U670 ( .A1(n626), .A2(n578), .ZN(n588) );
  NOR2_X1 U671 ( .A1(n769), .A2(n588), .ZN(n580) );
  XNOR2_X1 U672 ( .A(KEYINPUT114), .B(KEYINPUT42), .ZN(n579) );
  XNOR2_X1 U673 ( .A(KEYINPUT88), .B(KEYINPUT46), .ZN(n581) );
  XNOR2_X1 U674 ( .A(n581), .B(KEYINPUT64), .ZN(n582) );
  XNOR2_X1 U675 ( .A(n583), .B(n582), .ZN(n607) );
  INV_X1 U676 ( .A(n584), .ZN(n712) );
  NOR2_X2 U677 ( .A1(n712), .A2(n585), .ZN(n586) );
  INV_X1 U678 ( .A(KEYINPUT82), .ZN(n587) );
  INV_X1 U679 ( .A(n588), .ZN(n590) );
  NAND2_X1 U680 ( .A1(n590), .A2(n589), .ZN(n707) );
  NOR2_X1 U681 ( .A1(n707), .A2(KEYINPUT47), .ZN(n591) );
  OR2_X1 U682 ( .A1(n593), .A2(n592), .ZN(n617) );
  OR2_X1 U683 ( .A1(n551), .A2(n617), .ZN(n594) );
  NOR2_X1 U684 ( .A1(n595), .A2(n594), .ZN(n710) );
  XOR2_X1 U685 ( .A(KEYINPUT83), .B(n710), .Z(n596) );
  NOR2_X1 U686 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U687 ( .A(n598), .B(KEYINPUT73), .ZN(n605) );
  NAND2_X1 U688 ( .A1(n600), .A2(n599), .ZN(n602) );
  INV_X1 U689 ( .A(KEYINPUT36), .ZN(n601) );
  XNOR2_X1 U690 ( .A(n602), .B(n601), .ZN(n604) );
  AND2_X1 U691 ( .A1(n604), .A2(n603), .ZN(n717) );
  XNOR2_X1 U692 ( .A(n655), .B(KEYINPUT78), .ZN(n611) );
  NAND2_X1 U693 ( .A1(n612), .A2(n624), .ZN(n613) );
  XNOR2_X1 U694 ( .A(n613), .B(KEYINPUT74), .ZN(n620) );
  OR2_X2 U695 ( .A1(n620), .A2(n631), .ZN(n615) );
  INV_X1 U696 ( .A(KEYINPUT33), .ZN(n614) );
  XNOR2_X2 U697 ( .A(n615), .B(n614), .ZN(n760) );
  INV_X1 U698 ( .A(n622), .ZN(n616) );
  INV_X1 U699 ( .A(n617), .ZN(n618) );
  INV_X1 U700 ( .A(KEYINPUT91), .ZN(n619) );
  OR2_X1 U701 ( .A1(n620), .A2(n743), .ZN(n621) );
  XNOR2_X1 U702 ( .A(n621), .B(KEYINPUT103), .ZN(n748) );
  NAND2_X1 U703 ( .A1(n748), .A2(n440), .ZN(n623) );
  XNOR2_X1 U704 ( .A(n623), .B(KEYINPUT31), .ZN(n715) );
  AND2_X1 U705 ( .A1(n743), .A2(n624), .ZN(n625) );
  AND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U707 ( .A1(n440), .A2(n627), .ZN(n702) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n635) );
  AND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n634) );
  AND2_X1 U711 ( .A1(n635), .A2(n684), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n639) );
  INV_X1 U713 ( .A(KEYINPUT90), .ZN(n638) );
  BUF_X1 U714 ( .A(n642), .Z(n643) );
  INV_X1 U715 ( .A(n643), .ZN(n645) );
  INV_X1 U716 ( .A(KEYINPUT44), .ZN(n644) );
  AND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n649) );
  INV_X1 U718 ( .A(KEYINPUT92), .ZN(n646) );
  XNOR2_X1 U719 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U720 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n651), .A2(KEYINPUT2), .ZN(n652) );
  INV_X1 U722 ( .A(KEYINPUT65), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n654), .B(n653), .ZN(n659) );
  BUF_X1 U724 ( .A(n655), .Z(n792) );
  INV_X1 U725 ( .A(n792), .ZN(n729) );
  NAND2_X1 U726 ( .A1(n729), .A2(KEYINPUT2), .ZN(n657) );
  INV_X1 U727 ( .A(n776), .ZN(n730) );
  NOR2_X1 U728 ( .A1(n657), .A2(n730), .ZN(n734) );
  INV_X1 U729 ( .A(n734), .ZN(n658) );
  AND2_X2 U730 ( .A1(n659), .A2(n658), .ZN(n686) );
  NAND2_X1 U731 ( .A1(n686), .A2(G475), .ZN(n662) );
  XNOR2_X1 U732 ( .A(n662), .B(n661), .ZN(n664) );
  INV_X1 U733 ( .A(G952), .ZN(n663) );
  NAND2_X1 U734 ( .A1(n664), .A2(n690), .ZN(n666) );
  INV_X1 U735 ( .A(KEYINPUT60), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n666), .B(n665), .ZN(G60) );
  NAND2_X1 U737 ( .A1(n686), .A2(G210), .ZN(n670) );
  XNOR2_X1 U738 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U740 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U741 ( .A1(n671), .A2(n690), .ZN(n673) );
  XOR2_X1 U742 ( .A(KEYINPUT120), .B(KEYINPUT56), .Z(n672) );
  XNOR2_X1 U743 ( .A(n673), .B(n672), .ZN(G51) );
  NAND2_X1 U744 ( .A1(n686), .A2(G472), .ZN(n676) );
  XNOR2_X1 U745 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U746 ( .A1(n677), .A2(n690), .ZN(n679) );
  XOR2_X1 U747 ( .A(KEYINPUT115), .B(KEYINPUT63), .Z(n678) );
  XNOR2_X1 U748 ( .A(n679), .B(n678), .ZN(G57) );
  NAND2_X1 U749 ( .A1(n686), .A2(G478), .ZN(n681) );
  XNOR2_X1 U750 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U751 ( .A1(n682), .A2(n690), .ZN(n683) );
  XNOR2_X1 U752 ( .A(n683), .B(KEYINPUT121), .ZN(G63) );
  XNOR2_X1 U753 ( .A(n684), .B(G101), .ZN(G3) );
  XOR2_X1 U754 ( .A(n409), .B(G131), .Z(G33) );
  XOR2_X1 U755 ( .A(n643), .B(G122), .Z(G24) );
  NAND2_X1 U756 ( .A1(n692), .A2(G217), .ZN(n689) );
  XNOR2_X1 U757 ( .A(n687), .B(KEYINPUT122), .ZN(n688) );
  XNOR2_X1 U758 ( .A(n689), .B(n688), .ZN(n691) );
  INV_X1 U759 ( .A(n690), .ZN(n698) );
  NOR2_X1 U760 ( .A1(n691), .A2(n698), .ZN(G66) );
  NAND2_X1 U761 ( .A1(n692), .A2(G469), .ZN(n697) );
  BUF_X1 U762 ( .A(n693), .Z(n695) );
  XOR2_X1 U763 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n694) );
  XNOR2_X1 U764 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U765 ( .A(n697), .B(n696), .ZN(n699) );
  NOR2_X1 U766 ( .A1(n699), .A2(n698), .ZN(G54) );
  NAND2_X1 U767 ( .A1(n702), .A2(n712), .ZN(n700) );
  XNOR2_X1 U768 ( .A(n700), .B(G104), .ZN(G6) );
  XOR2_X1 U769 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n704) );
  NAND2_X1 U770 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U771 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U772 ( .A(G107), .B(n705), .ZN(G9) );
  XOR2_X1 U773 ( .A(G128), .B(KEYINPUT29), .Z(n709) );
  NAND2_X1 U774 ( .A1(n389), .A2(n701), .ZN(n708) );
  XNOR2_X1 U775 ( .A(n709), .B(n708), .ZN(G30) );
  XOR2_X1 U776 ( .A(G143), .B(n710), .Z(G45) );
  NAND2_X1 U777 ( .A1(n389), .A2(n712), .ZN(n711) );
  XNOR2_X1 U778 ( .A(n711), .B(G146), .ZN(G48) );
  NAND2_X1 U779 ( .A1(n715), .A2(n712), .ZN(n713) );
  XNOR2_X1 U780 ( .A(n713), .B(KEYINPUT116), .ZN(n714) );
  XNOR2_X1 U781 ( .A(G113), .B(n714), .ZN(G15) );
  NAND2_X1 U782 ( .A1(n715), .A2(n701), .ZN(n716) );
  XNOR2_X1 U783 ( .A(n716), .B(G116), .ZN(G18) );
  XOR2_X1 U784 ( .A(KEYINPUT37), .B(KEYINPUT117), .Z(n719) );
  XNOR2_X1 U785 ( .A(G125), .B(n717), .ZN(n718) );
  XNOR2_X1 U786 ( .A(n719), .B(n718), .ZN(G27) );
  NOR2_X1 U787 ( .A1(n729), .A2(KEYINPUT85), .ZN(n721) );
  XNOR2_X1 U788 ( .A(KEYINPUT2), .B(KEYINPUT81), .ZN(n726) );
  INV_X1 U789 ( .A(n726), .ZN(n720) );
  NOR2_X1 U790 ( .A1(n721), .A2(n720), .ZN(n723) );
  NAND2_X1 U791 ( .A1(n730), .A2(KEYINPUT84), .ZN(n722) );
  NAND2_X1 U792 ( .A1(n723), .A2(n722), .ZN(n728) );
  INV_X1 U793 ( .A(KEYINPUT85), .ZN(n724) );
  NAND2_X1 U794 ( .A1(n724), .A2(KEYINPUT84), .ZN(n725) );
  OR2_X1 U795 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U796 ( .A1(n728), .A2(n727), .ZN(n736) );
  NAND2_X1 U797 ( .A1(n729), .A2(KEYINPUT85), .ZN(n732) );
  OR2_X1 U798 ( .A1(n730), .A2(KEYINPUT84), .ZN(n731) );
  NAND2_X1 U799 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U800 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U801 ( .A1(n736), .A2(n735), .ZN(n773) );
  NAND2_X1 U802 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U803 ( .A(KEYINPUT50), .B(n739), .Z(n746) );
  NAND2_X1 U804 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U805 ( .A(KEYINPUT49), .B(n742), .Z(n744) );
  NAND2_X1 U806 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U807 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U808 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U809 ( .A(KEYINPUT51), .B(n749), .Z(n750) );
  NOR2_X1 U810 ( .A1(n769), .A2(n750), .ZN(n765) );
  NOR2_X1 U811 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U812 ( .A1(n754), .A2(n753), .ZN(n759) );
  NOR2_X1 U813 ( .A1(n364), .A2(n755), .ZN(n757) );
  XNOR2_X1 U814 ( .A(n757), .B(KEYINPUT118), .ZN(n758) );
  NOR2_X1 U815 ( .A1(n759), .A2(n758), .ZN(n762) );
  BUF_X1 U816 ( .A(n760), .Z(n761) );
  NOR2_X1 U817 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U818 ( .A(KEYINPUT119), .B(n763), .Z(n764) );
  NOR2_X1 U819 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U820 ( .A(n766), .B(KEYINPUT52), .ZN(n767) );
  NOR2_X1 U821 ( .A1(n768), .A2(n767), .ZN(n771) );
  NOR2_X1 U822 ( .A1(n769), .A2(n761), .ZN(n770) );
  NOR2_X1 U823 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U824 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U825 ( .A1(n774), .A2(n798), .ZN(n775) );
  XNOR2_X1 U826 ( .A(n775), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U827 ( .A1(n776), .A2(n793), .ZN(n780) );
  NAND2_X1 U828 ( .A1(n798), .A2(G224), .ZN(n777) );
  XNOR2_X1 U829 ( .A(KEYINPUT61), .B(n777), .ZN(n778) );
  NAND2_X1 U830 ( .A1(n778), .A2(G898), .ZN(n779) );
  NAND2_X1 U831 ( .A1(n780), .A2(n779), .ZN(n788) );
  NOR2_X1 U832 ( .A1(G898), .A2(n793), .ZN(n784) );
  XOR2_X1 U833 ( .A(G101), .B(KEYINPUT124), .Z(n782) );
  XNOR2_X1 U834 ( .A(n781), .B(n782), .ZN(n783) );
  NOR2_X1 U835 ( .A1(n784), .A2(n783), .ZN(n786) );
  XNOR2_X1 U836 ( .A(KEYINPUT123), .B(KEYINPUT125), .ZN(n785) );
  XNOR2_X1 U837 ( .A(n786), .B(n785), .ZN(n787) );
  XNOR2_X1 U838 ( .A(n788), .B(n787), .ZN(G69) );
  BUF_X1 U839 ( .A(n789), .Z(n790) );
  XNOR2_X1 U840 ( .A(n790), .B(n365), .ZN(n796) );
  XNOR2_X1 U841 ( .A(n792), .B(n796), .ZN(n794) );
  NAND2_X1 U842 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U843 ( .A(n795), .B(KEYINPUT126), .ZN(n801) );
  XNOR2_X1 U844 ( .A(n796), .B(G227), .ZN(n797) );
  NAND2_X1 U845 ( .A1(n797), .A2(G900), .ZN(n799) );
  NAND2_X1 U846 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U847 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U848 ( .A(KEYINPUT127), .B(n802), .Z(G72) );
  XOR2_X1 U849 ( .A(G137), .B(n803), .Z(G39) );
endmodule

