

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U555 ( .A(n726), .ZN(n706) );
  XNOR2_X2 U556 ( .A(n534), .B(KEYINPUT67), .ZN(n649) );
  XNOR2_X2 U557 ( .A(G543), .B(KEYINPUT0), .ZN(n534) );
  OR2_X2 U558 ( .A1(n682), .A2(n761), .ZN(n726) );
  NOR2_X1 U559 ( .A1(n719), .A2(n718), .ZN(n721) );
  AND2_X1 U560 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X2 U561 ( .A1(G651), .A2(G543), .ZN(n639) );
  XNOR2_X1 U562 ( .A(KEYINPUT32), .B(KEYINPUT97), .ZN(n522) );
  NAND2_X1 U563 ( .A1(n775), .A2(n774), .ZN(n523) );
  XOR2_X1 U564 ( .A(KEYINPUT87), .B(n763), .Z(n524) );
  INV_X1 U565 ( .A(KEYINPUT31), .ZN(n720) );
  XNOR2_X1 U566 ( .A(n734), .B(n522), .ZN(n741) );
  INV_X1 U567 ( .A(n954), .ZN(n744) );
  NOR2_X1 U568 ( .A1(n772), .A2(n744), .ZN(n745) );
  NAND2_X1 U569 ( .A1(G8), .A2(n726), .ZN(n772) );
  NOR2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  NOR2_X1 U571 ( .A1(G164), .A2(G1384), .ZN(n762) );
  XNOR2_X1 U572 ( .A(n577), .B(KEYINPUT75), .ZN(n578) );
  NOR2_X1 U573 ( .A1(n649), .A2(n538), .ZN(n640) );
  NOR2_X1 U574 ( .A1(G651), .A2(n649), .ZN(n648) );
  INV_X1 U575 ( .A(n603), .ZN(n686) );
  INV_X1 U576 ( .A(G2105), .ZN(n529) );
  AND2_X1 U577 ( .A1(n529), .A2(G2104), .ZN(n880) );
  NAND2_X1 U578 ( .A1(G102), .A2(n880), .ZN(n528) );
  XOR2_X1 U579 ( .A(KEYINPUT66), .B(n525), .Z(n526) );
  XNOR2_X2 U580 ( .A(n526), .B(KEYINPUT17), .ZN(n872) );
  NAND2_X1 U581 ( .A1(G138), .A2(n872), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n528), .A2(n527), .ZN(n533) );
  AND2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n874) );
  NAND2_X1 U584 ( .A1(G114), .A2(n874), .ZN(n531) );
  NOR2_X1 U585 ( .A1(G2104), .A2(n529), .ZN(n875) );
  NAND2_X1 U586 ( .A1(G126), .A2(n875), .ZN(n530) );
  NAND2_X1 U587 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U588 ( .A1(n533), .A2(n532), .ZN(G164) );
  AND2_X1 U589 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U590 ( .A1(G52), .A2(n648), .ZN(n537) );
  INV_X1 U591 ( .A(G651), .ZN(n538) );
  NOR2_X1 U592 ( .A1(G543), .A2(n538), .ZN(n535) );
  XOR2_X1 U593 ( .A(KEYINPUT1), .B(n535), .Z(n653) );
  NAND2_X1 U594 ( .A1(G64), .A2(n653), .ZN(n536) );
  NAND2_X1 U595 ( .A1(n537), .A2(n536), .ZN(n545) );
  XNOR2_X1 U596 ( .A(KEYINPUT70), .B(KEYINPUT9), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n640), .A2(G77), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n639), .A2(G90), .ZN(n539) );
  XOR2_X1 U599 ( .A(KEYINPUT69), .B(n539), .Z(n540) );
  NAND2_X1 U600 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U601 ( .A(n543), .B(n542), .Z(n544) );
  NOR2_X1 U602 ( .A1(n545), .A2(n544), .ZN(G171) );
  INV_X1 U603 ( .A(G171), .ZN(G301) );
  INV_X1 U604 ( .A(G57), .ZN(G237) );
  NAND2_X1 U605 ( .A1(G101), .A2(n880), .ZN(n546) );
  XOR2_X1 U606 ( .A(KEYINPUT23), .B(n546), .Z(n549) );
  NAND2_X1 U607 ( .A1(G113), .A2(n874), .ZN(n547) );
  XOR2_X1 U608 ( .A(KEYINPUT65), .B(n547), .Z(n548) );
  NAND2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n875), .A2(G125), .ZN(n551) );
  NAND2_X1 U611 ( .A1(G137), .A2(n872), .ZN(n550) );
  NAND2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U613 ( .A1(n553), .A2(n552), .ZN(G160) );
  NAND2_X1 U614 ( .A1(n639), .A2(G89), .ZN(n554) );
  XNOR2_X1 U615 ( .A(n554), .B(KEYINPUT4), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G76), .A2(n640), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U618 ( .A(n557), .B(KEYINPUT5), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n653), .A2(G63), .ZN(n558) );
  XNOR2_X1 U620 ( .A(n558), .B(KEYINPUT78), .ZN(n560) );
  NAND2_X1 U621 ( .A1(G51), .A2(n648), .ZN(n559) );
  NAND2_X1 U622 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT6), .B(n561), .Z(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U625 ( .A(n564), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U626 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U627 ( .A1(G7), .A2(G661), .ZN(n565) );
  XOR2_X1 U628 ( .A(n565), .B(KEYINPUT10), .Z(n817) );
  NAND2_X1 U629 ( .A1(n817), .A2(G567), .ZN(n566) );
  XNOR2_X1 U630 ( .A(n566), .B(KEYINPUT73), .ZN(n567) );
  XNOR2_X1 U631 ( .A(KEYINPUT11), .B(n567), .ZN(G234) );
  NAND2_X1 U632 ( .A1(n648), .A2(G43), .ZN(n568) );
  XNOR2_X1 U633 ( .A(KEYINPUT76), .B(n568), .ZN(n579) );
  NAND2_X1 U634 ( .A1(n653), .A2(G56), .ZN(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT14), .B(n569), .ZN(n576) );
  NAND2_X1 U636 ( .A1(G81), .A2(n639), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(KEYINPUT12), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT74), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G68), .A2(n640), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(KEYINPUT13), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n603) );
  NAND2_X1 U644 ( .A1(n686), .A2(G860), .ZN(G153) );
  NAND2_X1 U645 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U646 ( .A1(G66), .A2(n653), .ZN(n586) );
  NAND2_X1 U647 ( .A1(G79), .A2(n640), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G54), .A2(n648), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U650 ( .A1(G92), .A2(n639), .ZN(n582) );
  XNOR2_X1 U651 ( .A(KEYINPUT77), .B(n582), .ZN(n583) );
  NOR2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U654 ( .A(n587), .B(KEYINPUT15), .Z(n946) );
  INV_X1 U655 ( .A(G868), .ZN(n664) );
  NAND2_X1 U656 ( .A1(n946), .A2(n664), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U658 ( .A1(G53), .A2(n648), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G65), .A2(n653), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G91), .A2(n639), .ZN(n593) );
  NAND2_X1 U662 ( .A1(G78), .A2(n640), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U665 ( .A(KEYINPUT71), .B(n596), .Z(n952) );
  XOR2_X1 U666 ( .A(n952), .B(KEYINPUT72), .Z(G299) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U668 ( .A1(G286), .A2(n664), .ZN(n597) );
  NOR2_X1 U669 ( .A1(n598), .A2(n597), .ZN(G297) );
  INV_X1 U670 ( .A(G559), .ZN(n599) );
  NOR2_X1 U671 ( .A1(G860), .A2(n599), .ZN(n600) );
  XNOR2_X1 U672 ( .A(KEYINPUT79), .B(n600), .ZN(n601) );
  INV_X1 U673 ( .A(n946), .ZN(n891) );
  NAND2_X1 U674 ( .A1(n601), .A2(n891), .ZN(n602) );
  XNOR2_X1 U675 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U676 ( .A1(G868), .A2(n603), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G868), .A2(n891), .ZN(n604) );
  NOR2_X1 U678 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U679 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U680 ( .A1(G99), .A2(n880), .ZN(n608) );
  NAND2_X1 U681 ( .A1(G111), .A2(n874), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U683 ( .A(KEYINPUT80), .B(n609), .ZN(n614) );
  NAND2_X1 U684 ( .A1(G123), .A2(n875), .ZN(n610) );
  XNOR2_X1 U685 ( .A(n610), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U686 ( .A1(G135), .A2(n872), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U688 ( .A1(n614), .A2(n613), .ZN(n918) );
  XNOR2_X1 U689 ( .A(n918), .B(G2096), .ZN(n615) );
  INV_X1 U690 ( .A(G2100), .ZN(n835) );
  NAND2_X1 U691 ( .A1(n615), .A2(n835), .ZN(G156) );
  NAND2_X1 U692 ( .A1(G559), .A2(n891), .ZN(n616) );
  XOR2_X1 U693 ( .A(n616), .B(n686), .Z(n662) );
  NOR2_X1 U694 ( .A1(n662), .A2(G860), .ZN(n623) );
  NAND2_X1 U695 ( .A1(G55), .A2(n648), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G67), .A2(n653), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G93), .A2(n639), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G80), .A2(n640), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n665) );
  XNOR2_X1 U702 ( .A(n623), .B(n665), .ZN(G145) );
  NAND2_X1 U703 ( .A1(n639), .A2(G86), .ZN(n630) );
  NAND2_X1 U704 ( .A1(G48), .A2(n648), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G61), .A2(n653), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n640), .A2(G73), .ZN(n626) );
  XOR2_X1 U708 ( .A(KEYINPUT2), .B(n626), .Z(n627) );
  NOR2_X1 U709 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U711 ( .A(KEYINPUT81), .B(n631), .Z(G305) );
  NAND2_X1 U712 ( .A1(G85), .A2(n639), .ZN(n633) );
  NAND2_X1 U713 ( .A1(G72), .A2(n640), .ZN(n632) );
  NAND2_X1 U714 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U715 ( .A1(G60), .A2(n653), .ZN(n634) );
  XOR2_X1 U716 ( .A(KEYINPUT68), .B(n634), .Z(n635) );
  NOR2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U718 ( .A1(n648), .A2(G47), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n638), .A2(n637), .ZN(G290) );
  NAND2_X1 U720 ( .A1(G88), .A2(n639), .ZN(n642) );
  NAND2_X1 U721 ( .A1(G75), .A2(n640), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n647) );
  NAND2_X1 U723 ( .A1(G62), .A2(n653), .ZN(n643) );
  XNOR2_X1 U724 ( .A(n643), .B(KEYINPUT82), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n648), .A2(G50), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U727 ( .A1(n647), .A2(n646), .ZN(G166) );
  NAND2_X1 U728 ( .A1(G49), .A2(n648), .ZN(n651) );
  NAND2_X1 U729 ( .A1(G87), .A2(n649), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U732 ( .A1(G651), .A2(G74), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n655), .A2(n654), .ZN(G288) );
  XNOR2_X1 U734 ( .A(n665), .B(KEYINPUT19), .ZN(n656) );
  XNOR2_X1 U735 ( .A(n656), .B(KEYINPUT83), .ZN(n659) );
  XOR2_X1 U736 ( .A(G166), .B(G299), .Z(n657) );
  XNOR2_X1 U737 ( .A(G290), .B(n657), .ZN(n658) );
  XNOR2_X1 U738 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U739 ( .A(n660), .B(G288), .ZN(n661) );
  XNOR2_X1 U740 ( .A(G305), .B(n661), .ZN(n894) );
  XNOR2_X1 U741 ( .A(n662), .B(n894), .ZN(n663) );
  NAND2_X1 U742 ( .A1(n663), .A2(G868), .ZN(n667) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U744 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U745 ( .A(KEYINPUT84), .B(n668), .Z(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U750 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U752 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n674) );
  NAND2_X1 U753 ( .A1(G132), .A2(G82), .ZN(n673) );
  XNOR2_X1 U754 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U755 ( .A1(n675), .A2(G218), .ZN(n676) );
  NAND2_X1 U756 ( .A1(G96), .A2(n676), .ZN(n822) );
  NAND2_X1 U757 ( .A1(n822), .A2(G2106), .ZN(n680) );
  NAND2_X1 U758 ( .A1(G69), .A2(G120), .ZN(n677) );
  NOR2_X1 U759 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U760 ( .A1(G108), .A2(n678), .ZN(n821) );
  NAND2_X1 U761 ( .A1(n821), .A2(G567), .ZN(n679) );
  NAND2_X1 U762 ( .A1(n680), .A2(n679), .ZN(n844) );
  NAND2_X1 U763 ( .A1(G483), .A2(G661), .ZN(n681) );
  NOR2_X1 U764 ( .A1(n844), .A2(n681), .ZN(n820) );
  NAND2_X1 U765 ( .A1(n820), .A2(G36), .ZN(G176) );
  XOR2_X1 U766 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  INV_X1 U767 ( .A(n762), .ZN(n682) );
  NAND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n761) );
  NOR2_X1 U769 ( .A1(n706), .A2(G1348), .ZN(n684) );
  NOR2_X1 U770 ( .A1(G2067), .A2(n726), .ZN(n683) );
  NOR2_X1 U771 ( .A1(n684), .A2(n683), .ZN(n692) );
  NAND2_X1 U772 ( .A1(n692), .A2(n946), .ZN(n691) );
  INV_X1 U773 ( .A(G1996), .ZN(n824) );
  NOR2_X1 U774 ( .A1(n726), .A2(n824), .ZN(n685) );
  XNOR2_X1 U775 ( .A(n685), .B(KEYINPUT26), .ZN(n689) );
  NAND2_X1 U776 ( .A1(n726), .A2(G1341), .ZN(n687) );
  NAND2_X1 U777 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U778 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U779 ( .A1(n691), .A2(n690), .ZN(n694) );
  OR2_X1 U780 ( .A1(n692), .A2(n946), .ZN(n693) );
  NAND2_X1 U781 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U782 ( .A(KEYINPUT94), .B(n695), .Z(n700) );
  NAND2_X1 U783 ( .A1(n706), .A2(G2072), .ZN(n696) );
  XNOR2_X1 U784 ( .A(n696), .B(KEYINPUT27), .ZN(n698) );
  INV_X1 U785 ( .A(G1956), .ZN(n951) );
  NOR2_X1 U786 ( .A1(n951), .A2(n706), .ZN(n697) );
  NOR2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U788 ( .A1(n701), .A2(n952), .ZN(n699) );
  NAND2_X1 U789 ( .A1(n700), .A2(n699), .ZN(n704) );
  NOR2_X1 U790 ( .A1(n701), .A2(n952), .ZN(n702) );
  XOR2_X1 U791 ( .A(n702), .B(KEYINPUT28), .Z(n703) );
  NAND2_X1 U792 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U793 ( .A(KEYINPUT29), .B(n705), .Z(n710) );
  XNOR2_X1 U794 ( .A(G1961), .B(KEYINPUT93), .ZN(n985) );
  NAND2_X1 U795 ( .A1(n726), .A2(n985), .ZN(n708) );
  XNOR2_X1 U796 ( .A(G2078), .B(KEYINPUT25), .ZN(n998) );
  NAND2_X1 U797 ( .A1(n706), .A2(n998), .ZN(n707) );
  NAND2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n717) );
  NAND2_X1 U799 ( .A1(n717), .A2(G171), .ZN(n709) );
  NAND2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n723) );
  INV_X1 U801 ( .A(KEYINPUT92), .ZN(n712) );
  NOR2_X1 U802 ( .A1(G1966), .A2(n772), .ZN(n711) );
  XNOR2_X1 U803 ( .A(n712), .B(n711), .ZN(n736) );
  INV_X1 U804 ( .A(G8), .ZN(n731) );
  NOR2_X1 U805 ( .A1(G2084), .A2(n726), .ZN(n735) );
  NOR2_X1 U806 ( .A1(n731), .A2(n735), .ZN(n713) );
  AND2_X1 U807 ( .A1(n736), .A2(n713), .ZN(n715) );
  XNOR2_X1 U808 ( .A(KEYINPUT30), .B(KEYINPUT95), .ZN(n714) );
  XNOR2_X1 U809 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U810 ( .A1(n716), .A2(G168), .ZN(n719) );
  NOR2_X1 U811 ( .A1(G171), .A2(n717), .ZN(n718) );
  XNOR2_X1 U812 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n737) );
  AND2_X1 U814 ( .A1(G286), .A2(G8), .ZN(n724) );
  NAND2_X1 U815 ( .A1(n737), .A2(n724), .ZN(n733) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n772), .ZN(n725) );
  XNOR2_X1 U817 ( .A(n725), .B(KEYINPUT96), .ZN(n728) );
  NOR2_X1 U818 ( .A1(n726), .A2(G2090), .ZN(n727) );
  NOR2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n729), .A2(G303), .ZN(n730) );
  OR2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U822 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U823 ( .A1(G8), .A2(n735), .ZN(n739) );
  AND2_X1 U824 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U825 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U826 ( .A1(n741), .A2(n740), .ZN(n770) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n953) );
  NOR2_X1 U828 ( .A1(G303), .A2(G1971), .ZN(n742) );
  NOR2_X1 U829 ( .A1(n953), .A2(n742), .ZN(n743) );
  NAND2_X1 U830 ( .A1(n770), .A2(n743), .ZN(n746) );
  NAND2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n954) );
  XNOR2_X1 U832 ( .A(n747), .B(KEYINPUT64), .ZN(n748) );
  NOR2_X1 U833 ( .A1(KEYINPUT33), .A2(n748), .ZN(n751) );
  NAND2_X1 U834 ( .A1(n953), .A2(KEYINPUT33), .ZN(n749) );
  NOR2_X1 U835 ( .A1(n749), .A2(n772), .ZN(n750) );
  NOR2_X1 U836 ( .A1(n751), .A2(n750), .ZN(n765) );
  XOR2_X1 U837 ( .A(G1981), .B(G305), .Z(n942) );
  XNOR2_X1 U838 ( .A(KEYINPUT37), .B(G2067), .ZN(n808) );
  NAND2_X1 U839 ( .A1(G104), .A2(n880), .ZN(n753) );
  NAND2_X1 U840 ( .A1(G140), .A2(n872), .ZN(n752) );
  NAND2_X1 U841 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U842 ( .A(KEYINPUT34), .B(n754), .ZN(n759) );
  NAND2_X1 U843 ( .A1(G116), .A2(n874), .ZN(n756) );
  NAND2_X1 U844 ( .A1(G128), .A2(n875), .ZN(n755) );
  NAND2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U846 ( .A(KEYINPUT35), .B(n757), .Z(n758) );
  NOR2_X1 U847 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U848 ( .A(KEYINPUT36), .B(n760), .ZN(n887) );
  NOR2_X1 U849 ( .A1(n808), .A2(n887), .ZN(n937) );
  NOR2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n810) );
  NAND2_X1 U851 ( .A1(n937), .A2(n810), .ZN(n763) );
  AND2_X1 U852 ( .A1(n942), .A2(n524), .ZN(n764) );
  NAND2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n777) );
  NOR2_X1 U854 ( .A1(G1981), .A2(G305), .ZN(n766) );
  XOR2_X1 U855 ( .A(n766), .B(KEYINPUT24), .Z(n767) );
  OR2_X1 U856 ( .A1(n772), .A2(n767), .ZN(n775) );
  NOR2_X1 U857 ( .A1(G2090), .A2(G303), .ZN(n768) );
  NAND2_X1 U858 ( .A1(G8), .A2(n768), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U860 ( .A(n771), .B(KEYINPUT98), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n524), .A2(n523), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n798) );
  NAND2_X1 U864 ( .A1(G107), .A2(n874), .ZN(n779) );
  NAND2_X1 U865 ( .A1(G119), .A2(n875), .ZN(n778) );
  NAND2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U867 ( .A(KEYINPUT88), .B(n780), .Z(n784) );
  NAND2_X1 U868 ( .A1(n872), .A2(G131), .ZN(n782) );
  NAND2_X1 U869 ( .A1(G95), .A2(n880), .ZN(n781) );
  AND2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n858) );
  AND2_X1 U872 ( .A1(n858), .A2(G1991), .ZN(n795) );
  NAND2_X1 U873 ( .A1(G117), .A2(n874), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G129), .A2(n875), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n791) );
  XOR2_X1 U876 ( .A(KEYINPUT38), .B(KEYINPUT90), .Z(n788) );
  NAND2_X1 U877 ( .A1(G105), .A2(n880), .ZN(n787) );
  XNOR2_X1 U878 ( .A(n788), .B(n787), .ZN(n789) );
  XOR2_X1 U879 ( .A(KEYINPUT89), .B(n789), .Z(n790) );
  NOR2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n793) );
  NAND2_X1 U881 ( .A1(G141), .A2(n872), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n852) );
  AND2_X1 U883 ( .A1(n852), .A2(G1996), .ZN(n794) );
  NOR2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n926) );
  XNOR2_X1 U885 ( .A(KEYINPUT91), .B(n810), .ZN(n796) );
  NOR2_X1 U886 ( .A1(n926), .A2(n796), .ZN(n804) );
  INV_X1 U887 ( .A(n804), .ZN(n797) );
  NAND2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U889 ( .A(n799), .B(KEYINPUT99), .ZN(n801) );
  XNOR2_X1 U890 ( .A(G1986), .B(G290), .ZN(n957) );
  NAND2_X1 U891 ( .A1(n957), .A2(n810), .ZN(n800) );
  NAND2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n813) );
  NOR2_X1 U893 ( .A1(G1996), .A2(n852), .ZN(n915) );
  NOR2_X1 U894 ( .A1(G1986), .A2(G290), .ZN(n802) );
  NOR2_X1 U895 ( .A1(G1991), .A2(n858), .ZN(n919) );
  NOR2_X1 U896 ( .A1(n802), .A2(n919), .ZN(n803) );
  NOR2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U898 ( .A1(n915), .A2(n805), .ZN(n806) );
  XNOR2_X1 U899 ( .A(n806), .B(KEYINPUT39), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n807), .A2(n524), .ZN(n809) );
  NAND2_X1 U901 ( .A1(n808), .A2(n887), .ZN(n934) );
  NAND2_X1 U902 ( .A1(n809), .A2(n934), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U904 ( .A1(n813), .A2(n812), .ZN(n816) );
  XOR2_X1 U905 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n814) );
  XNOR2_X1 U906 ( .A(KEYINPUT40), .B(n814), .ZN(n815) );
  XNOR2_X1 U907 ( .A(n816), .B(n815), .ZN(G329) );
  NAND2_X1 U908 ( .A1(G2106), .A2(n817), .ZN(G217) );
  INV_X1 U909 ( .A(n817), .ZN(G223) );
  AND2_X1 U910 ( .A1(G15), .A2(G2), .ZN(n818) );
  NAND2_X1 U911 ( .A1(G661), .A2(n818), .ZN(G259) );
  NAND2_X1 U912 ( .A1(G3), .A2(G1), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n820), .A2(n819), .ZN(G188) );
  INV_X1 U915 ( .A(G132), .ZN(G219) );
  INV_X1 U916 ( .A(G120), .ZN(G236) );
  INV_X1 U917 ( .A(G96), .ZN(G221) );
  INV_X1 U918 ( .A(G82), .ZN(G220) );
  INV_X1 U919 ( .A(G69), .ZN(G235) );
  NOR2_X1 U920 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U921 ( .A(n823), .B(KEYINPUT103), .Z(G325) );
  INV_X1 U922 ( .A(G325), .ZN(G261) );
  XOR2_X1 U923 ( .A(n824), .B(KEYINPUT41), .Z(n834) );
  XNOR2_X1 U924 ( .A(G1976), .B(n951), .ZN(n826) );
  XNOR2_X1 U925 ( .A(G1991), .B(G1961), .ZN(n825) );
  XNOR2_X1 U926 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U927 ( .A(G1981), .B(G1971), .Z(n828) );
  XNOR2_X1 U928 ( .A(G1986), .B(G1966), .ZN(n827) );
  XNOR2_X1 U929 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U930 ( .A(n830), .B(n829), .Z(n832) );
  XNOR2_X1 U931 ( .A(KEYINPUT104), .B(G2474), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(G229) );
  XNOR2_X1 U934 ( .A(n835), .B(G2096), .ZN(n837) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(G2678), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U937 ( .A(KEYINPUT43), .B(G2090), .Z(n839) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U940 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2084), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(G227) );
  INV_X1 U943 ( .A(n844), .ZN(G319) );
  NAND2_X1 U944 ( .A1(G124), .A2(n875), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n845), .B(KEYINPUT44), .ZN(n847) );
  NAND2_X1 U946 ( .A1(n880), .A2(G100), .ZN(n846) );
  NAND2_X1 U947 ( .A1(n847), .A2(n846), .ZN(n851) );
  NAND2_X1 U948 ( .A1(n874), .A2(G112), .ZN(n849) );
  NAND2_X1 U949 ( .A1(G136), .A2(n872), .ZN(n848) );
  NAND2_X1 U950 ( .A1(n849), .A2(n848), .ZN(n850) );
  NOR2_X1 U951 ( .A1(n851), .A2(n850), .ZN(G162) );
  XOR2_X1 U952 ( .A(KEYINPUT46), .B(KEYINPUT107), .Z(n854) );
  XOR2_X1 U953 ( .A(n852), .B(KEYINPUT48), .Z(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U955 ( .A(n855), .B(KEYINPUT108), .Z(n857) );
  XNOR2_X1 U956 ( .A(G164), .B(KEYINPUT111), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n862) );
  XOR2_X1 U958 ( .A(n918), .B(G162), .Z(n860) );
  XOR2_X1 U959 ( .A(G160), .B(n858), .Z(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n889) );
  NAND2_X1 U962 ( .A1(G130), .A2(n875), .ZN(n871) );
  NAND2_X1 U963 ( .A1(n874), .A2(G118), .ZN(n863) );
  XNOR2_X1 U964 ( .A(KEYINPUT105), .B(n863), .ZN(n869) );
  NAND2_X1 U965 ( .A1(G106), .A2(n880), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G142), .A2(n872), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U968 ( .A(KEYINPUT45), .B(n866), .Z(n867) );
  XNOR2_X1 U969 ( .A(KEYINPUT106), .B(n867), .ZN(n868) );
  NOR2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n885) );
  NAND2_X1 U972 ( .A1(G139), .A2(n872), .ZN(n873) );
  XNOR2_X1 U973 ( .A(KEYINPUT109), .B(n873), .ZN(n884) );
  NAND2_X1 U974 ( .A1(G115), .A2(n874), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G127), .A2(n875), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n878), .B(KEYINPUT110), .ZN(n879) );
  XNOR2_X1 U978 ( .A(n879), .B(KEYINPUT47), .ZN(n882) );
  NAND2_X1 U979 ( .A1(n880), .A2(G103), .ZN(n881) );
  NAND2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n927) );
  XNOR2_X1 U982 ( .A(n885), .B(n927), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U984 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U985 ( .A1(G37), .A2(n890), .ZN(G395) );
  XOR2_X1 U986 ( .A(n686), .B(G286), .Z(n893) );
  XOR2_X1 U987 ( .A(G301), .B(n891), .Z(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n895) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U990 ( .A1(G37), .A2(n896), .ZN(G397) );
  XNOR2_X1 U991 ( .A(KEYINPUT49), .B(KEYINPUT112), .ZN(n898) );
  NOR2_X1 U992 ( .A1(G229), .A2(G227), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n910) );
  XOR2_X1 U994 ( .A(KEYINPUT102), .B(G2446), .Z(n900) );
  XNOR2_X1 U995 ( .A(G2443), .B(G2454), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U997 ( .A(n901), .B(G2451), .Z(n903) );
  XNOR2_X1 U998 ( .A(G1348), .B(G1341), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U1000 ( .A(G2435), .B(G2427), .Z(n905) );
  XNOR2_X1 U1001 ( .A(G2430), .B(G2438), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1003 ( .A(n907), .B(n906), .Z(n908) );
  NAND2_X1 U1004 ( .A1(G14), .A2(n908), .ZN(n913) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n913), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(G108), .ZN(G238) );
  INV_X1 U1011 ( .A(n913), .ZN(G401) );
  XOR2_X1 U1012 ( .A(G2090), .B(G162), .Z(n914) );
  NOR2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1014 ( .A(KEYINPUT51), .B(n916), .Z(n917) );
  XNOR2_X1 U1015 ( .A(KEYINPUT114), .B(n917), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n924) );
  XNOR2_X1 U1018 ( .A(G2084), .B(G160), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(KEYINPUT113), .B(n922), .ZN(n923) );
  NOR2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n933) );
  XNOR2_X1 U1022 ( .A(G2072), .B(n927), .ZN(n929) );
  XNOR2_X1 U1023 ( .A(G164), .B(G2078), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1025 ( .A(KEYINPUT50), .B(n930), .Z(n931) );
  XNOR2_X1 U1026 ( .A(KEYINPUT115), .B(n931), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n935) );
  NAND2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1029 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1030 ( .A(KEYINPUT52), .B(n938), .ZN(n939) );
  INV_X1 U1031 ( .A(KEYINPUT55), .ZN(n1016) );
  NAND2_X1 U1032 ( .A1(n939), .A2(n1016), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(n940), .A2(G29), .ZN(n1025) );
  XOR2_X1 U1034 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n941) );
  XOR2_X1 U1035 ( .A(G16), .B(n941), .Z(n970) );
  XNOR2_X1 U1036 ( .A(G1966), .B(G168), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(n944), .B(KEYINPUT57), .ZN(n945) );
  XOR2_X1 U1039 ( .A(KEYINPUT121), .B(n945), .Z(n968) );
  XOR2_X1 U1040 ( .A(G301), .B(G1961), .Z(n949) );
  XOR2_X1 U1041 ( .A(G1348), .B(n946), .Z(n947) );
  XNOR2_X1 U1042 ( .A(n947), .B(KEYINPUT122), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(n950), .B(KEYINPUT123), .ZN(n964) );
  XOR2_X1 U1045 ( .A(n952), .B(n951), .Z(n959) );
  INV_X1 U1046 ( .A(n953), .ZN(n955) );
  NAND2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1048 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1049 ( .A1(n959), .A2(n958), .ZN(n962) );
  XNOR2_X1 U1050 ( .A(G1971), .B(G303), .ZN(n960) );
  XNOR2_X1 U1051 ( .A(KEYINPUT124), .B(n960), .ZN(n961) );
  NOR2_X1 U1052 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1053 ( .A1(n964), .A2(n963), .ZN(n966) );
  XOR2_X1 U1054 ( .A(G1341), .B(n686), .Z(n965) );
  NOR2_X1 U1055 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1056 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1057 ( .A1(n970), .A2(n969), .ZN(n997) );
  INV_X1 U1058 ( .A(G16), .ZN(n995) );
  XOR2_X1 U1059 ( .A(G1971), .B(G22), .Z(n973) );
  XOR2_X1 U1060 ( .A(G24), .B(KEYINPUT126), .Z(n971) );
  XNOR2_X1 U1061 ( .A(n971), .B(G1986), .ZN(n972) );
  NAND2_X1 U1062 ( .A1(n973), .A2(n972), .ZN(n975) );
  XNOR2_X1 U1063 ( .A(G23), .B(G1976), .ZN(n974) );
  NOR2_X1 U1064 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1065 ( .A(KEYINPUT58), .B(n976), .Z(n992) );
  XOR2_X1 U1066 ( .A(G20), .B(G1956), .Z(n980) );
  XNOR2_X1 U1067 ( .A(G1341), .B(G19), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(G1981), .B(G6), .ZN(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n983) );
  XOR2_X1 U1071 ( .A(KEYINPUT59), .B(G1348), .Z(n981) );
  XNOR2_X1 U1072 ( .A(G4), .B(n981), .ZN(n982) );
  NOR2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(KEYINPUT60), .B(n984), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(n985), .B(G5), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n989) );
  XNOR2_X1 U1077 ( .A(G21), .B(G1966), .ZN(n988) );
  NOR2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(KEYINPUT125), .B(n990), .ZN(n991) );
  NOR2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(KEYINPUT61), .B(n993), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n1023) );
  XOR2_X1 U1084 ( .A(G29), .B(KEYINPUT118), .Z(n1019) );
  XOR2_X1 U1085 ( .A(G2090), .B(G35), .Z(n1012) );
  XNOR2_X1 U1086 ( .A(G27), .B(n998), .ZN(n1004) );
  XOR2_X1 U1087 ( .A(G32), .B(G1996), .Z(n999) );
  NAND2_X1 U1088 ( .A1(n999), .A2(G28), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(KEYINPUT116), .B(G2072), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(G33), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1008) );
  XOR2_X1 U1093 ( .A(G2067), .B(G26), .Z(n1006) );
  XOR2_X1 U1094 ( .A(G1991), .B(G25), .Z(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(n1009), .B(KEYINPUT117), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(n1010), .B(KEYINPUT53), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XNOR2_X1 U1100 ( .A(G34), .B(G2084), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT54), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XOR2_X1 U1103 ( .A(n1017), .B(n1016), .Z(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(G11), .ZN(n1021) );
  XOR2_X1 U1106 ( .A(KEYINPUT119), .B(n1021), .Z(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1109 ( .A(n1026), .B(KEYINPUT127), .ZN(n1027) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1027), .Z(G150) );
  INV_X1 U1111 ( .A(G150), .ZN(G311) );
endmodule

