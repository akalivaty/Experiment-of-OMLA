

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X2 U555 ( .A(n892), .Z(n521) );
  XOR2_X1 U556 ( .A(KEYINPUT17), .B(n532), .Z(n892) );
  INV_X1 U557 ( .A(n680), .ZN(n697) );
  XOR2_X1 U558 ( .A(n680), .B(KEYINPUT93), .Z(n677) );
  NOR2_X1 U559 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  NOR2_X2 U560 ( .A1(n542), .A2(n541), .ZN(G164) );
  NOR2_X1 U561 ( .A1(n551), .A2(n550), .ZN(G160) );
  XOR2_X1 U562 ( .A(KEYINPUT29), .B(n676), .Z(n522) );
  XNOR2_X1 U563 ( .A(KEYINPUT104), .B(n757), .ZN(n523) );
  INV_X1 U564 ( .A(KEYINPUT28), .ZN(n640) );
  XNOR2_X1 U565 ( .A(n689), .B(KEYINPUT30), .ZN(n690) );
  XNOR2_X1 U566 ( .A(n687), .B(KEYINPUT92), .ZN(n735) );
  NOR2_X1 U567 ( .A1(G651), .A2(n584), .ZN(n787) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n790) );
  NAND2_X1 U569 ( .A1(n758), .A2(n523), .ZN(n759) );
  NAND2_X1 U570 ( .A1(G85), .A2(n790), .ZN(n525) );
  XOR2_X1 U571 ( .A(G543), .B(KEYINPUT0), .Z(n584) );
  INV_X1 U572 ( .A(G651), .ZN(n526) );
  NOR2_X1 U573 ( .A1(n584), .A2(n526), .ZN(n791) );
  NAND2_X1 U574 ( .A1(G72), .A2(n791), .ZN(n524) );
  NAND2_X1 U575 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X1 U576 ( .A1(G543), .A2(n526), .ZN(n527) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n527), .Z(n786) );
  NAND2_X1 U578 ( .A1(G60), .A2(n786), .ZN(n529) );
  NAND2_X1 U579 ( .A1(G47), .A2(n787), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n530) );
  OR2_X1 U581 ( .A1(n531), .A2(n530), .ZN(G290) );
  NAND2_X1 U582 ( .A1(n521), .A2(G138), .ZN(n534) );
  INV_X1 U583 ( .A(KEYINPUT87), .ZN(n533) );
  XNOR2_X1 U584 ( .A(n534), .B(n533), .ZN(n537) );
  NAND2_X1 U585 ( .A1(G2104), .A2(G2105), .ZN(n535) );
  XNOR2_X1 U586 ( .A(n535), .B(KEYINPUT67), .ZN(n886) );
  NAND2_X1 U587 ( .A1(n886), .A2(G114), .ZN(n536) );
  NAND2_X1 U588 ( .A1(n537), .A2(n536), .ZN(n542) );
  INV_X1 U589 ( .A(G2105), .ZN(n538) );
  AND2_X1 U590 ( .A1(n538), .A2(G2104), .ZN(n890) );
  NAND2_X1 U591 ( .A1(G102), .A2(n890), .ZN(n540) );
  NOR2_X2 U592 ( .A1(G2104), .A2(n538), .ZN(n887) );
  NAND2_X1 U593 ( .A1(G126), .A2(n887), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U595 ( .A1(G137), .A2(n521), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G113), .A2(n886), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n551) );
  NAND2_X1 U598 ( .A1(n887), .A2(G125), .ZN(n545) );
  XNOR2_X1 U599 ( .A(KEYINPUT65), .B(n545), .ZN(n548) );
  NAND2_X1 U600 ( .A1(n890), .A2(G101), .ZN(n546) );
  XNOR2_X1 U601 ( .A(KEYINPUT23), .B(n546), .ZN(n547) );
  NOR2_X1 U602 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U603 ( .A(KEYINPUT66), .B(n549), .Z(n550) );
  NAND2_X1 U604 ( .A1(G64), .A2(n786), .ZN(n553) );
  NAND2_X1 U605 ( .A1(G52), .A2(n787), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U607 ( .A(KEYINPUT68), .B(n554), .ZN(n559) );
  NAND2_X1 U608 ( .A1(G90), .A2(n790), .ZN(n556) );
  NAND2_X1 U609 ( .A1(G77), .A2(n791), .ZN(n555) );
  NAND2_X1 U610 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U611 ( .A(KEYINPUT9), .B(n557), .Z(n558) );
  NOR2_X1 U612 ( .A1(n559), .A2(n558), .ZN(G171) );
  NAND2_X1 U613 ( .A1(G76), .A2(n791), .ZN(n563) );
  XOR2_X1 U614 ( .A(KEYINPUT4), .B(KEYINPUT71), .Z(n561) );
  NAND2_X1 U615 ( .A1(G89), .A2(n790), .ZN(n560) );
  XNOR2_X1 U616 ( .A(n561), .B(n560), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U618 ( .A(n564), .B(KEYINPUT5), .ZN(n565) );
  XNOR2_X1 U619 ( .A(n565), .B(KEYINPUT72), .ZN(n571) );
  NAND2_X1 U620 ( .A1(n786), .A2(G63), .ZN(n566) );
  XOR2_X1 U621 ( .A(KEYINPUT73), .B(n566), .Z(n568) );
  NAND2_X1 U622 ( .A1(n787), .A2(G51), .ZN(n567) );
  NAND2_X1 U623 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U624 ( .A(KEYINPUT6), .B(n569), .Z(n570) );
  NAND2_X1 U625 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U626 ( .A(n572), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G62), .A2(n786), .ZN(n574) );
  NAND2_X1 U629 ( .A1(G50), .A2(n787), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U631 ( .A(KEYINPUT80), .B(n575), .ZN(n578) );
  NAND2_X1 U632 ( .A1(G75), .A2(n791), .ZN(n576) );
  XNOR2_X1 U633 ( .A(KEYINPUT81), .B(n576), .ZN(n577) );
  NOR2_X1 U634 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U635 ( .A1(n790), .A2(G88), .ZN(n579) );
  NAND2_X1 U636 ( .A1(n580), .A2(n579), .ZN(G303) );
  NAND2_X1 U637 ( .A1(G49), .A2(n787), .ZN(n582) );
  NAND2_X1 U638 ( .A1(G74), .A2(G651), .ZN(n581) );
  NAND2_X1 U639 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U640 ( .A1(n786), .A2(n583), .ZN(n586) );
  NAND2_X1 U641 ( .A1(n584), .A2(G87), .ZN(n585) );
  NAND2_X1 U642 ( .A1(n586), .A2(n585), .ZN(G288) );
  XOR2_X1 U643 ( .A(KEYINPUT2), .B(KEYINPUT78), .Z(n588) );
  NAND2_X1 U644 ( .A1(G73), .A2(n791), .ZN(n587) );
  XNOR2_X1 U645 ( .A(n588), .B(n587), .ZN(n592) );
  NAND2_X1 U646 ( .A1(n786), .A2(G61), .ZN(n590) );
  NAND2_X1 U647 ( .A1(n790), .A2(G86), .ZN(n589) );
  NAND2_X1 U648 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U649 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U650 ( .A(KEYINPUT79), .B(n593), .Z(n595) );
  NAND2_X1 U651 ( .A1(n787), .A2(G48), .ZN(n594) );
  NAND2_X1 U652 ( .A1(n595), .A2(n594), .ZN(G305) );
  XOR2_X1 U653 ( .A(KEYINPUT88), .B(G1986), .Z(n596) );
  XNOR2_X1 U654 ( .A(G290), .B(n596), .ZN(n981) );
  NAND2_X1 U655 ( .A1(G131), .A2(n521), .ZN(n598) );
  NAND2_X1 U656 ( .A1(G95), .A2(n890), .ZN(n597) );
  NAND2_X1 U657 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U658 ( .A1(G107), .A2(n886), .ZN(n600) );
  NAND2_X1 U659 ( .A1(G119), .A2(n887), .ZN(n599) );
  NAND2_X1 U660 ( .A1(n600), .A2(n599), .ZN(n601) );
  OR2_X1 U661 ( .A1(n602), .A2(n601), .ZN(n878) );
  XOR2_X1 U662 ( .A(KEYINPUT89), .B(G1991), .Z(n956) );
  AND2_X1 U663 ( .A1(n878), .A2(n956), .ZN(n603) );
  XNOR2_X1 U664 ( .A(n603), .B(KEYINPUT90), .ZN(n613) );
  NAND2_X1 U665 ( .A1(G141), .A2(n521), .ZN(n605) );
  NAND2_X1 U666 ( .A1(G129), .A2(n887), .ZN(n604) );
  NAND2_X1 U667 ( .A1(n605), .A2(n604), .ZN(n611) );
  NAND2_X1 U668 ( .A1(G105), .A2(n890), .ZN(n606) );
  XNOR2_X1 U669 ( .A(n606), .B(KEYINPUT38), .ZN(n609) );
  NAND2_X1 U670 ( .A1(G117), .A2(n886), .ZN(n607) );
  XOR2_X1 U671 ( .A(KEYINPUT91), .B(n607), .Z(n608) );
  NAND2_X1 U672 ( .A1(n609), .A2(n608), .ZN(n610) );
  OR2_X1 U673 ( .A1(n611), .A2(n610), .ZN(n879) );
  AND2_X1 U674 ( .A1(G1996), .A2(n879), .ZN(n612) );
  NOR2_X1 U675 ( .A1(n613), .A2(n612), .ZN(n927) );
  NAND2_X1 U676 ( .A1(n981), .A2(n927), .ZN(n617) );
  NOR2_X1 U677 ( .A1(G1384), .A2(G164), .ZN(n615) );
  INV_X1 U678 ( .A(KEYINPUT64), .ZN(n614) );
  XNOR2_X1 U679 ( .A(n615), .B(n614), .ZN(n634) );
  INV_X1 U680 ( .A(n634), .ZN(n616) );
  NAND2_X1 U681 ( .A1(G160), .A2(G40), .ZN(n635) );
  NOR2_X1 U682 ( .A1(n616), .A2(n635), .ZN(n756) );
  NAND2_X1 U683 ( .A1(n617), .A2(n756), .ZN(n627) );
  NAND2_X1 U684 ( .A1(G140), .A2(n521), .ZN(n619) );
  NAND2_X1 U685 ( .A1(G104), .A2(n890), .ZN(n618) );
  NAND2_X1 U686 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U687 ( .A(KEYINPUT34), .B(n620), .ZN(n625) );
  NAND2_X1 U688 ( .A1(G116), .A2(n886), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G128), .A2(n887), .ZN(n621) );
  NAND2_X1 U690 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U691 ( .A(KEYINPUT35), .B(n623), .Z(n624) );
  NOR2_X1 U692 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U693 ( .A(KEYINPUT36), .B(n626), .ZN(n880) );
  XNOR2_X1 U694 ( .A(G2067), .B(KEYINPUT37), .ZN(n753) );
  NOR2_X1 U695 ( .A1(n880), .A2(n753), .ZN(n931) );
  NAND2_X1 U696 ( .A1(n931), .A2(n756), .ZN(n751) );
  NAND2_X1 U697 ( .A1(n627), .A2(n751), .ZN(n742) );
  NAND2_X1 U698 ( .A1(G65), .A2(n786), .ZN(n629) );
  NAND2_X1 U699 ( .A1(G53), .A2(n787), .ZN(n628) );
  NAND2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U701 ( .A1(G91), .A2(n790), .ZN(n631) );
  NAND2_X1 U702 ( .A1(G78), .A2(n791), .ZN(n630) );
  NAND2_X1 U703 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U704 ( .A1(n633), .A2(n632), .ZN(n988) );
  XOR2_X1 U705 ( .A(KEYINPUT97), .B(KEYINPUT27), .Z(n637) );
  NOR2_X2 U706 ( .A1(n635), .A2(n634), .ZN(n680) );
  NAND2_X1 U707 ( .A1(G2072), .A2(n677), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n637), .B(n636), .ZN(n639) );
  INV_X1 U709 ( .A(G1956), .ZN(n1006) );
  NOR2_X1 U710 ( .A1(n677), .A2(n1006), .ZN(n638) );
  NOR2_X1 U711 ( .A1(n639), .A2(n638), .ZN(n642) );
  NOR2_X1 U712 ( .A1(n988), .A2(n642), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n641), .B(n640), .ZN(n675) );
  NAND2_X1 U714 ( .A1(n988), .A2(n642), .ZN(n673) );
  NAND2_X1 U715 ( .A1(n680), .A2(G1996), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n643), .B(KEYINPUT26), .ZN(n645) );
  NAND2_X1 U717 ( .A1(G1341), .A2(n697), .ZN(n644) );
  NAND2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U719 ( .A(KEYINPUT98), .B(n646), .Z(n666) );
  NAND2_X1 U720 ( .A1(n790), .A2(G81), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n647), .B(KEYINPUT12), .ZN(n649) );
  NAND2_X1 U722 ( .A1(G68), .A2(n791), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U724 ( .A(n650), .B(KEYINPUT13), .ZN(n652) );
  NAND2_X1 U725 ( .A1(G43), .A2(n787), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U727 ( .A1(n786), .A2(G56), .ZN(n653) );
  XOR2_X1 U728 ( .A(KEYINPUT14), .B(n653), .Z(n654) );
  NOR2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n980) );
  NAND2_X1 U730 ( .A1(n666), .A2(n980), .ZN(n663) );
  NAND2_X1 U731 ( .A1(G66), .A2(n786), .ZN(n657) );
  NAND2_X1 U732 ( .A1(G54), .A2(n787), .ZN(n656) );
  NAND2_X1 U733 ( .A1(n657), .A2(n656), .ZN(n661) );
  NAND2_X1 U734 ( .A1(G92), .A2(n790), .ZN(n659) );
  NAND2_X1 U735 ( .A1(G79), .A2(n791), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U737 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U738 ( .A(n662), .B(KEYINPUT15), .ZN(n987) );
  NAND2_X1 U739 ( .A1(n663), .A2(n987), .ZN(n671) );
  NAND2_X1 U740 ( .A1(n697), .A2(G1348), .ZN(n665) );
  NAND2_X1 U741 ( .A1(G2067), .A2(n677), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n665), .A2(n664), .ZN(n669) );
  INV_X1 U743 ( .A(n980), .ZN(n772) );
  NOR2_X1 U744 ( .A1(n772), .A2(n987), .ZN(n667) );
  NAND2_X1 U745 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U746 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U747 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U748 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U749 ( .A1(n675), .A2(n674), .ZN(n676) );
  INV_X1 U750 ( .A(n677), .ZN(n679) );
  XOR2_X1 U751 ( .A(G2078), .B(KEYINPUT25), .Z(n678) );
  XNOR2_X1 U752 ( .A(KEYINPUT94), .B(n678), .ZN(n955) );
  NOR2_X1 U753 ( .A1(n679), .A2(n955), .ZN(n682) );
  NOR2_X1 U754 ( .A1(n680), .A2(G1961), .ZN(n681) );
  NOR2_X1 U755 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U756 ( .A(KEYINPUT95), .B(n683), .ZN(n686) );
  NAND2_X1 U757 ( .A1(G171), .A2(n686), .ZN(n684) );
  XNOR2_X1 U758 ( .A(n684), .B(KEYINPUT96), .ZN(n685) );
  NAND2_X1 U759 ( .A1(n522), .A2(n685), .ZN(n695) );
  NOR2_X1 U760 ( .A1(G171), .A2(n686), .ZN(n692) );
  NAND2_X1 U761 ( .A1(G8), .A2(n697), .ZN(n687) );
  NOR2_X1 U762 ( .A1(n735), .A2(G1966), .ZN(n709) );
  NOR2_X1 U763 ( .A1(G2084), .A2(n697), .ZN(n707) );
  NOR2_X1 U764 ( .A1(n709), .A2(n707), .ZN(n688) );
  NAND2_X1 U765 ( .A1(G8), .A2(n688), .ZN(n689) );
  NOR2_X1 U766 ( .A1(n690), .A2(G168), .ZN(n691) );
  NOR2_X1 U767 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U768 ( .A(KEYINPUT31), .B(n693), .Z(n694) );
  NAND2_X1 U769 ( .A1(n695), .A2(n694), .ZN(n711) );
  AND2_X1 U770 ( .A1(G286), .A2(G8), .ZN(n696) );
  NAND2_X1 U771 ( .A1(n711), .A2(n696), .ZN(n705) );
  INV_X1 U772 ( .A(G8), .ZN(n703) );
  NOR2_X1 U773 ( .A1(G2090), .A2(n697), .ZN(n698) );
  XNOR2_X1 U774 ( .A(n698), .B(KEYINPUT100), .ZN(n700) );
  NOR2_X1 U775 ( .A1(n735), .A2(G1971), .ZN(n699) );
  NOR2_X1 U776 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U777 ( .A1(n701), .A2(G303), .ZN(n702) );
  OR2_X1 U778 ( .A1(n703), .A2(n702), .ZN(n704) );
  AND2_X1 U779 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U780 ( .A(n706), .B(KEYINPUT32), .ZN(n714) );
  AND2_X1 U781 ( .A1(G8), .A2(n707), .ZN(n708) );
  NOR2_X1 U782 ( .A1(n709), .A2(n708), .ZN(n710) );
  AND2_X1 U783 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U784 ( .A(n712), .B(KEYINPUT99), .ZN(n713) );
  NAND2_X1 U785 ( .A1(n714), .A2(n713), .ZN(n734) );
  NOR2_X1 U786 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NOR2_X1 U787 ( .A1(G1971), .A2(G303), .ZN(n715) );
  NOR2_X1 U788 ( .A1(n974), .A2(n715), .ZN(n717) );
  INV_X1 U789 ( .A(KEYINPUT33), .ZN(n716) );
  AND2_X1 U790 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U791 ( .A1(n734), .A2(n718), .ZN(n727) );
  NAND2_X1 U792 ( .A1(n974), .A2(KEYINPUT33), .ZN(n719) );
  NOR2_X1 U793 ( .A1(n735), .A2(n719), .ZN(n721) );
  XOR2_X1 U794 ( .A(G1981), .B(G305), .Z(n983) );
  INV_X1 U795 ( .A(n983), .ZN(n720) );
  NOR2_X1 U796 ( .A1(n721), .A2(n720), .ZN(n725) );
  NAND2_X1 U797 ( .A1(G1976), .A2(G288), .ZN(n976) );
  INV_X1 U798 ( .A(n976), .ZN(n722) );
  NOR2_X1 U799 ( .A1(n735), .A2(n722), .ZN(n723) );
  OR2_X1 U800 ( .A1(KEYINPUT33), .A2(n723), .ZN(n724) );
  AND2_X1 U801 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U802 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U803 ( .A(n728), .B(KEYINPUT101), .ZN(n740) );
  NOR2_X1 U804 ( .A1(G1981), .A2(G305), .ZN(n729) );
  XNOR2_X1 U805 ( .A(KEYINPUT24), .B(n729), .ZN(n731) );
  INV_X1 U806 ( .A(n735), .ZN(n730) );
  NAND2_X1 U807 ( .A1(n731), .A2(n730), .ZN(n738) );
  NOR2_X1 U808 ( .A1(G2090), .A2(G303), .ZN(n732) );
  NAND2_X1 U809 ( .A1(G8), .A2(n732), .ZN(n733) );
  NAND2_X1 U810 ( .A1(n734), .A2(n733), .ZN(n736) );
  NAND2_X1 U811 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U813 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U814 ( .A1(n742), .A2(n741), .ZN(n743) );
  INV_X1 U815 ( .A(n743), .ZN(n758) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n879), .ZN(n940) );
  NOR2_X1 U817 ( .A1(n956), .A2(n878), .ZN(n930) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n744) );
  XNOR2_X1 U819 ( .A(KEYINPUT102), .B(n744), .ZN(n745) );
  NOR2_X1 U820 ( .A1(n930), .A2(n745), .ZN(n747) );
  INV_X1 U821 ( .A(n927), .ZN(n746) );
  NOR2_X1 U822 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U823 ( .A(KEYINPUT103), .B(n748), .Z(n749) );
  NOR2_X1 U824 ( .A1(n940), .A2(n749), .ZN(n750) );
  XNOR2_X1 U825 ( .A(n750), .B(KEYINPUT39), .ZN(n752) );
  NAND2_X1 U826 ( .A1(n752), .A2(n751), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n880), .A2(n753), .ZN(n926) );
  NAND2_X1 U828 ( .A1(n754), .A2(n926), .ZN(n755) );
  NAND2_X1 U829 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U830 ( .A(n759), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U831 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U832 ( .A(G57), .ZN(G237) );
  INV_X1 U833 ( .A(G69), .ZN(G235) );
  INV_X1 U834 ( .A(G108), .ZN(G238) );
  INV_X1 U835 ( .A(G120), .ZN(G236) );
  INV_X1 U836 ( .A(G132), .ZN(G219) );
  INV_X1 U837 ( .A(G82), .ZN(G220) );
  XOR2_X1 U838 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n761) );
  NAND2_X1 U839 ( .A1(G7), .A2(G661), .ZN(n760) );
  XNOR2_X1 U840 ( .A(n761), .B(n760), .ZN(G223) );
  XOR2_X1 U841 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n763) );
  INV_X1 U842 ( .A(G223), .ZN(n829) );
  NAND2_X1 U843 ( .A1(G567), .A2(n829), .ZN(n762) );
  XNOR2_X1 U844 ( .A(n763), .B(n762), .ZN(G234) );
  NAND2_X1 U845 ( .A1(n980), .A2(G860), .ZN(G153) );
  INV_X1 U846 ( .A(G171), .ZN(G301) );
  NAND2_X1 U847 ( .A1(G868), .A2(G301), .ZN(n765) );
  INV_X1 U848 ( .A(G868), .ZN(n810) );
  NAND2_X1 U849 ( .A1(n987), .A2(n810), .ZN(n764) );
  NAND2_X1 U850 ( .A1(n765), .A2(n764), .ZN(G284) );
  INV_X1 U851 ( .A(n988), .ZN(G299) );
  XNOR2_X1 U852 ( .A(KEYINPUT74), .B(n810), .ZN(n766) );
  NOR2_X1 U853 ( .A1(G286), .A2(n766), .ZN(n768) );
  NOR2_X1 U854 ( .A1(G868), .A2(G299), .ZN(n767) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U856 ( .A(KEYINPUT75), .B(n769), .Z(G297) );
  INV_X1 U857 ( .A(G860), .ZN(n798) );
  NAND2_X1 U858 ( .A1(n798), .A2(G559), .ZN(n770) );
  INV_X1 U859 ( .A(n987), .ZN(n796) );
  NAND2_X1 U860 ( .A1(n770), .A2(n796), .ZN(n771) );
  XNOR2_X1 U861 ( .A(n771), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U862 ( .A1(G868), .A2(n772), .ZN(n775) );
  NAND2_X1 U863 ( .A1(G868), .A2(n796), .ZN(n773) );
  NOR2_X1 U864 ( .A1(G559), .A2(n773), .ZN(n774) );
  NOR2_X1 U865 ( .A1(n775), .A2(n774), .ZN(G282) );
  NAND2_X1 U866 ( .A1(G111), .A2(n886), .ZN(n777) );
  NAND2_X1 U867 ( .A1(G99), .A2(n890), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U869 ( .A(KEYINPUT76), .B(n778), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G123), .A2(n887), .ZN(n779) );
  XNOR2_X1 U871 ( .A(n779), .B(KEYINPUT18), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n521), .A2(G135), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U874 ( .A1(n783), .A2(n782), .ZN(n929) );
  XNOR2_X1 U875 ( .A(n929), .B(G2096), .ZN(n785) );
  INV_X1 U876 ( .A(G2100), .ZN(n784) );
  NAND2_X1 U877 ( .A1(n785), .A2(n784), .ZN(G156) );
  NAND2_X1 U878 ( .A1(G67), .A2(n786), .ZN(n789) );
  NAND2_X1 U879 ( .A1(G55), .A2(n787), .ZN(n788) );
  NAND2_X1 U880 ( .A1(n789), .A2(n788), .ZN(n795) );
  NAND2_X1 U881 ( .A1(G93), .A2(n790), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G80), .A2(n791), .ZN(n792) );
  NAND2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n809) );
  NAND2_X1 U885 ( .A1(G559), .A2(n796), .ZN(n797) );
  XNOR2_X1 U886 ( .A(n797), .B(n980), .ZN(n807) );
  NAND2_X1 U887 ( .A1(n798), .A2(n807), .ZN(n799) );
  XNOR2_X1 U888 ( .A(n799), .B(KEYINPUT77), .ZN(n800) );
  XNOR2_X1 U889 ( .A(n809), .B(n800), .ZN(G145) );
  INV_X1 U890 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U891 ( .A(n809), .B(KEYINPUT19), .ZN(n801) );
  XNOR2_X1 U892 ( .A(n801), .B(KEYINPUT82), .ZN(n802) );
  XNOR2_X1 U893 ( .A(n802), .B(G288), .ZN(n805) );
  XNOR2_X1 U894 ( .A(n988), .B(G166), .ZN(n803) );
  XNOR2_X1 U895 ( .A(n803), .B(G290), .ZN(n804) );
  XNOR2_X1 U896 ( .A(n805), .B(n804), .ZN(n806) );
  XNOR2_X1 U897 ( .A(n806), .B(G305), .ZN(n903) );
  XNOR2_X1 U898 ( .A(n807), .B(n903), .ZN(n808) );
  NAND2_X1 U899 ( .A1(n808), .A2(G868), .ZN(n812) );
  NAND2_X1 U900 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U901 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U902 ( .A(KEYINPUT83), .B(n813), .ZN(G295) );
  NAND2_X1 U903 ( .A1(G2078), .A2(G2084), .ZN(n814) );
  XOR2_X1 U904 ( .A(KEYINPUT20), .B(n814), .Z(n815) );
  NAND2_X1 U905 ( .A1(G2090), .A2(n815), .ZN(n817) );
  XNOR2_X1 U906 ( .A(KEYINPUT84), .B(KEYINPUT21), .ZN(n816) );
  XNOR2_X1 U907 ( .A(n817), .B(n816), .ZN(n818) );
  NAND2_X1 U908 ( .A1(G2072), .A2(n818), .ZN(G158) );
  XOR2_X1 U909 ( .A(KEYINPUT85), .B(G44), .Z(n819) );
  XNOR2_X1 U910 ( .A(KEYINPUT3), .B(n819), .ZN(G218) );
  NOR2_X1 U911 ( .A1(G220), .A2(G219), .ZN(n820) );
  XOR2_X1 U912 ( .A(KEYINPUT22), .B(n820), .Z(n821) );
  NOR2_X1 U913 ( .A1(G218), .A2(n821), .ZN(n822) );
  NAND2_X1 U914 ( .A1(G96), .A2(n822), .ZN(n835) );
  NAND2_X1 U915 ( .A1(n835), .A2(G2106), .ZN(n827) );
  NOR2_X1 U916 ( .A1(G236), .A2(G238), .ZN(n824) );
  NOR2_X1 U917 ( .A1(G235), .A2(G237), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U919 ( .A(KEYINPUT86), .B(n825), .ZN(n836) );
  NAND2_X1 U920 ( .A1(n836), .A2(G567), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n858) );
  NAND2_X1 U922 ( .A1(G661), .A2(G483), .ZN(n828) );
  NOR2_X1 U923 ( .A1(n858), .A2(n828), .ZN(n834) );
  NAND2_X1 U924 ( .A1(n834), .A2(G36), .ZN(G176) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n829), .ZN(G217) );
  NAND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n830) );
  XOR2_X1 U927 ( .A(KEYINPUT106), .B(n830), .Z(n831) );
  NAND2_X1 U928 ( .A1(n831), .A2(G661), .ZN(n832) );
  XOR2_X1 U929 ( .A(KEYINPUT107), .B(n832), .Z(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U931 ( .A1(n834), .A2(n833), .ZN(G188) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  NOR2_X1 U934 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XOR2_X1 U936 ( .A(KEYINPUT111), .B(G1991), .Z(n838) );
  XNOR2_X1 U937 ( .A(G1981), .B(G1996), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U939 ( .A(n839), .B(KEYINPUT41), .Z(n841) );
  XNOR2_X1 U940 ( .A(G1956), .B(G1976), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U942 ( .A(G1986), .B(G1971), .Z(n843) );
  XNOR2_X1 U943 ( .A(G1966), .B(G1961), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U945 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U946 ( .A(KEYINPUT110), .B(G2474), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(G229) );
  XOR2_X1 U948 ( .A(G2100), .B(KEYINPUT109), .Z(n849) );
  XNOR2_X1 U949 ( .A(G2678), .B(KEYINPUT108), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U951 ( .A(KEYINPUT43), .B(G2090), .Z(n851) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U954 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U955 ( .A(KEYINPUT42), .B(G2096), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n857) );
  XOR2_X1 U957 ( .A(G2078), .B(G2084), .Z(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(G227) );
  INV_X1 U959 ( .A(n858), .ZN(G319) );
  NAND2_X1 U960 ( .A1(G124), .A2(n887), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n886), .A2(G112), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n861), .A2(n860), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G136), .A2(n521), .ZN(n863) );
  NAND2_X1 U965 ( .A1(G100), .A2(n890), .ZN(n862) );
  NAND2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U967 ( .A1(n865), .A2(n864), .ZN(G162) );
  XOR2_X1 U968 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n876) );
  NAND2_X1 U969 ( .A1(G115), .A2(n886), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G127), .A2(n887), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U972 ( .A(n868), .B(KEYINPUT47), .ZN(n870) );
  NAND2_X1 U973 ( .A1(G103), .A2(n890), .ZN(n869) );
  NAND2_X1 U974 ( .A1(n870), .A2(n869), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G139), .A2(n521), .ZN(n871) );
  XNOR2_X1 U976 ( .A(KEYINPUT115), .B(n871), .ZN(n872) );
  NOR2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U978 ( .A(KEYINPUT116), .B(n874), .Z(n935) );
  XNOR2_X1 U979 ( .A(n935), .B(KEYINPUT114), .ZN(n875) );
  XNOR2_X1 U980 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U981 ( .A(n878), .B(n877), .Z(n882) );
  XOR2_X1 U982 ( .A(n880), .B(n879), .Z(n881) );
  XNOR2_X1 U983 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U984 ( .A(n883), .B(G162), .Z(n885) );
  XNOR2_X1 U985 ( .A(G164), .B(G160), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n901) );
  NAND2_X1 U987 ( .A1(G118), .A2(n886), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G130), .A2(n887), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n898) );
  NAND2_X1 U990 ( .A1(n890), .A2(G106), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n891), .B(KEYINPUT112), .ZN(n894) );
  NAND2_X1 U992 ( .A1(G142), .A2(n521), .ZN(n893) );
  NAND2_X1 U993 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U994 ( .A(KEYINPUT45), .B(n895), .ZN(n896) );
  XNOR2_X1 U995 ( .A(KEYINPUT113), .B(n896), .ZN(n897) );
  NOR2_X1 U996 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U997 ( .A(n929), .B(n899), .Z(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U999 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U1000 ( .A(KEYINPUT117), .B(n903), .Z(n905) );
  XNOR2_X1 U1001 ( .A(G171), .B(G286), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n907) );
  XOR2_X1 U1003 ( .A(n987), .B(n980), .Z(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n908), .ZN(G397) );
  NOR2_X1 U1006 ( .A1(G229), .A2(G227), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n922) );
  XOR2_X1 U1009 ( .A(G2454), .B(G2435), .Z(n912) );
  XNOR2_X1 U1010 ( .A(G2438), .B(G2427), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n912), .B(n911), .ZN(n919) );
  XOR2_X1 U1012 ( .A(KEYINPUT105), .B(G2446), .Z(n914) );
  XNOR2_X1 U1013 ( .A(G2443), .B(G2430), .ZN(n913) );
  XNOR2_X1 U1014 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1015 ( .A(n915), .B(G2451), .Z(n917) );
  XNOR2_X1 U1016 ( .A(G1348), .B(G1341), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n917), .B(n916), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n919), .B(n918), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n920), .A2(G14), .ZN(n925) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n925), .ZN(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(n925), .ZN(G401) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n947) );
  XOR2_X1 U1027 ( .A(G2084), .B(G160), .Z(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(KEYINPUT119), .B(n934), .ZN(n945) );
  XOR2_X1 U1032 ( .A(G164), .B(G2078), .Z(n937) );
  XNOR2_X1 U1033 ( .A(G2072), .B(n935), .ZN(n936) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1035 ( .A(KEYINPUT50), .B(n938), .Z(n943) );
  XOR2_X1 U1036 ( .A(G2090), .B(G162), .Z(n939) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(KEYINPUT51), .B(n941), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(KEYINPUT52), .B(n948), .ZN(n949) );
  XOR2_X1 U1043 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n970) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n970), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(n950), .A2(G29), .ZN(n1032) );
  XOR2_X1 U1046 ( .A(G2084), .B(G34), .Z(n951) );
  XNOR2_X1 U1047 ( .A(KEYINPUT54), .B(n951), .ZN(n967) );
  XNOR2_X1 U1048 ( .A(G2090), .B(G35), .ZN(n965) );
  XOR2_X1 U1049 ( .A(G2067), .B(G26), .Z(n952) );
  NAND2_X1 U1050 ( .A1(n952), .A2(G28), .ZN(n962) );
  XNOR2_X1 U1051 ( .A(G1996), .B(G32), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(n955), .B(G27), .ZN(n958) );
  XNOR2_X1 U1055 ( .A(G25), .B(n956), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(KEYINPUT53), .B(n963), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(n968), .B(KEYINPUT121), .ZN(n969) );
  XOR2_X1 U1063 ( .A(n970), .B(n969), .Z(n972) );
  INV_X1 U1064 ( .A(G29), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n973), .A2(G11), .ZN(n1030) );
  XNOR2_X1 U1067 ( .A(G16), .B(KEYINPUT56), .ZN(n1000) );
  INV_X1 U1068 ( .A(n974), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1070 ( .A(KEYINPUT123), .B(n977), .Z(n979) );
  XNOR2_X1 U1071 ( .A(G1961), .B(G301), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n998) );
  XNOR2_X1 U1073 ( .A(n980), .B(G1341), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n996) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G168), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(n985), .B(KEYINPUT122), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(KEYINPUT57), .B(n986), .ZN(n994) );
  XNOR2_X1 U1079 ( .A(G1348), .B(n987), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(G166), .B(G1971), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(n988), .B(G1956), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1028) );
  INV_X1 U1088 ( .A(G16), .ZN(n1026) );
  XOR2_X1 U1089 ( .A(G1341), .B(G19), .Z(n1005) );
  XOR2_X1 U1090 ( .A(KEYINPUT125), .B(G4), .Z(n1002) );
  XNOR2_X1 U1091 ( .A(G1348), .B(KEYINPUT59), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(n1002), .B(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(KEYINPUT124), .B(n1003), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1010) );
  XOR2_X1 U1095 ( .A(G1981), .B(G6), .Z(n1008) );
  XNOR2_X1 U1096 ( .A(n1006), .B(G20), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(KEYINPUT60), .B(n1011), .Z(n1013) );
  XNOR2_X1 U1100 ( .A(G1966), .B(G21), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT126), .B(n1014), .ZN(n1023) );
  XNOR2_X1 U1103 ( .A(G1961), .B(G5), .ZN(n1021) );
  XNOR2_X1 U1104 ( .A(G1971), .B(G22), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(G23), .B(G1976), .ZN(n1015) );
  NOR2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XOR2_X1 U1107 ( .A(G1986), .B(G24), .Z(n1017) );
  NAND2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1109 ( .A(KEYINPUT58), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1112 ( .A(KEYINPUT61), .B(n1024), .Z(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1117 ( .A(n1033), .B(KEYINPUT127), .ZN(n1034) );
  XNOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1034), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

