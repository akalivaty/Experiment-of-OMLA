//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n203), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  INV_X1    g0024(.A(G97), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n201), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(new_n224), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  AOI21_X1  g0045(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n246));
  INV_X1    g0046(.A(G274), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n248));
  NOR3_X1   g0048(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n248), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n249), .B1(G226), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G222), .A2(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G223), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n255), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n259), .B(new_n246), .C1(G77), .C2(new_n255), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G190), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n263), .B1(G200), .B2(new_n261), .ZN(new_n264));
  OAI21_X1  g0064(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n265));
  INV_X1    g0065(.A(G150), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT65), .B1(G20), .B2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NOR3_X1   g0068(.A1(KEYINPUT65), .A2(G20), .A3(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT8), .B(G58), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT64), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n201), .A2(KEYINPUT64), .A3(KEYINPUT8), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n207), .A2(G33), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n265), .B1(new_n266), .B2(new_n270), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n215), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G50), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n279), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(G1), .B2(new_n207), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n284), .B1(new_n286), .B2(new_n283), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(KEYINPUT9), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT9), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(new_n280), .B2(new_n288), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n264), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT10), .ZN(new_n294));
  INV_X1    g0094(.A(new_n289), .ZN(new_n295));
  INV_X1    g0095(.A(new_n261), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G169), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n298), .A2(KEYINPUT66), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n298), .A2(KEYINPUT66), .B1(new_n300), .B2(new_n296), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n294), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n224), .A2(G1698), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n255), .B(new_n304), .C1(G226), .C2(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G97), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n251), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(G1), .A2(G13), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n247), .B1(new_n309), .B2(new_n250), .ZN(new_n310));
  INV_X1    g0110(.A(new_n248), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n219), .B2(new_n252), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT13), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n308), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT13), .B1(new_n307), .B2(new_n313), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(KEYINPUT69), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT69), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n319), .B(KEYINPUT13), .C1(new_n307), .C2(new_n313), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(G169), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT14), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT14), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n318), .A2(new_n323), .A3(G169), .A4(new_n320), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n316), .A2(G179), .A3(new_n317), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n276), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n328));
  OAI21_X1  g0128(.A(G50), .B1(new_n268), .B2(new_n269), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n285), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n330), .A2(KEYINPUT11), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(KEYINPUT11), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n279), .B1(new_n206), .B2(G20), .ZN(new_n333));
  OR3_X1    g0133(.A1(new_n281), .A2(KEYINPUT12), .A3(G68), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT12), .B1(new_n281), .B2(G68), .ZN(new_n335));
  AOI22_X1  g0135(.A1(G68), .A2(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n331), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n326), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n316), .A2(G190), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n337), .B1(new_n339), .B2(new_n317), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n318), .A2(G200), .A3(new_n320), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT67), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT15), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G87), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(new_n327), .B1(G20), .B2(G77), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n270), .B2(new_n271), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n279), .ZN(new_n351));
  INV_X1    g0151(.A(G77), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n282), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n333), .A2(G77), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G200), .ZN(new_n356));
  INV_X1    g0156(.A(G244), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n312), .B1(new_n357), .B2(new_n252), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(G232), .A2(G1698), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n257), .A2(G238), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n255), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT3), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G33), .ZN(new_n364));
  INV_X1    g0164(.A(G33), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT3), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G107), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n362), .A2(new_n246), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n356), .B1(new_n359), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n344), .B1(new_n355), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n359), .A2(G190), .A3(new_n370), .ZN(new_n373));
  INV_X1    g0173(.A(new_n370), .ZN(new_n374));
  OAI21_X1  g0174(.A(G200), .B1(new_n374), .B2(new_n358), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n354), .A2(new_n353), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n375), .A2(KEYINPUT67), .A3(new_n351), .A4(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n372), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n359), .A2(new_n370), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT68), .B1(new_n379), .B2(G179), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT68), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n359), .A2(new_n381), .A3(new_n300), .A4(new_n370), .ZN(new_n382));
  INV_X1    g0182(.A(G169), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n380), .A2(new_n355), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  OR3_X1    g0187(.A1(new_n303), .A2(new_n343), .A3(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(G257), .A2(G1698), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n257), .A2(G264), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n255), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G303), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n367), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n246), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G41), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n206), .B(G45), .C1(new_n395), .C2(KEYINPUT5), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT77), .ZN(new_n397));
  INV_X1    g0197(.A(G45), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(G1), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT77), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT5), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G41), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n401), .A2(G41), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n397), .A2(new_n403), .A3(new_n405), .A4(new_n310), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT83), .ZN(new_n407));
  OAI211_X1 g0207(.A(G270), .B(new_n251), .C1(new_n396), .C2(new_n404), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n407), .B1(new_n406), .B2(new_n408), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n394), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G283), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n412), .B(new_n207), .C1(G33), .C2(new_n225), .ZN(new_n413));
  INV_X1    g0213(.A(G116), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G20), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n279), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT20), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n416), .B(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n206), .A2(G33), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n281), .A2(new_n419), .A3(new_n215), .A4(new_n278), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G116), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(G116), .B2(new_n282), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n383), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n411), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT21), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(G190), .B(new_n394), .C1(new_n409), .C2(new_n410), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n418), .A2(new_n422), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n394), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n406), .A2(new_n408), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT83), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n427), .B(new_n429), .C1(new_n434), .C2(new_n356), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(G179), .A3(new_n428), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n411), .A2(new_n423), .A3(KEYINPUT21), .ZN(new_n437));
  AND4_X1   g0237(.A1(new_n426), .A2(new_n435), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n364), .A2(new_n366), .A3(new_n207), .A4(G87), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT22), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT22), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n255), .A2(new_n441), .A3(new_n207), .A4(G87), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT85), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n207), .B2(G107), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT23), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT23), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n444), .B(new_n447), .C1(new_n207), .C2(G107), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n446), .A2(new_n448), .B1(G116), .B2(new_n327), .ZN(new_n449));
  XOR2_X1   g0249(.A(KEYINPUT84), .B(KEYINPUT24), .Z(new_n450));
  AND3_X1   g0250(.A1(new_n443), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n443), .B2(new_n449), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n279), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(G264), .B(new_n251), .C1(new_n396), .C2(new_n404), .ZN(new_n454));
  NOR2_X1   g0254(.A1(G250), .A2(G1698), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n226), .B2(G1698), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(new_n255), .B1(G33), .B2(G294), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n406), .B(new_n454), .C1(new_n457), .C2(new_n251), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n356), .ZN(new_n459));
  INV_X1    g0259(.A(new_n455), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n226), .A2(G1698), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n460), .A2(new_n364), .A3(new_n366), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G294), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n251), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n465), .A2(new_n262), .A3(new_n406), .A4(new_n454), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n285), .A2(KEYINPUT75), .A3(new_n419), .A4(new_n281), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT75), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n420), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n470), .A3(G107), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n281), .A2(G107), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT25), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n453), .A2(new_n467), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n458), .A2(G169), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT86), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n465), .A2(G179), .A3(new_n406), .A4(new_n454), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n477), .B1(new_n476), .B2(new_n478), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n453), .A2(new_n474), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n475), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT76), .B1(new_n367), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n412), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G250), .A2(G1698), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n255), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n357), .A2(G1698), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(new_n364), .A3(new_n366), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT76), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n255), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n485), .A2(new_n489), .A3(new_n493), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n246), .ZN(new_n498));
  OAI211_X1 g0298(.A(G257), .B(new_n251), .C1(new_n396), .C2(new_n404), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n406), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n498), .A2(KEYINPUT78), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT78), .B1(new_n498), .B2(new_n501), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n383), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT71), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n365), .B2(KEYINPUT3), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n363), .A2(KEYINPUT71), .A3(G33), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(new_n366), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n207), .A2(KEYINPUT7), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT7), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n255), .B2(G20), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n368), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n368), .A2(KEYINPUT6), .A3(G97), .ZN(new_n515));
  XNOR2_X1  g0315(.A(G97), .B(G107), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT6), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI22_X1  g0318(.A1(new_n518), .A2(new_n207), .B1(new_n352), .B2(new_n270), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n279), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n468), .A2(new_n470), .A3(G97), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n282), .A2(new_n225), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n498), .A2(new_n300), .A3(new_n501), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT78), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n485), .A2(new_n496), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n412), .B1(new_n367), .B2(new_n487), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT4), .B1(new_n255), .B2(new_n490), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n251), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n527), .B1(new_n532), .B2(new_n500), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n500), .B1(new_n246), .B2(new_n497), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT78), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n535), .A3(G190), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n356), .B1(new_n498), .B2(new_n501), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n524), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n504), .A2(new_n526), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n348), .B(KEYINPUT82), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(new_n470), .A3(new_n468), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT19), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n207), .B1(new_n306), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n220), .A2(new_n225), .A3(new_n368), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n364), .A2(new_n366), .A3(new_n207), .A4(G68), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n542), .B1(new_n276), .B2(new_n225), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n279), .ZN(new_n549));
  INV_X1    g0349(.A(new_n348), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n282), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n541), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n399), .B(new_n247), .C1(KEYINPUT79), .C2(new_n221), .ZN(new_n553));
  NAND2_X1  g0353(.A1(KEYINPUT79), .A2(G250), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n398), .B2(G1), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n553), .A2(KEYINPUT80), .A3(new_n251), .A4(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n206), .A2(new_n247), .A3(G45), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n221), .A2(KEYINPUT79), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n555), .B(new_n251), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT80), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n365), .A2(new_n414), .ZN(new_n563));
  NOR2_X1   g0363(.A1(G238), .A2(G1698), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n357), .B2(G1698), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n563), .B1(new_n565), .B2(new_n255), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT81), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n246), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n219), .A2(new_n257), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n357), .A2(G1698), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n364), .A2(new_n569), .A3(new_n366), .A4(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n563), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n562), .B(new_n300), .C1(new_n568), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n571), .A2(new_n572), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n251), .B1(new_n576), .B2(KEYINPUT81), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(new_n573), .B1(new_n556), .B2(new_n561), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n552), .B(new_n575), .C1(new_n578), .C2(G169), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n562), .B(G190), .C1(new_n568), .C2(new_n574), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n468), .A2(new_n470), .A3(G87), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n581), .A2(new_n549), .A3(new_n551), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n580), .B(new_n582), .C1(new_n578), .C2(new_n356), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n438), .A2(new_n483), .A3(new_n539), .A4(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n275), .A2(new_n333), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n281), .B2(new_n275), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(G159), .B1(new_n268), .B2(new_n269), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G58), .A2(G68), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n203), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G20), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT70), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G159), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT65), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(new_n207), .A3(new_n365), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n594), .B1(new_n596), .B2(new_n267), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n207), .B1(new_n203), .B2(new_n590), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT70), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n202), .B1(new_n511), .B2(new_n513), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT16), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n509), .B1(new_n364), .B2(new_n366), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n365), .A2(KEYINPUT3), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n363), .A2(G33), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n207), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n605), .B1(new_n608), .B2(new_n512), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT16), .B1(new_n609), .B2(new_n202), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n589), .A2(new_n592), .A3(KEYINPUT70), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n599), .B1(new_n597), .B2(new_n598), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n279), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n588), .B1(new_n604), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT72), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT16), .ZN(new_n617));
  AOI21_X1  g0417(.A(G20), .B1(new_n364), .B2(new_n366), .ZN(new_n618));
  OAI22_X1  g0418(.A1(new_n618), .A2(KEYINPUT7), .B1(new_n255), .B2(new_n509), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n619), .B2(G68), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n285), .B1(new_n601), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n617), .B1(new_n613), .B2(new_n602), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n587), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT72), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OR2_X1    g0425(.A1(G223), .A2(G1698), .ZN(new_n626));
  INV_X1    g0426(.A(G226), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G1698), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n364), .A2(new_n626), .A3(new_n366), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(G33), .A2(G87), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT73), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n629), .A2(KEYINPUT73), .A3(new_n630), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n246), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n312), .B1(new_n224), .B2(new_n252), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G169), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n251), .B1(new_n631), .B2(new_n632), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n636), .B1(new_n640), .B2(new_n634), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G179), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n616), .A2(new_n625), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT18), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n635), .A2(new_n262), .A3(new_n637), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(G200), .B2(new_n641), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT74), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT17), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n623), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  AOI211_X1 g0452(.A(G190), .B(new_n636), .C1(new_n640), .C2(new_n634), .ZN(new_n653));
  AOI21_X1  g0453(.A(G200), .B1(new_n635), .B2(new_n637), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n615), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g0456(.A(KEYINPUT74), .B(KEYINPUT17), .Z(new_n657));
  OAI21_X1  g0457(.A(new_n652), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT18), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n616), .A2(new_n625), .A3(new_n659), .A4(new_n643), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n645), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n388), .A2(new_n585), .A3(new_n661), .ZN(G372));
  NOR2_X1   g0462(.A1(new_n388), .A2(new_n661), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n504), .A2(new_n526), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n536), .A2(new_n538), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n664), .A2(new_n584), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n436), .A2(new_n437), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n453), .A2(new_n474), .B1(new_n476), .B2(new_n478), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT21), .B1(new_n411), .B2(new_n423), .ZN(new_n669));
  OR3_X1    g0469(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT87), .ZN(new_n671));
  INV_X1    g0471(.A(new_n475), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n666), .A2(new_n670), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n664), .A2(new_n672), .A3(new_n584), .A4(new_n665), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT87), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n579), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n579), .A2(new_n583), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n678), .B1(new_n664), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n524), .A2(new_n525), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n533), .A2(new_n535), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(new_n383), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n683), .A2(new_n584), .A3(KEYINPUT26), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n677), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n673), .A2(new_n676), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n663), .A2(new_n686), .ZN(new_n687));
  AOI211_X1 g0487(.A(new_n300), .B(new_n636), .C1(new_n640), .C2(new_n634), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n383), .B1(new_n635), .B2(new_n637), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT18), .B1(new_n623), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n615), .A2(new_n643), .A3(new_n659), .ZN(new_n692));
  INV_X1    g0492(.A(new_n385), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n326), .A2(new_n337), .B1(new_n342), .B2(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n623), .A2(new_n647), .A3(new_n651), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n657), .B1(new_n623), .B2(new_n647), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n691), .B(new_n692), .C1(new_n694), .C2(new_n697), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n698), .A2(new_n294), .B1(new_n299), .B2(new_n301), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n687), .A2(new_n699), .ZN(G369));
  AND2_X1   g0500(.A1(new_n436), .A2(new_n437), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n426), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n703), .A2(KEYINPUT88), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(KEYINPUT88), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(KEYINPUT27), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT27), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n704), .A2(new_n708), .A3(new_n705), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(new_n709), .A3(G213), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT89), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n707), .A2(new_n709), .A3(KEYINPUT89), .A4(G213), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G343), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n428), .ZN(new_n717));
  MUX2_X1   g0517(.A(new_n702), .B(new_n438), .S(new_n717), .Z(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G330), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n476), .A2(new_n478), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT86), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n482), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n672), .A2(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n716), .A2(new_n482), .ZN(new_n726));
  INV_X1    g0526(.A(new_n716), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n725), .A2(new_n726), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n720), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n668), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n702), .A2(new_n727), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n483), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n729), .A2(new_n730), .A3(new_n733), .ZN(G399));
  INV_X1    g0534(.A(new_n210), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G41), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n544), .A2(G116), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(G1), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT90), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n739), .A2(new_n740), .B1(new_n213), .B2(new_n737), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n740), .B2(new_n739), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT91), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT28), .Z(new_n744));
  INV_X1    g0544(.A(G330), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT94), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(new_n585), .B2(new_n716), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n664), .A2(new_n584), .A3(new_n665), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n725), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n749), .A2(KEYINPUT94), .A3(new_n438), .A4(new_n727), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT30), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n576), .A2(KEYINPUT81), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(new_n246), .A3(new_n573), .ZN(new_n754));
  INV_X1    g0554(.A(new_n454), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n464), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n754), .A2(new_n562), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT92), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT92), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n754), .A2(new_n759), .A3(new_n562), .A4(new_n756), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n758), .A2(G179), .A3(new_n434), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n752), .B1(new_n761), .B2(new_n682), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n754), .A2(new_n562), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n300), .ZN(new_n764));
  OAI21_X1  g0564(.A(KEYINPUT93), .B1(new_n764), .B2(new_n434), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT93), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n411), .A2(new_n766), .A3(new_n300), .A4(new_n763), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n534), .B1(new_n406), .B2(new_n756), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AND3_X1   g0569(.A1(new_n434), .A2(new_n760), .A3(G179), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n502), .A2(new_n503), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n770), .A2(new_n771), .A3(KEYINPUT30), .A4(new_n758), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n762), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  AND3_X1   g0573(.A1(new_n773), .A2(KEYINPUT31), .A3(new_n716), .ZN(new_n774));
  AOI21_X1  g0574(.A(KEYINPUT31), .B1(new_n773), .B2(new_n716), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n745), .B1(new_n751), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n686), .A2(new_n727), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(KEYINPUT95), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT29), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT95), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n686), .A2(new_n781), .A3(new_n727), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n701), .A2(new_n426), .A3(new_n724), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n784), .A2(new_n539), .A3(new_n584), .A4(new_n672), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n685), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(KEYINPUT29), .A3(new_n727), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n777), .B1(new_n783), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n744), .B1(new_n788), .B2(G1), .ZN(G364));
  AND2_X1   g0589(.A1(new_n207), .A2(G13), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n206), .B1(new_n790), .B2(G45), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n736), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n718), .A2(G330), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n720), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G13), .A2(G33), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT97), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n718), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n215), .B1(G20), .B2(new_n383), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n207), .A2(G179), .ZN(new_n803));
  NOR2_X1   g0603(.A1(G190), .A2(G200), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n594), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT32), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n356), .A2(G190), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n803), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n367), .B(new_n808), .C1(G107), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n262), .A2(G200), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n300), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G20), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n225), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(new_n807), .B2(new_n806), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n262), .A2(new_n356), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n803), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n220), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n207), .A2(new_n300), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n804), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n823), .A2(new_n283), .B1(new_n824), .B2(new_n352), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n822), .A2(new_n809), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n821), .B(new_n825), .C1(G68), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT98), .ZN(new_n829));
  AND3_X1   g0629(.A1(new_n822), .A2(new_n829), .A3(new_n813), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n829), .B1(new_n822), .B2(new_n813), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G58), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n812), .A2(new_n818), .A3(new_n828), .A4(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n823), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n836), .A2(G326), .B1(new_n811), .B2(G283), .ZN(new_n837));
  INV_X1    g0637(.A(new_n824), .ZN(new_n838));
  INV_X1    g0638(.A(new_n805), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G311), .A2(new_n838), .B1(new_n839), .B2(G329), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n367), .B1(new_n820), .B2(new_n392), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G294), .B2(new_n815), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n833), .A2(G322), .ZN(new_n844));
  XNOR2_X1  g0644(.A(KEYINPUT33), .B(G317), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n845), .A2(KEYINPUT99), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(KEYINPUT99), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n846), .A2(new_n847), .A3(new_n827), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n841), .A2(new_n843), .A3(new_n844), .A4(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n802), .B1(new_n835), .B2(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n793), .B(KEYINPUT96), .Z(new_n851));
  NAND2_X1  g0651(.A1(new_n210), .A2(new_n255), .ZN(new_n852));
  INV_X1    g0652(.A(G355), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n852), .A2(new_n853), .B1(G116), .B2(new_n210), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n735), .A2(new_n255), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n398), .B2(new_n214), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n241), .A2(new_n398), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n799), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(new_n801), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n851), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n800), .A2(new_n850), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n795), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(G396));
  NAND4_X1  g0666(.A1(new_n712), .A2(new_n355), .A3(G343), .A4(new_n713), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n378), .A2(new_n385), .A3(new_n867), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n385), .A2(new_n867), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n779), .A2(new_n782), .A3(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n870), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n686), .A2(new_n727), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n777), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n793), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n875), .B2(new_n874), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n802), .A2(new_n797), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n851), .B1(G77), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(G283), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n414), .A2(new_n824), .B1(new_n826), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT100), .ZN(new_n882));
  INV_X1    g0682(.A(G294), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n882), .B1(new_n883), .B2(new_n832), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n836), .A2(G303), .B1(new_n839), .B2(G311), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n368), .B2(new_n820), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n367), .B1(new_n810), .B2(new_n220), .ZN(new_n887));
  NOR4_X1   g0687(.A1(new_n884), .A2(new_n817), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n888), .A2(KEYINPUT101), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(KEYINPUT101), .ZN(new_n890));
  AOI22_X1  g0690(.A1(G137), .A2(new_n836), .B1(new_n838), .B2(G159), .ZN(new_n891));
  INV_X1    g0691(.A(G143), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n891), .B1(new_n266), .B2(new_n826), .C1(new_n832), .C2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n894), .A2(KEYINPUT34), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n255), .B1(new_n820), .B2(new_n283), .ZN(new_n896));
  INV_X1    g0696(.A(G132), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n810), .A2(new_n202), .B1(new_n805), .B2(new_n897), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n896), .B(new_n898), .C1(G58), .C2(new_n815), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT34), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n899), .B1(new_n893), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n889), .B(new_n890), .C1(new_n895), .C2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n879), .B1(new_n902), .B2(new_n801), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n872), .B2(new_n797), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n877), .A2(new_n904), .ZN(G384));
  INV_X1    g0705(.A(new_n518), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n906), .A2(KEYINPUT35), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(KEYINPUT35), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n907), .A2(G116), .A3(new_n216), .A4(new_n908), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT36), .Z(new_n910));
  NAND3_X1  g0710(.A1(new_n214), .A2(G77), .A3(new_n590), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n283), .A2(G68), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n206), .B(G13), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n751), .A2(new_n776), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n716), .A2(new_n337), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n343), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n338), .A2(new_n342), .A3(new_n916), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n870), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n605), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n202), .B1(new_n513), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n617), .B1(new_n613), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n587), .B1(new_n621), .B2(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(new_n714), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n661), .A2(new_n926), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n615), .A2(new_n655), .B1(new_n924), .B2(new_n714), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n924), .A2(new_n690), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT37), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT102), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(KEYINPUT102), .B(KEYINPUT37), .C1(new_n928), .C2(new_n929), .ZN(new_n933));
  INV_X1    g0733(.A(new_n714), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n616), .A2(new_n625), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT37), .B1(new_n623), .B2(new_n647), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n644), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n932), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n927), .A2(new_n938), .A3(KEYINPUT38), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT38), .B1(new_n927), .B2(new_n938), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n915), .B(new_n920), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT40), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n915), .A2(new_n920), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n927), .A2(new_n938), .A3(KEYINPUT38), .ZN(new_n944));
  INV_X1    g0744(.A(new_n935), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n691), .A2(new_n692), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n945), .B1(new_n697), .B2(new_n946), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n644), .A2(new_n935), .A3(new_n936), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT37), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n621), .A2(new_n622), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n950), .A2(new_n588), .B1(new_n639), .B2(new_n642), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n656), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n949), .B1(new_n952), .B2(new_n935), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n947), .B1(new_n948), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT38), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n942), .B1(new_n944), .B2(new_n956), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n941), .A2(new_n942), .B1(new_n943), .B2(new_n957), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n958), .A2(new_n663), .A3(new_n915), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n958), .B1(new_n663), .B2(new_n915), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n959), .A2(new_n960), .A3(new_n745), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n918), .A2(new_n919), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n716), .A2(new_n385), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n963), .B1(new_n873), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n927), .A2(new_n938), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n955), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n944), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n966), .A2(new_n969), .B1(new_n946), .B2(new_n714), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n944), .A2(new_n956), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT39), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n968), .A2(KEYINPUT39), .A3(new_n944), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n338), .A2(new_n716), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n970), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n783), .A2(new_n663), .A3(new_n787), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n699), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n977), .B(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n961), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n206), .B2(new_n790), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n961), .A2(new_n980), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n914), .B1(new_n982), .B2(new_n983), .ZN(G367));
  NAND2_X1  g0784(.A1(new_n716), .A2(new_n524), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n539), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n683), .A2(new_n716), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n733), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n664), .B1(new_n986), .B2(new_n724), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n989), .A2(KEYINPUT42), .B1(new_n727), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(KEYINPUT42), .B2(new_n989), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT43), .ZN(new_n993));
  OR3_X1    g0793(.A1(new_n727), .A2(new_n579), .A3(new_n582), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n584), .B1(new_n727), .B2(new_n582), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n992), .B1(new_n993), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n729), .A2(new_n988), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n736), .B(new_n1003), .Z(new_n1004));
  INV_X1    g0804(.A(new_n988), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1005), .A2(new_n730), .A3(new_n733), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT45), .Z(new_n1007));
  AOI21_X1  g0807(.A(new_n1005), .B1(new_n730), .B2(new_n733), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT44), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(new_n729), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n720), .A2(KEYINPUT104), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n733), .B1(new_n728), .B2(new_n732), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1012), .B(new_n1013), .Z(new_n1014));
  NAND3_X1  g0814(.A1(new_n1011), .A2(new_n788), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1004), .B1(new_n1015), .B2(new_n788), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1002), .B1(new_n792), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n856), .A2(new_n237), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n861), .B1(new_n210), .B2(new_n550), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n820), .A2(new_n414), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT46), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT107), .Z(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G303), .B2(new_n833), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G107), .A2(new_n815), .B1(new_n838), .B2(G283), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT105), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n367), .B1(new_n883), .B2(new_n826), .C1(new_n1020), .C2(KEYINPUT46), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n810), .A2(new_n225), .ZN(new_n1027));
  XOR2_X1   g0827(.A(KEYINPUT106), .B(G311), .Z(new_n1028));
  XNOR2_X1  g0828(.A(KEYINPUT108), .B(G317), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n823), .A2(new_n1028), .B1(new_n805), .B2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1026), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1023), .A2(new_n1025), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n820), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT109), .B(G137), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G58), .A2(new_n1033), .B1(new_n839), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n283), .B2(new_n824), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G150), .B2(new_n833), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n823), .A2(new_n892), .B1(new_n826), .B2(new_n594), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n367), .B(new_n1039), .C1(G77), .C2(new_n811), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(new_n202), .C2(new_n816), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1032), .A2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT47), .Z(new_n1043));
  OAI221_X1 g0843(.A(new_n851), .B1(new_n1018), .B2(new_n1019), .C1(new_n1043), .C2(new_n802), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1044), .A2(KEYINPUT110), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(KEYINPUT110), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(new_n799), .C2(new_n996), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1017), .A2(new_n1047), .ZN(G387));
  NAND2_X1  g0848(.A1(new_n1014), .A2(new_n792), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n540), .A2(new_n815), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n275), .B2(new_n826), .C1(new_n283), .C2(new_n832), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n836), .A2(G159), .B1(new_n839), .B2(G150), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1033), .A2(G77), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(new_n202), .C2(new_n824), .ZN(new_n1054));
  NOR4_X1   g0854(.A1(new_n1051), .A2(new_n1054), .A3(new_n367), .A4(new_n1027), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT112), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1028), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n827), .A2(new_n1057), .B1(new_n836), .B2(G322), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n392), .B2(new_n824), .C1(new_n832), .C2(new_n1029), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT48), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G283), .A2(new_n815), .B1(new_n1033), .B2(G294), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT113), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(KEYINPUT49), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n255), .B1(new_n839), .B2(G326), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(new_n414), .C2(new_n810), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1065), .A2(KEYINPUT49), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1056), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n801), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n851), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n852), .A2(new_n738), .B1(G107), .B2(new_n210), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n234), .A2(new_n398), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n738), .ZN(new_n1075));
  AOI211_X1 g0875(.A(G45), .B(new_n1075), .C1(G68), .C2(G77), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n271), .A2(G50), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT50), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n856), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1073), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1080), .A2(KEYINPUT111), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n862), .B1(new_n1080), .B2(KEYINPUT111), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1072), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1071), .B(new_n1083), .C1(new_n728), .C2(new_n799), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1014), .A2(new_n788), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n736), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1014), .A2(new_n788), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1049), .B(new_n1084), .C1(new_n1086), .C2(new_n1087), .ZN(G393));
  INV_X1    g0888(.A(new_n1011), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT114), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n791), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n1090), .B2(new_n1089), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1089), .A2(new_n1085), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1093), .A2(new_n736), .A3(new_n1015), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n816), .A2(new_n352), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n824), .A2(new_n271), .B1(new_n805), .B2(new_n892), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n283), .A2(new_n826), .B1(new_n820), .B2(new_n202), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n255), .B1(new_n810), .B2(new_n220), .ZN(new_n1098));
  NOR4_X1   g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n833), .A2(G159), .B1(G150), .B2(new_n836), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT51), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1099), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1104), .A2(KEYINPUT115), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(KEYINPUT115), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n833), .A2(G311), .B1(G317), .B2(new_n836), .ZN(new_n1108));
  XOR2_X1   g0908(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n1109));
  XNOR2_X1  g0909(.A(new_n1108), .B(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G294), .A2(new_n838), .B1(new_n839), .B2(G322), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n880), .B2(new_n820), .C1(new_n392), .C2(new_n826), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n367), .B1(new_n810), .B2(new_n368), .C1(new_n816), .C2(new_n414), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1107), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n801), .B1(new_n1106), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n862), .B1(G97), .B2(new_n735), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n855), .A2(new_n244), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1072), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1116), .B(new_n1119), .C1(new_n1005), .C2(new_n799), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1092), .A2(new_n1094), .A3(new_n1120), .ZN(G390));
  NAND3_X1  g0921(.A1(new_n777), .A2(new_n872), .A3(new_n962), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n975), .B1(new_n944), .B2(new_n956), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT117), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n716), .B(new_n870), .C1(new_n685), .C2(new_n785), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n962), .B1(new_n1126), .B2(new_n964), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1125), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n975), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n873), .A2(new_n965), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n962), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1131), .A2(new_n1133), .B1(new_n973), .B2(new_n974), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1123), .B1(new_n1130), .B2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n939), .A2(new_n940), .A3(new_n972), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT39), .B1(new_n944), .B2(new_n956), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n966), .A2(new_n975), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1138), .B(new_n1122), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1140), .A2(new_n791), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n796), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n878), .B1(new_n274), .B2(new_n273), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n824), .A2(new_n225), .B1(new_n810), .B2(new_n202), .ZN(new_n1144));
  OR4_X1    g0944(.A1(new_n255), .A2(new_n1095), .A3(new_n821), .A4(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G107), .A2(new_n827), .B1(new_n839), .B2(G294), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n880), .B2(new_n823), .C1(new_n832), .C2(new_n414), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n820), .A2(new_n266), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT53), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n367), .B1(new_n811), .B2(G50), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(new_n594), .C2(new_n816), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT54), .B(G143), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G128), .A2(new_n836), .B1(new_n838), .B2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n827), .A2(new_n1035), .B1(new_n839), .B2(G125), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n897), .C2(new_n832), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n1145), .A2(new_n1147), .B1(new_n1151), .B2(new_n1156), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1143), .B(new_n1072), .C1(new_n801), .C2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1141), .B1(new_n1142), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT118), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n872), .B1(new_n777), .B2(new_n1160), .ZN(new_n1161));
  AOI211_X1 g0961(.A(KEYINPUT118), .B(new_n745), .C1(new_n751), .C2(new_n776), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n963), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1126), .A2(new_n964), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1122), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n962), .B1(new_n777), .B2(new_n872), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1132), .B1(new_n1123), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n663), .A2(new_n777), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n978), .A2(new_n699), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n1140), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1169), .A2(new_n1135), .A3(new_n1139), .A4(new_n1172), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(new_n736), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1159), .A2(new_n1176), .ZN(G378));
  NAND2_X1  g0977(.A1(new_n941), .A2(new_n942), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n957), .A2(new_n915), .A3(new_n920), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(G330), .A3(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n295), .A2(new_n714), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n294), .A2(new_n302), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1184), .B1(new_n294), .B2(new_n302), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1182), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1187), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(new_n1185), .A3(new_n1181), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1180), .A2(KEYINPUT123), .A3(new_n1191), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1188), .A2(new_n1190), .A3(KEYINPUT122), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT122), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n958), .A2(new_n1195), .A3(G330), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT123), .B1(new_n1180), .B2(new_n1191), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n977), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1180), .A2(new_n1191), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT123), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n977), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1202), .A2(new_n1203), .A3(new_n1196), .A4(new_n1192), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1199), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n796), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n793), .B1(G50), .B2(new_n878), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT121), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n540), .A2(new_n838), .B1(G97), .B2(new_n827), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT120), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G41), .B(new_n255), .C1(new_n836), .C2(G116), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n880), .B2(new_n805), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1053), .B1(new_n201), .B2(new_n810), .C1(new_n816), .C2(new_n202), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1210), .B(new_n1214), .C1(new_n368), .C2(new_n832), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1216), .A2(KEYINPUT58), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(G33), .A2(G41), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT119), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n283), .C1(G41), .C2(new_n255), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1216), .A2(KEYINPUT58), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G125), .A2(new_n836), .B1(new_n827), .B2(G132), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G137), .A2(new_n838), .B1(new_n1033), .B2(new_n1153), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(G128), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1224), .B1(new_n266), .B2(new_n816), .C1(new_n1225), .C2(new_n832), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n810), .A2(new_n594), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1219), .B(new_n1229), .C1(G124), .C2(new_n839), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1217), .A2(new_n1220), .A3(new_n1221), .A4(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1208), .B1(new_n1232), .B2(new_n801), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1205), .A2(new_n792), .B1(new_n1206), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT57), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1175), .B2(new_n1172), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1205), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n736), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1175), .A2(new_n1172), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT57), .B1(new_n1205), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1234), .B1(new_n1238), .B2(new_n1240), .ZN(G375));
  INV_X1    g1041(.A(KEYINPUT125), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n791), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n963), .A2(new_n796), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n851), .B1(G68), .B2(new_n878), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G159), .A2(new_n1033), .B1(new_n827), .B2(new_n1153), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n897), .B2(new_n823), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n833), .B2(new_n1035), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n824), .A2(new_n266), .B1(new_n805), .B2(new_n1225), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n367), .B(new_n1249), .C1(G58), .C2(new_n811), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1248), .B(new_n1250), .C1(new_n283), .C2(new_n816), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1050), .B1(new_n880), .B2(new_n832), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT124), .Z(new_n1253));
  AOI22_X1  g1053(.A1(G294), .A2(new_n836), .B1(new_n1033), .B2(G97), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G116), .A2(new_n827), .B1(new_n839), .B2(G303), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n838), .A2(G107), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n255), .B1(new_n811), .B2(G77), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1251), .B1(new_n1253), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1245), .B1(new_n1259), .B2(new_n801), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1244), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1242), .B1(new_n1243), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1167), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1122), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1132), .A2(new_n1265), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1266));
  OAI211_X1 g1066(.A(KEYINPUT125), .B(new_n1261), .C1(new_n1266), .C2(new_n791), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1004), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1166), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1173), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1271), .ZN(new_n1272));
  XOR2_X1   g1072(.A(new_n1272), .B(KEYINPUT126), .Z(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(G381));
  NOR2_X1   g1074(.A1(G393), .A2(G396), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(G390), .A2(G384), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(G387), .ZN(new_n1278));
  INV_X1    g1078(.A(G378), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1273), .A2(new_n1277), .A3(new_n1278), .A4(new_n1279), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1280), .A2(G375), .ZN(G407));
  NAND2_X1  g1081(.A1(new_n715), .A2(G213), .ZN(new_n1282));
  OR3_X1    g1082(.A1(G375), .A2(G378), .A3(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(G407), .A2(G213), .A3(new_n1283), .ZN(G409));
  OAI211_X1 g1084(.A(G378), .B(new_n1234), .C1(new_n1238), .C2(new_n1240), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1205), .A2(new_n1269), .A3(new_n1239), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1234), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1279), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1266), .A2(KEYINPUT60), .A3(new_n1171), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT60), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1270), .A2(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1290), .A2(new_n1292), .A3(new_n736), .A4(new_n1173), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1268), .A2(new_n1293), .A3(G384), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(G384), .B1(new_n1268), .B2(new_n1293), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1289), .A2(new_n1282), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(KEYINPUT62), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1289), .A2(new_n1282), .ZN(new_n1300));
  OAI21_X1  g1100(.A(KEYINPUT127), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1268), .A2(new_n1293), .ZN(new_n1302));
  INV_X1    g1102(.A(G384), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT127), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(new_n1305), .A3(new_n1294), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n715), .A2(G213), .A3(G2897), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1301), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1307), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1297), .A2(new_n1305), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1300), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT61), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1289), .A2(new_n1314), .A3(new_n1282), .A4(new_n1297), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1299), .A2(new_n1312), .A3(new_n1313), .A4(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(G390), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(G393), .A2(G396), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1317), .B1(new_n1319), .B2(new_n1275), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(G390), .A2(new_n1276), .A3(new_n1318), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1320), .A2(new_n1278), .A3(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1278), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1316), .A2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT61), .B1(new_n1300), .B2(new_n1311), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1298), .A2(new_n1328), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1289), .A2(KEYINPUT63), .A3(new_n1282), .A4(new_n1297), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1324), .A2(new_n1327), .A3(new_n1329), .A4(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1326), .A2(new_n1331), .ZN(G405));
  NAND2_X1  g1132(.A1(G375), .A2(new_n1279), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1285), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1334), .A2(new_n1297), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1297), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1325), .B1(new_n1335), .B2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1335), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1339), .A2(new_n1324), .A3(new_n1336), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1338), .A2(new_n1340), .ZN(G402));
endmodule


