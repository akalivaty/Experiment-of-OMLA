

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  INV_X1 U324 ( .A(n529), .ZN(n531) );
  XNOR2_X1 U325 ( .A(n471), .B(KEYINPUT122), .ZN(n582) );
  XOR2_X1 U326 ( .A(G36GAT), .B(G190GAT), .Z(n387) );
  INV_X1 U327 ( .A(KEYINPUT95), .ZN(n333) );
  XNOR2_X1 U328 ( .A(n467), .B(KEYINPUT48), .ZN(n529) );
  XNOR2_X1 U329 ( .A(n334), .B(n333), .ZN(n335) );
  NOR2_X1 U330 ( .A1(n494), .A2(n372), .ZN(n530) );
  XNOR2_X1 U331 ( .A(n336), .B(n335), .ZN(n340) );
  INV_X1 U332 ( .A(n582), .ZN(n584) );
  INV_X1 U333 ( .A(KEYINPUT59), .ZN(n474) );
  XOR2_X1 U334 ( .A(KEYINPUT41), .B(n576), .Z(n566) );
  XOR2_X1 U335 ( .A(n346), .B(n345), .Z(n522) );
  XNOR2_X1 U336 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U337 ( .A(n452), .B(KEYINPUT40), .ZN(n453) );
  XNOR2_X1 U338 ( .A(n477), .B(n476), .ZN(G1352GAT) );
  XNOR2_X1 U339 ( .A(n454), .B(n453), .ZN(G1330GAT) );
  XNOR2_X1 U340 ( .A(G134GAT), .B(KEYINPUT81), .ZN(n292) );
  XNOR2_X1 U341 ( .A(n292), .B(KEYINPUT0), .ZN(n359) );
  XOR2_X1 U342 ( .A(KEYINPUT92), .B(G155GAT), .Z(n294) );
  XNOR2_X1 U343 ( .A(G120GAT), .B(G148GAT), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U345 ( .A(G57GAT), .B(KEYINPUT93), .Z(n296) );
  XNOR2_X1 U346 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U348 ( .A(n298), .B(n297), .Z(n309) );
  XOR2_X1 U349 ( .A(KEYINPUT1), .B(KEYINPUT91), .Z(n300) );
  XNOR2_X1 U350 ( .A(KEYINPUT6), .B(KEYINPUT90), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n307) );
  XOR2_X1 U352 ( .A(G113GAT), .B(G1GAT), .Z(n424) );
  XOR2_X1 U353 ( .A(G85GAT), .B(G162GAT), .Z(n302) );
  XNOR2_X1 U354 ( .A(G29GAT), .B(G127GAT), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U356 ( .A(n424), .B(n303), .Z(n305) );
  NAND2_X1 U357 ( .A1(G225GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n359), .B(n310), .ZN(n312) );
  XNOR2_X1 U362 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n311) );
  XOR2_X1 U363 ( .A(n311), .B(KEYINPUT2), .Z(n322) );
  XOR2_X1 U364 ( .A(n312), .B(n322), .Z(n520) );
  XOR2_X1 U365 ( .A(G22GAT), .B(G155GAT), .Z(n398) );
  XOR2_X1 U366 ( .A(KEYINPUT89), .B(KEYINPUT23), .Z(n314) );
  XNOR2_X1 U367 ( .A(KEYINPUT24), .B(KEYINPUT87), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U369 ( .A(n398), .B(n315), .Z(n317) );
  NAND2_X1 U370 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U372 ( .A(n318), .B(G204GAT), .Z(n321) );
  XNOR2_X1 U373 ( .A(G50GAT), .B(KEYINPUT74), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n319), .B(G162GAT), .ZN(n383) );
  XNOR2_X1 U375 ( .A(n383), .B(KEYINPUT22), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n330) );
  XOR2_X1 U378 ( .A(KEYINPUT21), .B(G218GAT), .Z(n325) );
  XNOR2_X1 U379 ( .A(KEYINPUT88), .B(G211GAT), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U381 ( .A(G197GAT), .B(n326), .Z(n344) );
  XOR2_X1 U382 ( .A(G78GAT), .B(G148GAT), .Z(n328) );
  XNOR2_X1 U383 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n440) );
  XNOR2_X1 U385 ( .A(n344), .B(n440), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n560) );
  XOR2_X1 U387 ( .A(n387), .B(KEYINPUT94), .Z(n332) );
  NAND2_X1 U388 ( .A1(G226GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U390 ( .A(G169GAT), .B(G8GAT), .Z(n423) );
  XNOR2_X1 U391 ( .A(n423), .B(KEYINPUT96), .ZN(n334) );
  XOR2_X1 U392 ( .A(G92GAT), .B(G64GAT), .Z(n338) );
  XNOR2_X1 U393 ( .A(G176GAT), .B(KEYINPUT73), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U395 ( .A(G204GAT), .B(n339), .Z(n449) );
  XOR2_X1 U396 ( .A(n340), .B(n449), .Z(n346) );
  XOR2_X1 U397 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n342) );
  XNOR2_X1 U398 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U400 ( .A(KEYINPUT17), .B(n343), .Z(n363) );
  XNOR2_X1 U401 ( .A(n363), .B(n344), .ZN(n345) );
  INV_X1 U402 ( .A(n522), .ZN(n499) );
  XOR2_X1 U403 ( .A(G176GAT), .B(G99GAT), .Z(n348) );
  XNOR2_X1 U404 ( .A(G43GAT), .B(G190GAT), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U406 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n350) );
  XNOR2_X1 U407 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U409 ( .A(n352), .B(n351), .Z(n357) );
  XOR2_X1 U410 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n354) );
  NAND2_X1 U411 ( .A1(G227GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U413 ( .A(G113GAT), .B(n355), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U415 ( .A(G120GAT), .B(G71GAT), .Z(n436) );
  XOR2_X1 U416 ( .A(n358), .B(n436), .Z(n361) );
  XOR2_X1 U417 ( .A(G15GAT), .B(G127GAT), .Z(n399) );
  XNOR2_X1 U418 ( .A(n359), .B(n399), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U420 ( .A(n363), .B(n362), .Z(n524) );
  INV_X1 U421 ( .A(n524), .ZN(n563) );
  NOR2_X1 U422 ( .A1(n499), .A2(n563), .ZN(n364) );
  XOR2_X1 U423 ( .A(KEYINPUT99), .B(n364), .Z(n365) );
  NOR2_X1 U424 ( .A1(n560), .A2(n365), .ZN(n366) );
  XOR2_X1 U425 ( .A(KEYINPUT25), .B(n366), .Z(n370) );
  XNOR2_X1 U426 ( .A(n522), .B(KEYINPUT97), .ZN(n367) );
  XNOR2_X1 U427 ( .A(KEYINPUT27), .B(n367), .ZN(n372) );
  NAND2_X1 U428 ( .A1(n563), .A2(n560), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n368), .B(KEYINPUT26), .ZN(n548) );
  NOR2_X1 U430 ( .A1(n372), .A2(n548), .ZN(n369) );
  NOR2_X1 U431 ( .A1(n370), .A2(n369), .ZN(n371) );
  NOR2_X1 U432 ( .A1(n520), .A2(n371), .ZN(n376) );
  XOR2_X1 U433 ( .A(n560), .B(KEYINPUT28), .Z(n502) );
  INV_X1 U434 ( .A(n502), .ZN(n534) );
  INV_X1 U435 ( .A(n520), .ZN(n494) );
  NAND2_X1 U436 ( .A1(n530), .A2(n563), .ZN(n373) );
  NOR2_X1 U437 ( .A1(n534), .A2(n373), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n374), .B(KEYINPUT98), .ZN(n375) );
  NOR2_X1 U439 ( .A1(n376), .A2(n375), .ZN(n481) );
  XOR2_X1 U440 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n378) );
  XNOR2_X1 U441 ( .A(KEYINPUT64), .B(KEYINPUT11), .ZN(n377) );
  XNOR2_X1 U442 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U443 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n380) );
  XNOR2_X1 U444 ( .A(G134GAT), .B(KEYINPUT75), .ZN(n379) );
  XNOR2_X1 U445 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U446 ( .A(n382), .B(n381), .Z(n393) );
  XOR2_X1 U447 ( .A(G92GAT), .B(n383), .Z(n385) );
  NAND2_X1 U448 ( .A1(G232GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n391) );
  XNOR2_X1 U450 ( .A(G99GAT), .B(G85GAT), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n386), .B(KEYINPUT71), .ZN(n439) );
  XOR2_X1 U452 ( .A(n387), .B(n439), .Z(n389) );
  XNOR2_X1 U453 ( .A(G218GAT), .B(G106GAT), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U457 ( .A(KEYINPUT67), .B(KEYINPUT7), .Z(n395) );
  XNOR2_X1 U458 ( .A(G43GAT), .B(G29GAT), .ZN(n394) );
  XNOR2_X1 U459 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U460 ( .A(KEYINPUT8), .B(n396), .ZN(n433) );
  XOR2_X1 U461 ( .A(n397), .B(n433), .Z(n572) );
  XOR2_X1 U462 ( .A(n572), .B(KEYINPUT36), .Z(n583) );
  NOR2_X1 U463 ( .A1(n481), .A2(n583), .ZN(n417) );
  XOR2_X1 U464 ( .A(n398), .B(G78GAT), .Z(n401) );
  XNOR2_X1 U465 ( .A(n399), .B(G211GAT), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n406) );
  XNOR2_X1 U467 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n402), .B(KEYINPUT68), .ZN(n435) );
  XOR2_X1 U469 ( .A(n435), .B(KEYINPUT79), .Z(n404) );
  NAND2_X1 U470 ( .A1(G231GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U471 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U472 ( .A(n406), .B(n405), .Z(n408) );
  XNOR2_X1 U473 ( .A(G183GAT), .B(G71GAT), .ZN(n407) );
  XNOR2_X1 U474 ( .A(n408), .B(n407), .ZN(n416) );
  XOR2_X1 U475 ( .A(KEYINPUT14), .B(G64GAT), .Z(n410) );
  XNOR2_X1 U476 ( .A(G1GAT), .B(G8GAT), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U478 ( .A(KEYINPUT15), .B(KEYINPUT78), .Z(n412) );
  XNOR2_X1 U479 ( .A(KEYINPUT12), .B(KEYINPUT80), .ZN(n411) );
  XNOR2_X1 U480 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U481 ( .A(n414), .B(n413), .Z(n415) );
  XOR2_X1 U482 ( .A(n416), .B(n415), .Z(n478) );
  NAND2_X1 U483 ( .A1(n417), .A2(n478), .ZN(n418) );
  XOR2_X1 U484 ( .A(KEYINPUT37), .B(n418), .Z(n519) );
  XOR2_X1 U485 ( .A(G22GAT), .B(G141GAT), .Z(n420) );
  XNOR2_X1 U486 ( .A(G15GAT), .B(G197GAT), .ZN(n419) );
  XNOR2_X1 U487 ( .A(n420), .B(n419), .ZN(n432) );
  XOR2_X1 U488 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n422) );
  XNOR2_X1 U489 ( .A(KEYINPUT65), .B(KEYINPUT29), .ZN(n421) );
  XNOR2_X1 U490 ( .A(n422), .B(n421), .ZN(n428) );
  XOR2_X1 U491 ( .A(G36GAT), .B(G50GAT), .Z(n426) );
  XNOR2_X1 U492 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U493 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U494 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U495 ( .A1(G229GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U496 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U497 ( .A(n432), .B(n431), .ZN(n434) );
  XOR2_X1 U498 ( .A(n434), .B(n433), .Z(n504) );
  INV_X1 U499 ( .A(n504), .ZN(n564) );
  XOR2_X1 U500 ( .A(n435), .B(KEYINPUT31), .Z(n438) );
  XNOR2_X1 U501 ( .A(n436), .B(KEYINPUT69), .ZN(n437) );
  XNOR2_X1 U502 ( .A(n438), .B(n437), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n440), .B(n439), .ZN(n446) );
  XOR2_X1 U504 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n442) );
  NAND2_X1 U505 ( .A1(G230GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U506 ( .A(n442), .B(n441), .ZN(n444) );
  INV_X1 U507 ( .A(KEYINPUT72), .ZN(n443) );
  XNOR2_X1 U508 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U509 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U510 ( .A(n448), .B(n447), .ZN(n450) );
  XOR2_X1 U511 ( .A(n450), .B(n449), .Z(n462) );
  NAND2_X1 U512 ( .A1(n564), .A2(n462), .ZN(n483) );
  NOR2_X1 U513 ( .A1(n519), .A2(n483), .ZN(n451) );
  XOR2_X1 U514 ( .A(KEYINPUT38), .B(n451), .Z(n501) );
  NOR2_X1 U515 ( .A1(n501), .A2(n563), .ZN(n454) );
  INV_X1 U516 ( .A(G43GAT), .ZN(n452) );
  XOR2_X1 U517 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n473) );
  INV_X1 U518 ( .A(n572), .ZN(n459) );
  INV_X1 U519 ( .A(n478), .ZN(n580) );
  XNOR2_X1 U520 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n456) );
  INV_X1 U521 ( .A(n462), .ZN(n576) );
  NAND2_X1 U522 ( .A1(n564), .A2(n566), .ZN(n455) );
  XNOR2_X1 U523 ( .A(n456), .B(n455), .ZN(n457) );
  NOR2_X1 U524 ( .A1(n580), .A2(n457), .ZN(n458) );
  NAND2_X1 U525 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U526 ( .A(n460), .B(KEYINPUT47), .ZN(n466) );
  NOR2_X1 U527 ( .A1(n478), .A2(n583), .ZN(n461) );
  XNOR2_X1 U528 ( .A(n461), .B(KEYINPUT45), .ZN(n463) );
  NAND2_X1 U529 ( .A1(n463), .A2(n462), .ZN(n464) );
  NOR2_X1 U530 ( .A1(n564), .A2(n464), .ZN(n465) );
  NOR2_X1 U531 ( .A1(n466), .A2(n465), .ZN(n467) );
  XOR2_X1 U532 ( .A(n522), .B(KEYINPUT120), .Z(n468) );
  NOR2_X1 U533 ( .A1(n529), .A2(n468), .ZN(n469) );
  XNOR2_X1 U534 ( .A(n469), .B(KEYINPUT54), .ZN(n470) );
  NAND2_X1 U535 ( .A1(n470), .A2(n494), .ZN(n559) );
  NOR2_X1 U536 ( .A1(n548), .A2(n559), .ZN(n471) );
  NAND2_X1 U537 ( .A1(n582), .A2(n564), .ZN(n472) );
  XNOR2_X1 U538 ( .A(n473), .B(n472), .ZN(n477) );
  XNOR2_X1 U539 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n475) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n485) );
  NOR2_X1 U541 ( .A1(n478), .A2(n572), .ZN(n479) );
  XOR2_X1 U542 ( .A(KEYINPUT16), .B(n479), .Z(n480) );
  NOR2_X1 U543 ( .A1(n481), .A2(n480), .ZN(n482) );
  XOR2_X1 U544 ( .A(KEYINPUT100), .B(n482), .Z(n505) );
  NOR2_X1 U545 ( .A1(n505), .A2(n483), .ZN(n492) );
  NAND2_X1 U546 ( .A1(n520), .A2(n492), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n485), .B(n484), .ZN(G1324GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n487) );
  NAND2_X1 U549 ( .A1(n492), .A2(n522), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U551 ( .A(G8GAT), .B(n488), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U553 ( .A1(n492), .A2(n524), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U555 ( .A(G15GAT), .B(n491), .Z(G1326GAT) );
  NAND2_X1 U556 ( .A1(n534), .A2(n492), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n493), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U558 ( .A1(n494), .A2(n501), .ZN(n498) );
  XOR2_X1 U559 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n496) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n495) );
  XNOR2_X1 U561 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U563 ( .A1(n499), .A2(n501), .ZN(n500) );
  XOR2_X1 U564 ( .A(G36GAT), .B(n500), .Z(G1329GAT) );
  NOR2_X1 U565 ( .A1(n502), .A2(n501), .ZN(n503) );
  XOR2_X1 U566 ( .A(G50GAT), .B(n503), .Z(G1331GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n507) );
  NAND2_X1 U568 ( .A1(n504), .A2(n566), .ZN(n518) );
  NOR2_X1 U569 ( .A1(n505), .A2(n518), .ZN(n513) );
  NAND2_X1 U570 ( .A1(n513), .A2(n520), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n508), .Z(G1332GAT) );
  XOR2_X1 U573 ( .A(G64GAT), .B(KEYINPUT107), .Z(n510) );
  NAND2_X1 U574 ( .A1(n513), .A2(n522), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n513), .A2(n524), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n511), .B(KEYINPUT108), .ZN(n512) );
  XNOR2_X1 U578 ( .A(G71GAT), .B(n512), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U580 ( .A1(n513), .A2(n534), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(n517) );
  XOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT110), .Z(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NOR2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n526) );
  NAND2_X1 U585 ( .A1(n520), .A2(n526), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n526), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n526), .A2(n524), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U591 ( .A1(n534), .A2(n526), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  XOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT113), .Z(n536) );
  NAND2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n547) );
  NOR2_X1 U596 ( .A1(n563), .A2(n547), .ZN(n532) );
  XOR2_X1 U597 ( .A(KEYINPUT112), .B(n532), .Z(n533) );
  NOR2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n542), .A2(n564), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U602 ( .A1(n542), .A2(n566), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n540) );
  NAND2_X1 U605 ( .A1(n542), .A2(n580), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n544) );
  NAND2_X1 U609 ( .A1(n542), .A2(n572), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n546) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT115), .Z(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  XOR2_X1 U613 ( .A(G141GAT), .B(KEYINPUT117), .Z(n550) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n556), .A2(n564), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1344GAT) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n554) );
  XOR2_X1 U618 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n552) );
  NAND2_X1 U619 ( .A1(n556), .A2(n566), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U622 ( .A1(n580), .A2(n556), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n555), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U624 ( .A(G162GAT), .B(KEYINPUT119), .Z(n558) );
  NAND2_X1 U625 ( .A1(n556), .A2(n572), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G1347GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT55), .ZN(n562) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n564), .A2(n573), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n568) );
  NAND2_X1 U633 ( .A1(n573), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(n569), .ZN(G1349GAT) );
  XOR2_X1 U636 ( .A(G183GAT), .B(KEYINPUT121), .Z(n571) );
  NAND2_X1 U637 ( .A1(n573), .A2(n580), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(G1350GAT) );
  XNOR2_X1 U639 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1351GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n578) );
  NAND2_X1 U643 ( .A1(n576), .A2(n582), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U645 ( .A(G204GAT), .B(n579), .Z(G1353GAT) );
  NAND2_X1 U646 ( .A1(n582), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(G218GAT), .B(n587), .Z(G1355GAT) );
endmodule

