//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1194, new_n1195,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT65), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  INV_X1    g0010(.A(G116), .ZN(new_n211));
  INV_X1    g0011(.A(G270), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n214), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n213), .B(new_n218), .C1(G50), .C2(G226), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G87), .A2(G250), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G97), .A2(G257), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT66), .B(G238), .Z(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G68), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  AND2_X1   g0024(.A1(G107), .A2(G264), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n207), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n203), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n210), .B(new_n227), .C1(new_n230), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n212), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  INV_X1    g0042(.A(G50), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n214), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n251));
  INV_X1    g0051(.A(G274), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n251), .ZN(new_n257));
  INV_X1    g0057(.A(G238), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G226), .A2(G1698), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(new_n215), .B2(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n260), .A2(new_n265), .B1(G33), .B2(G97), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n254), .B1(new_n257), .B2(new_n258), .C1(new_n266), .C2(new_n256), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT13), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT70), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n268), .B(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n267), .A2(KEYINPUT13), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT71), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT71), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(new_n267), .B2(KEYINPUT13), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n270), .A2(G179), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n268), .ZN(new_n277));
  OR2_X1    g0077(.A1(new_n277), .A2(new_n271), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT14), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(new_n279), .A3(G169), .ZN(new_n280));
  OAI21_X1  g0080(.A(G169), .B1(new_n277), .B2(new_n271), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT14), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n276), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n228), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n250), .B2(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G68), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n287), .B(KEYINPUT72), .ZN(new_n288));
  INV_X1    g0088(.A(G13), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(G1), .ZN(new_n290));
  INV_X1    g0090(.A(G68), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G20), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT12), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n295), .A2(new_n243), .B1(new_n229), .B2(G68), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n229), .A2(G33), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(new_n216), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n285), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n299), .A2(KEYINPUT11), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(KEYINPUT11), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n288), .B(new_n293), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n283), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT18), .ZN(new_n305));
  XOR2_X1   g0105(.A(KEYINPUT8), .B(G58), .Z(new_n306));
  NAND2_X1  g0106(.A1(new_n290), .A2(G20), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n286), .B2(new_n306), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n263), .A2(new_n229), .A3(new_n264), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT7), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT73), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n229), .A4(new_n264), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n315), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT73), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(G68), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n214), .A2(new_n291), .ZN(new_n320));
  OAI21_X1  g0120(.A(G20), .B1(new_n320), .B2(new_n202), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n294), .A2(G159), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT16), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n284), .A2(new_n228), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n313), .A2(new_n315), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n323), .B1(new_n329), .B2(G68), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n328), .B1(new_n330), .B2(KEYINPUT16), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n310), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G169), .ZN(new_n333));
  OR2_X1    g0133(.A1(G223), .A2(G1698), .ZN(new_n334));
  INV_X1    g0134(.A(G1698), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n265), .B(new_n334), .C1(G226), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G87), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n256), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n253), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n257), .A2(new_n215), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n333), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n256), .B1(new_n336), .B2(new_n337), .ZN(new_n344));
  INV_X1    g0144(.A(G179), .ZN(new_n345));
  NOR4_X1   g0145(.A1(new_n344), .A2(new_n341), .A3(new_n345), .A4(new_n253), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n305), .B1(new_n332), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT16), .B1(new_n319), .B2(new_n324), .ZN(new_n349));
  AND2_X1   g0149(.A1(KEYINPUT3), .A2(G33), .ZN(new_n350));
  NOR2_X1   g0150(.A1(KEYINPUT3), .A2(G33), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT7), .B1(new_n352), .B2(new_n229), .ZN(new_n353));
  OAI21_X1  g0153(.A(G68), .B1(new_n353), .B2(new_n317), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(KEYINPUT16), .A3(new_n324), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n285), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n309), .B1(new_n349), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n340), .A2(G179), .A3(new_n342), .ZN(new_n358));
  NOR3_X1   g0158(.A1(new_n344), .A2(new_n341), .A3(new_n253), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n333), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(KEYINPUT18), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n348), .A2(KEYINPUT74), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G200), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n359), .A2(G190), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n332), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT17), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n332), .A2(KEYINPUT17), .A3(new_n364), .A4(new_n365), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n357), .A2(new_n360), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT74), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(new_n305), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n362), .A2(new_n368), .A3(new_n369), .A4(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n270), .A2(G190), .A3(new_n275), .ZN(new_n374));
  INV_X1    g0174(.A(new_n302), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n278), .A2(G200), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n307), .A2(G77), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n286), .A2(G77), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n306), .A2(new_n294), .B1(G20), .B2(G77), .ZN(new_n381));
  XOR2_X1   g0181(.A(KEYINPUT15), .B(G87), .Z(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n381), .B1(new_n297), .B2(new_n383), .ZN(new_n384));
  AOI211_X1 g0184(.A(new_n379), .B(new_n380), .C1(new_n384), .C2(new_n285), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n222), .A2(G1698), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n386), .B(new_n265), .C1(new_n215), .C2(G1698), .ZN(new_n387));
  INV_X1    g0187(.A(G107), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n256), .B1(new_n352), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n253), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n257), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G244), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OR3_X1    g0193(.A1(new_n393), .A2(KEYINPUT67), .A3(G179), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT67), .B1(new_n393), .B2(G179), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n385), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n333), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NOR4_X1   g0199(.A1(new_n304), .A2(new_n373), .A3(new_n378), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n335), .A2(G222), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G223), .A2(G1698), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n265), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(new_n339), .C1(G77), .C2(new_n265), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n391), .A2(G226), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n254), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(G190), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  XOR2_X1   g0208(.A(new_n408), .B(KEYINPUT68), .Z(new_n409));
  OAI21_X1  g0209(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n410));
  INV_X1    g0210(.A(G150), .ZN(new_n411));
  INV_X1    g0211(.A(new_n306), .ZN(new_n412));
  OAI221_X1 g0212(.A(new_n410), .B1(new_n411), .B2(new_n295), .C1(new_n412), .C2(new_n297), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n285), .B1(G50), .B2(new_n286), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(G50), .B2(new_n307), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT9), .ZN(new_n416));
  OR2_X1    g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n406), .A2(G200), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n415), .B2(new_n416), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n409), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT10), .B1(new_n418), .B2(KEYINPUT69), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n420), .B(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n406), .A2(new_n333), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n406), .A2(G179), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n415), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n393), .A2(G200), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(new_n385), .C1(new_n407), .C2(new_n393), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n423), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n400), .A2(new_n429), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n430), .A2(KEYINPUT75), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(KEYINPUT75), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n217), .A2(G1698), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n265), .B(new_n435), .C1(G238), .C2(G1698), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n262), .A2(new_n211), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n256), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G45), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n440), .A2(new_n252), .A3(G1), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(G250), .B1(new_n440), .B2(G1), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n339), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n333), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n345), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT19), .ZN(new_n449));
  INV_X1    g0249(.A(G97), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT76), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT76), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G97), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n449), .B1(new_n454), .B2(new_n297), .ZN(new_n455));
  NAND3_X1  g0255(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n229), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT76), .B(G97), .ZN(new_n458));
  INV_X1    g0258(.A(G87), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n388), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n457), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n265), .A2(new_n229), .A3(G68), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n455), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n250), .A2(G13), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(new_n229), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n463), .A2(new_n285), .B1(new_n465), .B2(new_n383), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT80), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n328), .B(new_n307), .C1(G1), .C2(new_n262), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n382), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n467), .B1(new_n466), .B2(new_n470), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n447), .B(new_n448), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n446), .A2(G200), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n469), .A2(G87), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n445), .A2(G190), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n474), .A2(new_n466), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n290), .A2(G20), .A3(new_n388), .ZN(new_n479));
  XNOR2_X1  g0279(.A(new_n479), .B(KEYINPUT25), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n469), .B2(G107), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n229), .B(G87), .C1(new_n350), .C2(new_n351), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT22), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT22), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n265), .A2(new_n485), .A3(new_n229), .A4(G87), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n484), .A2(new_n486), .B1(new_n229), .B2(new_n437), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT24), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT83), .B1(new_n388), .B2(G20), .ZN(new_n489));
  XOR2_X1   g0289(.A(new_n489), .B(KEYINPUT23), .Z(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n488), .B1(new_n487), .B2(new_n490), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n285), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT84), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n484), .A2(new_n486), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n437), .A2(new_n229), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(new_n490), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT24), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n491), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(KEYINPUT84), .A3(new_n285), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n482), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n440), .A2(G1), .ZN(new_n504));
  XNOR2_X1  g0304(.A(KEYINPUT5), .B(G41), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n339), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n506), .A2(G264), .ZN(new_n507));
  OR2_X1    g0307(.A1(G250), .A2(G1698), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n265), .B(new_n508), .C1(G257), .C2(new_n335), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G294), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n256), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n505), .A2(new_n441), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT85), .B1(new_n514), .B2(G190), .ZN(new_n515));
  INV_X1    g0315(.A(new_n513), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n507), .A2(new_n511), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT85), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(new_n407), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n515), .B(new_n519), .C1(G200), .C2(new_n517), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n478), .B1(new_n503), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n469), .A2(G116), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n465), .A2(new_n211), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n284), .A2(new_n228), .B1(G20), .B2(new_n211), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n451), .A2(new_n453), .A3(new_n262), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  AND3_X1   g0326(.A1(KEYINPUT79), .A2(G33), .A3(G283), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT79), .B1(G33), .B2(G283), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n229), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(KEYINPUT20), .B(new_n524), .C1(new_n526), .C2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G283), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT79), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(KEYINPUT79), .A2(G33), .A3(G283), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n525), .A2(new_n536), .A3(new_n229), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT20), .B1(new_n537), .B2(new_n524), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n522), .B(new_n523), .C1(new_n531), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n335), .A2(G257), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G264), .A2(G1698), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n540), .B(new_n541), .C1(new_n350), .C2(new_n351), .ZN(new_n542));
  INV_X1    g0342(.A(G303), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n263), .A2(new_n543), .A3(new_n264), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT81), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT81), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(new_n547), .A3(new_n544), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n339), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n516), .B1(new_n506), .B2(G270), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n539), .A2(G169), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(KEYINPUT82), .A2(KEYINPUT21), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n553), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n539), .A2(G169), .A3(new_n551), .A4(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n551), .A2(new_n345), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n539), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n554), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT84), .B1(new_n501), .B2(new_n285), .ZN(new_n560));
  AOI211_X1 g0360(.A(new_n495), .B(new_n328), .C1(new_n500), .C2(new_n491), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n481), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n514), .A2(new_n333), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n517), .A2(new_n345), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n559), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n539), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n551), .A2(G200), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n568), .B(new_n569), .C1(new_n407), .C2(new_n551), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n458), .A2(KEYINPUT6), .A3(new_n388), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT6), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n450), .A2(new_n388), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G97), .A2(G107), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(G20), .B1(G77), .B2(new_n294), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n316), .A2(G107), .A3(new_n318), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n328), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n468), .A2(new_n450), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n307), .A2(G97), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT77), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT78), .B1(new_n583), .B2(KEYINPUT4), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n335), .B(G244), .C1(KEYINPUT78), .C2(KEYINPUT4), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n584), .B1(new_n352), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(G244), .B1(KEYINPUT78), .B2(KEYINPUT4), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(G1698), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT78), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(KEYINPUT77), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(new_n265), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n265), .A2(G250), .A3(G1698), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n586), .A2(new_n592), .A3(new_n593), .A4(new_n536), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n339), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n506), .A2(G257), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n513), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G200), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n582), .B(new_n598), .C1(new_n407), .C2(new_n597), .ZN(new_n599));
  INV_X1    g0399(.A(new_n580), .ZN(new_n600));
  INV_X1    g0400(.A(new_n581), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n577), .A2(new_n578), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n600), .B(new_n601), .C1(new_n602), .C2(new_n328), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n597), .A2(new_n333), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n595), .A2(new_n513), .A3(new_n596), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n345), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n599), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n521), .A2(new_n567), .A3(new_n570), .A4(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n434), .A2(new_n609), .ZN(G372));
  INV_X1    g0410(.A(new_n426), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n303), .B1(new_n378), .B2(new_n398), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n368), .A2(new_n369), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT87), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n357), .A2(new_n615), .A3(new_n360), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n357), .B2(new_n360), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n616), .A2(new_n617), .A3(KEYINPUT88), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT88), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT87), .B1(new_n332), .B2(new_n347), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n357), .A2(new_n615), .A3(new_n360), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n305), .B1(new_n618), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT88), .B1(new_n616), .B2(new_n617), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n620), .A2(new_n619), .A3(new_n621), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(KEYINPUT18), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n614), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n611), .B1(new_n629), .B2(new_n423), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n554), .A2(new_n558), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n556), .B(new_n631), .C1(new_n503), .C2(new_n565), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n632), .A2(new_n521), .A3(new_n608), .ZN(new_n633));
  INV_X1    g0433(.A(new_n473), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n478), .B2(new_n607), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n637), .A2(KEYINPUT26), .A3(new_n473), .A4(new_n477), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n634), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT86), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n633), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI211_X1 g0441(.A(KEYINPUT86), .B(new_n634), .C1(new_n636), .C2(new_n638), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n630), .B1(new_n434), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g0444(.A(new_n644), .B(KEYINPUT89), .Z(G369));
  INV_X1    g0445(.A(KEYINPUT27), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n290), .B2(new_n229), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n464), .A2(KEYINPUT27), .A3(G20), .ZN(new_n648));
  INV_X1    g0448(.A(G213), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G343), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT90), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(new_n568), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n559), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n570), .ZN(new_n655));
  XOR2_X1   g0455(.A(new_n655), .B(KEYINPUT91), .Z(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G330), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n562), .A2(new_n566), .A3(new_n652), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n503), .A2(new_n520), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n503), .B2(new_n652), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n562), .A2(new_n566), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n559), .A2(new_n652), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n658), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n665), .A2(new_n669), .ZN(G399));
  INV_X1    g0470(.A(new_n208), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n458), .A2(G116), .A3(new_n460), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G1), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n231), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n605), .A2(new_n517), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n678), .A2(new_n345), .A3(new_n551), .A4(new_n446), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n557), .A2(new_n605), .A3(new_n512), .A4(new_n445), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n446), .A2(new_n551), .A3(new_n345), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(KEYINPUT30), .A3(new_n512), .A4(new_n605), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n679), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n652), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT31), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n609), .B2(new_n686), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n687), .A2(new_n688), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n633), .ZN(new_n695));
  INV_X1    g0495(.A(new_n639), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n652), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT29), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n652), .B1(new_n641), .B2(new_n642), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(KEYINPUT29), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n694), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n677), .B1(new_n701), .B2(G1), .ZN(G364));
  NOR2_X1   g0502(.A1(new_n289), .A2(G20), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G45), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n673), .A2(G1), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n657), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(G330), .ZN(new_n707));
  INV_X1    g0507(.A(new_n656), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(G13), .A2(G33), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT92), .Z(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n229), .ZN(new_n712));
  XOR2_X1   g0512(.A(new_n712), .B(KEYINPUT93), .Z(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n655), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n228), .B1(G20), .B2(new_n333), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n229), .A2(new_n345), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G200), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G190), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n229), .A2(G179), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n723), .A2(new_n407), .A3(new_n363), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI221_X1 g0525(.A(new_n265), .B1(new_n721), .B2(new_n291), .C1(new_n459), .C2(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n723), .A2(G190), .A3(new_n363), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n388), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G190), .A2(G200), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n722), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G159), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT32), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n718), .A2(new_n730), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n733), .A2(new_n734), .B1(new_n216), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n729), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n718), .A2(G190), .A3(new_n363), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n737), .B1(new_n214), .B2(new_n738), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n726), .B(new_n739), .C1(new_n734), .C2(new_n733), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n407), .A2(G179), .A3(G200), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n229), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n743), .A2(KEYINPUT94), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(KEYINPUT94), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G97), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n719), .A2(new_n407), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n740), .B(new_n748), .C1(new_n243), .C2(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT95), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n265), .B1(new_n724), .B2(G303), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT96), .ZN(new_n754));
  INV_X1    g0554(.A(new_n731), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n727), .A2(G283), .B1(G329), .B2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G317), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT33), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n757), .A2(KEYINPUT33), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n720), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G294), .A2(new_n743), .B1(new_n749), .B2(G326), .ZN(new_n761));
  AND4_X1   g0561(.A1(new_n754), .A2(new_n756), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  INV_X1    g0563(.A(G322), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n762), .B1(new_n763), .B2(new_n735), .C1(new_n764), .C2(new_n738), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n717), .B1(new_n752), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n714), .A2(new_n716), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n245), .A2(G45), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n671), .A2(new_n265), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(new_n440), .B2(new_n232), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n768), .A2(new_n771), .B1(new_n211), .B2(new_n671), .ZN(new_n772));
  NAND3_X1  g0572(.A1(G355), .A2(new_n208), .A3(new_n265), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n705), .B(new_n766), .C1(new_n767), .C2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n709), .B1(new_n715), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(G396));
  NAND3_X1  g0577(.A1(new_n396), .A2(new_n397), .A3(new_n652), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n652), .A2(new_n385), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n428), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n778), .B1(new_n399), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n652), .B(new_n782), .C1(new_n641), .C2(new_n642), .ZN(new_n783));
  INV_X1    g0583(.A(new_n699), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n781), .B(KEYINPUT99), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(new_n693), .ZN(new_n787));
  INV_X1    g0587(.A(new_n705), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n725), .A2(new_n243), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n352), .B1(new_n743), .B2(G58), .ZN(new_n791));
  INV_X1    g0591(.A(new_n738), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G137), .A2(new_n749), .B1(new_n792), .B2(G143), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n793), .B1(new_n411), .B2(new_n721), .C1(new_n732), .C2(new_n735), .ZN(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n791), .B1(new_n291), .B2(new_n728), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G132), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n798), .B2(new_n731), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n790), .B(new_n799), .C1(new_n795), .C2(new_n794), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n750), .A2(new_n543), .ZN(new_n801));
  INV_X1    g0601(.A(new_n735), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G116), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n727), .A2(G87), .ZN(new_n804));
  INV_X1    g0604(.A(G294), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n738), .A2(new_n805), .B1(new_n731), .B2(new_n763), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n265), .B(new_n806), .C1(G107), .C2(new_n724), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n748), .A2(new_n803), .A3(new_n804), .A4(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n801), .B(new_n808), .C1(G283), .C2(new_n720), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n716), .B1(new_n800), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n716), .A2(new_n710), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n216), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n781), .A2(new_n711), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n810), .A2(new_n788), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT98), .Z(new_n815));
  NOR2_X1   g0615(.A1(new_n789), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G384));
  NOR2_X1   g0617(.A1(new_n303), .A2(new_n686), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT101), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n330), .A2(KEYINPUT16), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n309), .B1(new_n356), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n360), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n366), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n650), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n819), .B1(new_n366), .B2(new_n822), .ZN(new_n826));
  OAI21_X1  g0626(.A(KEYINPUT37), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n357), .A2(new_n650), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n366), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(KEYINPUT37), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n370), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n824), .ZN(new_n833));
  AND3_X1   g0633(.A1(new_n373), .A2(KEYINPUT100), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(KEYINPUT100), .B1(new_n373), .B2(new_n833), .ZN(new_n835));
  OAI211_X1 g0635(.A(KEYINPUT38), .B(new_n832), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT39), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n623), .A2(new_n613), .A3(new_n626), .ZN(new_n838));
  INV_X1    g0638(.A(new_n828), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n620), .A2(new_n621), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT37), .B1(new_n840), .B2(new_n829), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n838), .A2(new_n839), .B1(new_n831), .B2(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n836), .B(new_n837), .C1(new_n842), .C2(KEYINPUT38), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT38), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n837), .B1(new_n847), .B2(new_n836), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n844), .A2(new_n848), .A3(KEYINPUT102), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT102), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n373), .A2(new_n833), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT100), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n373), .A2(KEYINPUT100), .A3(new_n833), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT38), .B1(new_n855), .B2(new_n832), .ZN(new_n856));
  INV_X1    g0656(.A(new_n836), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT39), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n850), .B1(new_n858), .B2(new_n843), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n818), .B1(new_n849), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n628), .A2(new_n650), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n302), .B(new_n686), .C1(new_n378), .C2(new_n283), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n686), .A2(new_n302), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n303), .A2(new_n377), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n783), .B2(new_n778), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n847), .A2(new_n836), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n861), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n860), .A2(KEYINPUT103), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT103), .ZN(new_n871));
  INV_X1    g0671(.A(new_n818), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT102), .B1(new_n844), .B2(new_n848), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n858), .A2(new_n850), .A3(new_n843), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n869), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n433), .A2(new_n700), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n630), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n878), .B(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n836), .B1(new_n842), .B2(KEYINPUT38), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT104), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n687), .B2(new_n688), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n685), .A2(KEYINPUT104), .A3(KEYINPUT31), .A4(new_n686), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n690), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n865), .A2(new_n782), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT40), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT105), .B1(new_n887), .B2(new_n888), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n781), .B1(new_n862), .B2(new_n864), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT105), .ZN(new_n894));
  OAI221_X1 g0694(.A(new_n893), .B1(new_n894), .B2(KEYINPUT40), .C1(new_n690), .C2(new_n886), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n868), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n690), .A2(new_n886), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n433), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n897), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(G330), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n881), .B(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n250), .B2(new_n703), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n211), .B1(new_n576), .B2(KEYINPUT35), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(new_n230), .C1(KEYINPUT35), .C2(new_n576), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT36), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n231), .A2(new_n216), .A3(new_n320), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n201), .A2(new_n291), .ZN(new_n908));
  OAI211_X1 g0708(.A(G1), .B(new_n289), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n903), .A2(new_n906), .A3(new_n909), .ZN(G367));
  NAND2_X1  g0710(.A1(new_n704), .A2(G1), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n599), .B(new_n607), .C1(new_n582), .C2(new_n652), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT107), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n912), .B(new_n913), .C1(new_n607), .C2(new_n652), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n637), .A2(KEYINPUT107), .A3(new_n686), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n669), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n917), .B(KEYINPUT45), .Z(new_n918));
  NAND2_X1  g0718(.A1(new_n669), .A2(new_n916), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT44), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n665), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n921), .B(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT110), .B1(new_n663), .B2(new_n667), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n657), .B(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n668), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n701), .B1(new_n923), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n672), .B(KEYINPUT41), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n911), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n922), .A2(new_n916), .ZN(new_n934));
  INV_X1    g0734(.A(new_n916), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n926), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT42), .Z(new_n937));
  OAI21_X1  g0737(.A(new_n607), .B1(new_n916), .B2(new_n662), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT108), .Z(new_n939));
  OAI21_X1  g0739(.A(new_n937), .B1(new_n686), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT109), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n652), .B1(new_n466), .B2(new_n475), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT106), .Z(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n473), .B2(new_n477), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n473), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n946), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n940), .B2(new_n941), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n947), .A2(KEYINPUT43), .A3(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(KEYINPUT43), .B(new_n940), .C1(new_n947), .C2(new_n949), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n934), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n950), .A2(new_n951), .A3(new_n934), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n933), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n767), .B1(new_n208), .B2(new_n383), .C1(new_n240), .C2(new_n770), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n792), .A2(G150), .B1(new_n802), .B2(new_n201), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n957), .B1(new_n732), .B2(new_n721), .C1(new_n746), .C2(new_n291), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n352), .B(new_n958), .C1(G143), .C2(new_n749), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n755), .A2(G137), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n961), .B1(new_n214), .B2(new_n725), .C1(new_n216), .C2(new_n728), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n750), .A2(new_n763), .ZN(new_n963));
  INV_X1    g0763(.A(G283), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n738), .A2(new_n543), .B1(new_n735), .B2(new_n964), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n265), .B(new_n965), .C1(G294), .C2(new_n720), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n724), .A2(G116), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT46), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n743), .A2(G107), .B1(G317), .B2(new_n755), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n727), .A2(new_n458), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n966), .A2(new_n968), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n962), .B1(new_n963), .B2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT47), .Z(new_n973));
  OAI211_X1 g0773(.A(new_n788), .B(new_n956), .C1(new_n973), .C2(new_n717), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n946), .A2(new_n713), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n955), .A2(new_n977), .ZN(G387));
  OAI21_X1  g0778(.A(new_n788), .B1(new_n663), .B2(new_n713), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n720), .A2(G311), .B1(new_n802), .B2(G303), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n757), .B2(new_n738), .C1(new_n764), .C2(new_n750), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT48), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n982), .B1(new_n964), .B2(new_n742), .C1(new_n805), .C2(new_n725), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT49), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n265), .B1(new_n755), .B2(G326), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n984), .B(new_n985), .C1(new_n211), .C2(new_n728), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n746), .A2(new_n383), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n725), .A2(new_n216), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n728), .A2(new_n450), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n265), .B1(new_n731), .B2(new_n411), .ZN(new_n990));
  NOR4_X1   g0790(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n792), .A2(G50), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n720), .A2(new_n306), .B1(new_n802), .B2(G68), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT112), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n749), .A2(G159), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n991), .A2(new_n992), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n717), .B1(new_n986), .B2(new_n996), .ZN(new_n997));
  OR3_X1    g0797(.A1(new_n412), .A2(KEYINPUT50), .A3(G50), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT50), .B1(new_n412), .B2(G50), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n998), .A2(new_n440), .A3(new_n674), .A4(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n291), .A2(new_n216), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n769), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT111), .Z(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n440), .B2(new_n237), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n265), .A2(new_n208), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1004), .B1(G107), .B2(new_n208), .C1(new_n674), .C2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n979), .B(new_n997), .C1(new_n767), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n929), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1007), .B1(new_n1008), .B2(new_n911), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n672), .B1(new_n1008), .B2(new_n701), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n701), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n929), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1009), .B1(new_n1010), .B2(new_n1012), .ZN(G393));
  AOI22_X1  g0813(.A1(G317), .A2(new_n749), .B1(new_n792), .B2(G311), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT52), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n265), .B(new_n1015), .C1(G294), .C2(new_n802), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n742), .A2(new_n211), .B1(new_n764), .B2(new_n731), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1017), .B(new_n729), .C1(G303), .C2(new_n720), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1016), .B(new_n1018), .C1(new_n964), .C2(new_n725), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT113), .Z(new_n1020));
  AOI22_X1  g0820(.A1(G150), .A2(new_n749), .B1(new_n792), .B2(G159), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT51), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G68), .B2(new_n724), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n802), .A2(new_n306), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n747), .A2(G77), .B1(G87), .B2(new_n727), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n352), .B1(new_n755), .B2(G143), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n201), .B2(new_n720), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n716), .B1(new_n1020), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n454), .A2(new_n208), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n248), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n767), .B1(new_n1031), .B2(new_n770), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1029), .B(new_n788), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT114), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n713), .B2(new_n935), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1008), .A2(new_n701), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n673), .B1(new_n1039), .B2(new_n923), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n923), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n1012), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1038), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n911), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(G390));
  OAI21_X1  g0845(.A(KEYINPUT115), .B1(new_n867), .B2(new_n818), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n783), .A2(new_n778), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n865), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT115), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n1049), .A3(new_n872), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n873), .A2(new_n874), .A3(new_n1046), .A4(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n399), .A2(new_n780), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n697), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n399), .B2(new_n652), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n882), .B(new_n872), .C1(new_n1054), .C2(new_n866), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n887), .A2(new_n707), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n893), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n693), .A2(new_n888), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n898), .A2(KEYINPUT116), .A3(G330), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT116), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n887), .B2(new_n707), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n785), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1060), .B1(new_n1064), .B2(new_n866), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n1054), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n865), .B1(new_n694), .B2(new_n782), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1058), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1047), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n433), .A2(G330), .A3(new_n898), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1071), .A2(new_n630), .A3(new_n879), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1051), .A2(new_n1055), .A3(new_n1060), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1059), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1071), .A2(new_n630), .A3(new_n879), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n1051), .A2(new_n1055), .A3(new_n1060), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1068), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1075), .A2(new_n1080), .A3(new_n672), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1059), .A2(new_n1074), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n911), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n873), .A2(new_n711), .A3(new_n874), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n746), .A2(new_n216), .B1(new_n211), .B2(new_n738), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT119), .Z(new_n1086));
  AOI21_X1  g0886(.A(new_n265), .B1(new_n724), .B2(G87), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT118), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n728), .A2(new_n291), .B1(new_n731), .B2(new_n805), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n388), .B2(new_n721), .C1(new_n964), .C2(new_n750), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n458), .B2(new_n802), .ZN(new_n1092));
  XOR2_X1   g0892(.A(KEYINPUT54), .B(G143), .Z(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1094), .A2(new_n735), .B1(new_n798), .B2(new_n738), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n724), .A2(G150), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1096), .B(new_n1097), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1095), .B(new_n1098), .C1(G159), .C2(new_n747), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n749), .A2(G128), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n201), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n728), .A2(new_n1101), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n352), .B(new_n1102), .C1(G137), .C2(new_n720), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1099), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G125), .B2(new_n755), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n716), .B1(new_n1092), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1084), .A2(new_n788), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n412), .B2(new_n811), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1081), .A2(new_n1083), .A3(new_n1109), .ZN(G378));
  NAND2_X1  g0910(.A1(new_n423), .A2(new_n426), .ZN(new_n1111));
  XOR2_X1   g0911(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n415), .A2(new_n650), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1112), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n423), .A2(new_n426), .A3(new_n1116), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1113), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1115), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n707), .B(new_n1120), .C1(new_n891), .C2(new_n896), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n897), .A2(G330), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1120), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT103), .B1(new_n860), .B2(new_n869), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n875), .A2(new_n871), .A3(new_n876), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1120), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n897), .B2(G330), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(new_n1121), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(new_n870), .A3(new_n877), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n911), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1129), .A2(new_n711), .B1(new_n1101), .B2(new_n811), .ZN(new_n1135));
  INV_X1    g0935(.A(G124), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n262), .B1(new_n731), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n747), .A2(G150), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n749), .A2(G125), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n792), .A2(G128), .B1(new_n802), .B2(G137), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n724), .A2(new_n1093), .B1(new_n720), .B2(G132), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  AOI211_X1 g0942(.A(G41), .B(new_n1137), .C1(new_n1142), .C2(KEYINPUT59), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(KEYINPUT59), .B2(new_n1142), .C1(new_n732), .C2(new_n728), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n243), .B1(new_n350), .B2(G41), .ZN(new_n1145));
  AOI21_X1  g0945(.A(G41), .B1(new_n792), .B2(G107), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n383), .B2(new_n735), .C1(new_n211), .C2(new_n750), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n352), .B1(new_n731), .B2(new_n964), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G97), .B2(new_n720), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1149), .B1(new_n214), .B2(new_n728), .C1(new_n216), .C2(new_n725), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1147), .B(new_n1150), .C1(G68), .C2(new_n747), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT58), .Z(new_n1152));
  AND3_X1   g0952(.A1(new_n1144), .A2(new_n1145), .A3(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1135), .B(new_n788), .C1(new_n717), .C2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT120), .Z(new_n1155));
  NAND2_X1  g0955(.A1(new_n1134), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1080), .A2(new_n1072), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1133), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT57), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n673), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1133), .A2(new_n1157), .A3(KEYINPUT57), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1156), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(G375));
  AOI21_X1  g0963(.A(new_n705), .B1(new_n291), .B2(new_n811), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT122), .Z(new_n1165));
  NOR2_X1   g0965(.A1(new_n725), .A2(new_n450), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n987), .B1(G77), .B2(new_n727), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n735), .A2(new_n388), .B1(new_n731), .B2(new_n543), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n265), .B(new_n1168), .C1(G116), .C2(new_n720), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(new_n964), .C2(new_n738), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1166), .B(new_n1170), .C1(G294), .C2(new_n749), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n750), .A2(new_n798), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT123), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n1172), .A2(new_n1173), .B1(new_n732), .B2(new_n725), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n265), .B1(new_n721), .B2(new_n1094), .C1(new_n214), .C2(new_n728), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(G137), .C2(new_n792), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n747), .A2(G50), .B1(G150), .B2(new_n802), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G128), .B2(new_n755), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1171), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(new_n717), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1165), .B(new_n1182), .C1(new_n710), .C2(new_n866), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n911), .B(KEYINPUT121), .Z(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n1070), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n931), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1185), .B1(new_n1186), .B2(new_n1077), .ZN(G381));
  NOR2_X1   g0987(.A1(G375), .A2(G378), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n955), .A2(new_n1189), .A3(new_n977), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(G381), .A2(G384), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(G393), .A2(G396), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(G407));
  INV_X1    g0993(.A(G378), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1162), .A2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g0995(.A(G407), .B(G213), .C1(G343), .C2(new_n1195), .ZN(G409));
  INV_X1    g0996(.A(KEYINPUT127), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(G393), .B(new_n776), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1189), .B1(new_n955), .B2(new_n977), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1198), .B1(new_n1190), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(G387), .A2(G390), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n955), .A2(new_n1189), .A3(new_n977), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1198), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1157), .A2(new_n931), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1133), .B1(new_n1206), .B2(new_n1184), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G378), .B1(new_n1207), .B2(new_n1154), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT124), .B1(new_n1162), .B2(G378), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1131), .A2(new_n870), .A3(new_n877), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n870), .A2(new_n877), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1076), .B1(new_n1082), .B2(new_n1077), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1159), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(new_n672), .A3(new_n1161), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1134), .A2(new_n1155), .ZN(new_n1217));
  AND4_X1   g1017(.A1(KEYINPUT124), .A2(new_n1216), .A3(G378), .A4(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1209), .B1(new_n1210), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT62), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1073), .B1(new_n1221), .B2(KEYINPUT60), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT125), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(KEYINPUT60), .ZN(new_n1225));
  OAI211_X1 g1025(.A(KEYINPUT125), .B(new_n1073), .C1(new_n1221), .C2(KEYINPUT60), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1224), .A2(new_n672), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1227), .A2(G384), .A3(new_n1185), .ZN(new_n1228));
  AOI21_X1  g1028(.A(G384), .B1(new_n1227), .B2(new_n1185), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n649), .A2(G343), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1219), .A2(new_n1220), .A3(new_n1230), .A4(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT61), .ZN(new_n1234));
  OAI211_X1 g1034(.A(G2897), .B(new_n1231), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1229), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1227), .A2(G384), .A3(new_n1185), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1231), .A2(G2897), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1235), .A2(new_n1239), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1132), .A2(new_n1128), .B1(new_n1080), .B2(new_n1072), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n672), .B1(new_n1241), .B2(KEYINPUT57), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1161), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1217), .B(G378), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT124), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1216), .A2(KEYINPUT124), .A3(G378), .A4(new_n1217), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1208), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1240), .B1(new_n1248), .B2(new_n1231), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1233), .A2(new_n1234), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1230), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1248), .A2(new_n1251), .A3(new_n1231), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  XOR2_X1   g1053(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1205), .B1(new_n1250), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1231), .B1(new_n1257), .B2(new_n1209), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1249), .A2(KEYINPUT63), .B1(new_n1258), .B2(new_n1230), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1219), .A2(KEYINPUT63), .A3(new_n1230), .A4(new_n1232), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1205), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1259), .A2(new_n1261), .A3(KEYINPUT61), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1197), .B1(new_n1256), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1233), .A2(new_n1234), .A3(new_n1249), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1254), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1252), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1264), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1249), .A2(KEYINPUT63), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1234), .B1(new_n1269), .B2(new_n1252), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1268), .B(KEYINPUT127), .C1(new_n1270), .C2(new_n1261), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1263), .A2(new_n1271), .ZN(G405));
  OAI21_X1  g1072(.A(new_n1257), .B1(G378), .B2(new_n1162), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1264), .B(new_n1273), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(new_n1230), .ZN(G402));
endmodule


