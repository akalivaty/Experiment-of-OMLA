//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n567, new_n568, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(G137), .A3(new_n466), .ZN(new_n467));
  XOR2_X1   g042(.A(new_n467), .B(KEYINPUT66), .Z(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n466), .A2(G2104), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n474), .A2(G2105), .B1(G101), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT67), .ZN(G160));
  NOR2_X1   g053(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n466), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n466), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI22_X1  g060(.A1(new_n482), .A2(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(G2105), .B1(new_n479), .B2(new_n481), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT69), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(new_n488), .B2(G124), .ZN(G162));
  NAND3_X1  g064(.A1(new_n465), .A2(G126), .A3(G2105), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n466), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n466), .A2(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT70), .B1(new_n472), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n466), .A2(G138), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n496), .B(new_n497), .C1(new_n471), .C2(new_n470), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n495), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n494), .B1(new_n463), .B2(new_n464), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT72), .B(KEYINPUT4), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n499), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n495), .A2(KEYINPUT71), .A3(KEYINPUT4), .A4(new_n498), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n493), .B1(new_n503), .B2(new_n504), .ZN(G164));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(new_n508), .ZN(new_n512));
  NAND3_X1  g087(.A1(KEYINPUT73), .A2(KEYINPUT6), .A3(G651), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(G50), .A2(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT74), .B(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n506), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n514), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n509), .B1(new_n518), .B2(KEYINPUT75), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n515), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n512), .A2(new_n513), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT75), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT76), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(new_n523), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n518), .A2(KEYINPUT75), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n526), .A2(new_n527), .A3(new_n528), .A4(new_n509), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(new_n529), .ZN(G166));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n521), .A2(new_n506), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n534), .B1(new_n536), .B2(G89), .ZN(new_n537));
  INV_X1    g112(.A(G51), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n514), .A2(KEYINPUT77), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT77), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n521), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(G543), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n537), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(KEYINPUT78), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(KEYINPUT78), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(G168));
  AND3_X1   g121(.A1(new_n539), .A2(G543), .A3(new_n541), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G52), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(new_n506), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n536), .A2(G90), .B1(new_n552), .B2(G651), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n548), .A2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  AOI22_X1  g130(.A1(new_n547), .A2(G43), .B1(G81), .B2(new_n536), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n550), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT79), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n508), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n561), .B1(new_n560), .B2(new_n559), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT80), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT81), .ZN(G188));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(KEYINPUT82), .B2(KEYINPUT9), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n547), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n572), .B(new_n573), .C1(new_n542), .C2(new_n575), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n550), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n536), .A2(G91), .B1(new_n581), .B2(G651), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n577), .A2(new_n578), .A3(new_n582), .ZN(G299));
  INV_X1    g158(.A(G168), .ZN(G286));
  AND2_X1   g159(.A1(new_n525), .A2(new_n529), .ZN(G303));
  OAI21_X1  g160(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n586));
  INV_X1    g161(.A(G87), .ZN(new_n587));
  INV_X1    g162(.A(G49), .ZN(new_n588));
  OAI221_X1 g163(.A(new_n586), .B1(new_n587), .B2(new_n535), .C1(new_n542), .C2(new_n588), .ZN(G288));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n590), .A2(new_n535), .B1(new_n591), .B2(new_n508), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  AND2_X1   g168(.A1(G48), .A2(G543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n521), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n521), .A2(KEYINPUT83), .A3(new_n594), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n593), .A2(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n536), .A2(G85), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G47), .ZN(new_n603));
  OAI221_X1 g178(.A(new_n601), .B1(new_n508), .B2(new_n602), .C1(new_n542), .C2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n521), .A2(G92), .A3(new_n506), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT10), .Z(new_n607));
  AOI22_X1  g182(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n508), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n547), .A2(G54), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n605), .B1(new_n613), .B2(G868), .ZN(G284));
  XOR2_X1   g189(.A(G284), .B(KEYINPUT84), .Z(G321));
  NOR2_X1   g190(.A1(G299), .A2(G868), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g192(.A(new_n616), .B1(G168), .B2(G868), .ZN(G280));
  XOR2_X1   g193(.A(KEYINPUT85), .B(G559), .Z(new_n619));
  OAI21_X1  g194(.A(new_n613), .B1(G860), .B2(new_n619), .ZN(G148));
  NAND2_X1  g195(.A1(new_n613), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n465), .A2(new_n475), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2100), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n488), .A2(G123), .ZN(new_n629));
  INV_X1    g204(.A(new_n482), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G135), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT87), .ZN(new_n633));
  AND2_X1   g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  OR3_X1    g210(.A1(new_n466), .A2(KEYINPUT86), .A3(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(KEYINPUT86), .B1(new_n466), .B2(G111), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n629), .B(new_n631), .C1(new_n634), .C2(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(G2096), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(G2096), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n628), .A2(new_n640), .A3(new_n641), .ZN(G156));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT89), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n644), .B(new_n646), .Z(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT88), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2430), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n647), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT90), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XNOR2_X1  g236(.A(G2084), .B(G2090), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT91), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(G2072), .A2(G2078), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n442), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT17), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT92), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n666), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n663), .B(new_n672), .C1(new_n667), .C2(new_n669), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n663), .A2(new_n666), .A3(new_n669), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT18), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT94), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT20), .Z(new_n687));
  NAND2_X1  g262(.A1(new_n680), .A2(new_n681), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n682), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n687), .B(new_n689), .C1(new_n685), .C2(new_n688), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT95), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n694), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n692), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n696), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n697), .A2(new_n701), .ZN(G229));
  OR2_X1    g277(.A1(G6), .A2(G16), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(G305), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT32), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1981), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(G23), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n586), .B1(new_n535), .B2(new_n587), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n547), .B2(G49), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n708), .B1(new_n710), .B2(new_n704), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT97), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n707), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT34), .ZN(new_n718));
  NOR2_X1   g293(.A1(G16), .A2(G22), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G166), .B2(G16), .ZN(new_n720));
  INV_X1    g295(.A(G1971), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n717), .A2(new_n718), .A3(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G24), .B(G290), .S(G16), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1986), .ZN(new_n725));
  OR2_X1    g300(.A1(G25), .A2(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n488), .A2(G119), .ZN(new_n727));
  OAI21_X1  g302(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n728));
  INV_X1    g303(.A(G107), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G2105), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT96), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n630), .A2(G131), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n727), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n726), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT35), .B(G1991), .Z(new_n738));
  AND2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n725), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n723), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n718), .B1(new_n717), .B2(new_n722), .ZN(new_n743));
  OAI21_X1  g318(.A(KEYINPUT36), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n743), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n745), .A2(new_n746), .A3(new_n723), .A4(new_n741), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(new_n466), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT25), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G139), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n750), .B(new_n753), .C1(new_n482), .C2(new_n754), .ZN(new_n755));
  MUX2_X1   g330(.A(G33), .B(new_n755), .S(G29), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2072), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n639), .A2(new_n736), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT31), .B(G11), .Z(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT106), .B(G28), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(KEYINPUT30), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n760), .B2(KEYINPUT30), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR4_X1   g338(.A1(new_n757), .A2(new_n758), .A3(new_n759), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(G160), .A2(G29), .ZN(new_n765));
  INV_X1    g340(.A(G34), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(KEYINPUT24), .ZN(new_n767));
  AOI21_X1  g342(.A(G29), .B1(new_n766), .B2(KEYINPUT24), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(KEYINPUT99), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(KEYINPUT99), .B2(new_n768), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT100), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n765), .A2(G2084), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(KEYINPUT101), .ZN(new_n773));
  INV_X1    g348(.A(G1348), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n613), .A2(G16), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G4), .B2(G16), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n764), .B(new_n773), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n704), .A2(G19), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n563), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1341), .ZN(new_n780));
  INV_X1    g355(.A(G2078), .ZN(new_n781));
  NOR2_X1   g356(.A1(G164), .A2(new_n736), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G27), .B2(new_n736), .ZN(new_n783));
  NOR2_X1   g358(.A1(G168), .A2(new_n704), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n704), .B2(G21), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT105), .B(G1966), .Z(new_n786));
  OAI221_X1 g361(.A(new_n780), .B1(new_n781), .B2(new_n783), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n783), .A2(new_n781), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n772), .B2(KEYINPUT101), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n777), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n785), .A2(new_n786), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT107), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n785), .A2(KEYINPUT107), .A3(new_n786), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n488), .A2(G128), .ZN(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n796));
  INV_X1    g371(.A(G116), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G2105), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n630), .B2(G140), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(KEYINPUT98), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT98), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n795), .A2(new_n802), .A3(new_n799), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G29), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n736), .A2(G26), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT28), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G2067), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n805), .A2(G2067), .A3(new_n807), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n793), .A2(new_n794), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(G2084), .B1(new_n765), .B2(new_n771), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n774), .B2(new_n776), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n704), .A2(G20), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT23), .Z(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G299), .B2(G16), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1956), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n704), .A2(G5), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G171), .B2(new_n704), .ZN(new_n820));
  INV_X1    g395(.A(G1961), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n814), .A2(new_n818), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(G29), .A2(G35), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G162), .B2(G29), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G2090), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT108), .B(KEYINPUT29), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n790), .A2(new_n812), .A3(new_n823), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n736), .A2(G32), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n475), .A2(G105), .ZN(new_n831));
  NAND3_X1  g406(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT103), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT26), .Z(new_n834));
  AOI211_X1 g409(.A(new_n831), .B(new_n834), .C1(G141), .C2(new_n630), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n488), .A2(KEYINPUT102), .A3(G129), .ZN(new_n836));
  AOI21_X1  g411(.A(KEYINPUT102), .B1(new_n488), .B2(G129), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT104), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT104), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n840), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n830), .B1(new_n843), .B2(new_n736), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT27), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(G1996), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(G1996), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n829), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n748), .A2(new_n848), .ZN(G311));
  AND3_X1   g424(.A1(new_n748), .A2(new_n848), .A3(KEYINPUT109), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT109), .B1(new_n748), .B2(new_n848), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(G150));
  NAND2_X1  g427(.A1(new_n536), .A2(G93), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  INV_X1    g429(.A(G55), .ZN(new_n855));
  OAI221_X1 g430(.A(new_n853), .B1(new_n508), .B2(new_n854), .C1(new_n542), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT37), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n613), .A2(G559), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT38), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n856), .A2(KEYINPUT110), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n856), .A2(KEYINPUT110), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n563), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n861), .A2(new_n564), .A3(new_n862), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n860), .B(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n868));
  INV_X1    g443(.A(G860), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n867), .B2(KEYINPUT39), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n858), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT111), .Z(G145));
  INV_X1    g447(.A(KEYINPUT115), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT112), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n755), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT4), .B1(new_n501), .B2(new_n497), .ZN(new_n876));
  INV_X1    g451(.A(new_n498), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n500), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n501), .A2(new_n502), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n504), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n493), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n875), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n804), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n875), .B(G164), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(new_n801), .A3(new_n803), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n842), .ZN(new_n888));
  INV_X1    g463(.A(new_n626), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT113), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n735), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n727), .A2(KEYINPUT113), .A3(new_n734), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(G106), .A2(G2105), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n895), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n896));
  INV_X1    g471(.A(G142), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n896), .B1(new_n482), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(new_n488), .B2(G130), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n891), .A2(new_n889), .A3(new_n892), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n894), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n899), .ZN(new_n902));
  INV_X1    g477(.A(new_n900), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(new_n893), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n884), .A2(new_n839), .A3(new_n841), .A4(new_n886), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n888), .A2(new_n901), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n906), .A2(KEYINPUT114), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(KEYINPUT114), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n639), .B(G160), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(G162), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n888), .A2(new_n905), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n904), .A2(new_n901), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n907), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n912), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n906), .ZN(new_n916));
  AOI21_X1  g491(.A(G37), .B1(new_n916), .B2(new_n910), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n873), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n914), .A2(new_n917), .A3(new_n873), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(KEYINPUT40), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n922));
  INV_X1    g497(.A(new_n920), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n922), .B1(new_n923), .B2(new_n918), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n921), .A2(new_n924), .ZN(G395));
  AND2_X1   g500(.A1(new_n864), .A2(new_n865), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(new_n621), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n612), .B(G299), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT116), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(KEYINPUT41), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n927), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT116), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n927), .A2(new_n937), .A3(new_n929), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n931), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT42), .ZN(new_n940));
  XNOR2_X1  g515(.A(G166), .B(G288), .ZN(new_n941));
  XNOR2_X1  g516(.A(G290), .B(G305), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n941), .B(new_n942), .Z(new_n943));
  INV_X1    g518(.A(KEYINPUT42), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n931), .A2(new_n936), .A3(new_n944), .A4(new_n938), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n940), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n943), .B1(new_n940), .B2(new_n945), .ZN(new_n947));
  OAI21_X1  g522(.A(G868), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G868), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n856), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(G295));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n950), .ZN(G331));
  NAND2_X1  g527(.A1(G286), .A2(G171), .ZN(new_n953));
  NAND2_X1  g528(.A1(G168), .A2(G301), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(new_n866), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n953), .A2(new_n954), .B1(new_n864), .B2(new_n865), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n932), .B(new_n934), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n926), .A2(new_n954), .A3(new_n953), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n955), .A2(new_n866), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n929), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n943), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT117), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT117), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n958), .A2(new_n961), .A3(new_n964), .A4(new_n943), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n943), .B1(new_n958), .B2(new_n961), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(G37), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT118), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT44), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n966), .A2(new_n968), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n970), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n971), .A2(new_n974), .A3(KEYINPUT44), .A4(new_n970), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(G397));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n882), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n468), .A2(G40), .A3(new_n476), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT119), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n984), .B(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n843), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n804), .B(new_n809), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n842), .A2(G1996), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n735), .B(new_n738), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n989), .A2(new_n990), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(G290), .B(G1986), .Z(new_n995));
  AOI21_X1  g570(.A(new_n987), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1956), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n880), .B2(new_n881), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n983), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR3_X1   g575(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n997), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT57), .ZN(new_n1003));
  XNOR2_X1  g578(.A(G299), .B(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n981), .B1(G164), .B2(G1384), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n882), .A2(KEYINPUT45), .A3(new_n979), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT56), .B(G2072), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n983), .A4(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1002), .A2(new_n1004), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1004), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n774), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n998), .A2(new_n983), .A3(new_n809), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n612), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1009), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT61), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1002), .A2(new_n1004), .A3(new_n1008), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n1010), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT123), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT123), .B(new_n1015), .C1(new_n1016), .C2(new_n1010), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1010), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1022), .A2(new_n1009), .A3(KEYINPUT61), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1005), .A2(new_n1006), .A3(new_n988), .A4(new_n983), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n983), .A2(new_n998), .ZN(new_n1025));
  XOR2_X1   g600(.A(KEYINPUT58), .B(G1341), .Z(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n563), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT59), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1011), .A2(new_n1012), .A3(KEYINPUT60), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n612), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT60), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1011), .A2(new_n1012), .A3(KEYINPUT60), .A4(new_n613), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1023), .A2(new_n1030), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1014), .B1(new_n1021), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT124), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT124), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1041), .B(new_n1014), .C1(new_n1021), .C2(new_n1038), .ZN(new_n1042));
  NAND4_X1  g617(.A1(G303), .A2(KEYINPUT120), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n525), .A2(new_n529), .A3(G8), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1043), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1005), .A2(new_n983), .A3(new_n1006), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1050), .A2(new_n721), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1000), .A2(new_n1001), .A3(G2090), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1049), .B(G8), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1976), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT52), .B1(G288), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n710), .A2(G1976), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1025), .A2(new_n1055), .A3(G8), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G8), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n983), .B2(new_n998), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1061), .A2(KEYINPUT121), .A3(new_n1056), .A4(new_n1055), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1056), .ZN(new_n1064));
  INV_X1    g639(.A(new_n599), .ZN(new_n1065));
  OAI21_X1  g640(.A(G1981), .B1(new_n1065), .B2(new_n592), .ZN(new_n1066));
  INV_X1    g641(.A(G1981), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n593), .A2(new_n1067), .A3(new_n599), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1066), .A2(KEYINPUT49), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT49), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1064), .A2(KEYINPUT52), .B1(new_n1071), .B2(new_n1061), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1053), .A2(new_n1063), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1052), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1050), .A2(new_n721), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1049), .B1(new_n1076), .B2(G8), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1005), .A2(new_n1006), .A3(new_n781), .A4(new_n983), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n980), .A2(KEYINPUT50), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n998), .A2(new_n999), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n983), .A3(new_n1082), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1080), .A2(KEYINPUT53), .B1(new_n1083), .B2(new_n821), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1079), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(G301), .A3(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1088), .A2(G1961), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1086), .ZN(new_n1090));
  OAI21_X1  g665(.A(G171), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT51), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1050), .A2(new_n786), .ZN(new_n1097));
  INV_X1    g672(.A(G2084), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1081), .A2(new_n1098), .A3(new_n983), .A4(new_n1082), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(G168), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1060), .B1(KEYINPUT125), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1096), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(G8), .A3(G286), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1100), .A2(new_n1102), .A3(new_n1096), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1087), .A2(new_n1091), .A3(KEYINPUT54), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1078), .A2(new_n1094), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1040), .A2(new_n1042), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1049), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1113), .B1(new_n1114), .B2(new_n1060), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1063), .A2(new_n1072), .ZN(new_n1116));
  AOI211_X1 g691(.A(new_n1060), .B(G286), .C1(new_n1097), .C2(new_n1099), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1115), .A2(new_n1053), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(KEYINPUT122), .A2(KEYINPUT63), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1063), .A2(new_n1072), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1060), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(new_n1122), .B2(new_n1049), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1119), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1123), .A2(new_n1115), .A3(new_n1124), .A4(new_n1117), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1073), .A2(new_n1091), .A3(new_n1077), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1104), .A2(new_n1128), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1107), .A2(new_n1106), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT62), .B1(new_n1130), .B2(new_n1103), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1127), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1053), .A2(new_n1121), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1061), .A2(new_n1071), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(new_n1054), .A3(new_n710), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1068), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1061), .B2(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1126), .A2(new_n1132), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n996), .B1(new_n1112), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n986), .A2(new_n988), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT46), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n987), .B1(new_n990), .B2(new_n843), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT47), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1143), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1140), .B(KEYINPUT46), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT47), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT126), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1144), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1146), .A2(new_n1147), .A3(KEYINPUT47), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n727), .A2(new_n734), .A3(new_n738), .ZN(new_n1155));
  OAI22_X1  g730(.A1(new_n1154), .A2(new_n1155), .B1(G2067), .B2(new_n804), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n993), .A2(new_n986), .ZN(new_n1157));
  NOR2_X1   g732(.A1(G290), .A2(G1986), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n986), .A2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT48), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1156), .A2(new_n986), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1149), .A2(new_n1153), .A3(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT127), .B1(new_n1139), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1149), .A2(new_n1153), .A3(new_n1161), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1126), .A2(new_n1132), .A3(new_n1137), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1110), .B1(KEYINPUT124), .B2(new_n1039), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1166), .B1(new_n1167), .B2(new_n1042), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1164), .B(new_n1165), .C1(new_n1168), .C2(new_n996), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1163), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g745(.A1(G227), .A2(new_n461), .ZN(new_n1172));
  NAND4_X1  g746(.A1(new_n697), .A2(new_n701), .A3(new_n660), .A4(new_n1172), .ZN(new_n1173));
  AOI21_X1  g747(.A(new_n1173), .B1(new_n974), .B2(new_n970), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n919), .A2(new_n920), .ZN(new_n1175));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n1175), .ZN(G225));
  INV_X1    g750(.A(G225), .ZN(G308));
endmodule


