//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  AOI22_X1  g002(.A1(new_n203), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n206), .A2(KEYINPUT26), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(new_n207), .B2(new_n203), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT27), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n210), .A2(KEYINPUT68), .A3(G183gat), .ZN(new_n211));
  AND2_X1   g010(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n209), .B(new_n211), .C1(new_n212), .C2(new_n210), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT28), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT27), .B(G183gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(KEYINPUT28), .A3(new_n209), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n208), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G226gat), .A2(G233gat), .ZN(new_n220));
  INV_X1    g019(.A(G183gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(new_n209), .A3(KEYINPUT64), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G183gat), .B2(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT24), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(G183gat), .A3(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n225), .A2(new_n230), .A3(KEYINPUT65), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT65), .B1(new_n225), .B2(new_n230), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT66), .B(KEYINPUT23), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT67), .B1(new_n234), .B2(new_n203), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n236));
  INV_X1    g035(.A(G169gat), .ZN(new_n237));
  INV_X1    g036(.A(G176gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(KEYINPUT23), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(KEYINPUT66), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n236), .B(new_n239), .C1(new_n241), .C2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n206), .B1(KEYINPUT23), .B2(new_n203), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n235), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT25), .B1(new_n233), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n235), .A2(new_n244), .A3(new_n245), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n227), .A2(new_n229), .ZN(new_n249));
  NOR2_X1   g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT25), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n219), .B(new_n220), .C1(new_n247), .C2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G197gat), .B(G204gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT22), .ZN(new_n255));
  INV_X1    g054(.A(G211gat), .ZN(new_n256));
  INV_X1    g055(.A(G218gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(G211gat), .B(G218gat), .Z(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n225), .A2(new_n230), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n205), .B1(new_n239), .B2(new_n242), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n239), .B1(new_n241), .B2(new_n243), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n265), .B1(new_n266), .B2(KEYINPUT67), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n225), .A2(new_n230), .A3(KEYINPUT65), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n264), .A2(new_n267), .A3(new_n244), .A4(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT25), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n252), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n218), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n220), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(KEYINPUT29), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n253), .B(new_n261), .C1(new_n273), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT75), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n252), .B1(new_n270), .B2(new_n269), .ZN(new_n278));
  OAI22_X1  g077(.A1(new_n278), .A2(new_n218), .B1(KEYINPUT29), .B2(new_n274), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT75), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n279), .A2(new_n280), .A3(new_n261), .A4(new_n253), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n253), .B1(new_n273), .B2(new_n275), .ZN(new_n283));
  INV_X1    g082(.A(new_n261), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT74), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n283), .A2(new_n287), .A3(new_n284), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n282), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G8gat), .B(G36gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT76), .ZN(new_n291));
  XNOR2_X1  g090(.A(G64gat), .B(G92gat), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n291), .B(new_n292), .Z(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n293), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n282), .A2(new_n295), .A3(new_n286), .A4(new_n288), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(KEYINPUT30), .A3(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G1gat), .B(G29gat), .Z(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(KEYINPUT0), .ZN(new_n299));
  XNOR2_X1  g098(.A(G57gat), .B(G85gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n301), .B(KEYINPUT85), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT80), .ZN(new_n304));
  OR2_X1    g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT2), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT77), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT2), .ZN(new_n309));
  NAND2_X1  g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n305), .A2(new_n307), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G162gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G155gat), .ZN(new_n313));
  INV_X1    g112(.A(G155gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G162gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT78), .B(G155gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n306), .B1(new_n318), .B2(G162gat), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n305), .A2(new_n313), .A3(new_n315), .A4(new_n310), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n317), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n304), .B1(new_n321), .B2(KEYINPUT3), .ZN(new_n322));
  AND2_X1   g121(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n324));
  OAI21_X1  g123(.A(G162gat), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT2), .ZN(new_n326));
  AND4_X1   g125(.A1(new_n313), .A2(new_n305), .A3(new_n315), .A4(new_n310), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n326), .A2(new_n327), .B1(new_n316), .B2(new_n311), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(KEYINPUT80), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G127gat), .B(G134gat), .ZN(new_n332));
  INV_X1    g131(.A(G113gat), .ZN(new_n333));
  INV_X1    g132(.A(G120gat), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT1), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT69), .B(G120gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G113gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n335), .B1(new_n333), .B2(new_n334), .ZN(new_n339));
  INV_X1    g138(.A(new_n332), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n336), .A2(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n321), .A2(KEYINPUT79), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n313), .A2(new_n315), .ZN(new_n344));
  XOR2_X1   g143(.A(G141gat), .B(G148gat), .Z(new_n345));
  OR2_X1    g144(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n312), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n344), .B(new_n345), .C1(new_n348), .C2(new_n306), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n317), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n343), .A2(KEYINPUT3), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n331), .A2(new_n342), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n341), .A2(new_n328), .A3(KEYINPUT4), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT4), .B1(new_n341), .B2(new_n328), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n353), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n343), .A2(new_n342), .A3(new_n351), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n328), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n354), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT5), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT81), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(new_n360), .ZN(new_n364));
  INV_X1    g163(.A(new_n354), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT5), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n358), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n357), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(KEYINPUT5), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n303), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT40), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n354), .B1(new_n353), .B2(new_n357), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT39), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n302), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT39), .B1(new_n364), .B2(new_n365), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n373), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n379), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n381), .A2(KEYINPUT40), .A3(new_n302), .A4(new_n376), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n372), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n289), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT30), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(new_n295), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n297), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(G78gat), .B(G106gat), .Z(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(G50gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G22gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n261), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n328), .B1(new_n396), .B2(new_n329), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT80), .B1(new_n328), .B2(new_n329), .ZN(new_n398));
  AND4_X1   g197(.A1(KEYINPUT80), .A2(new_n349), .A3(new_n329), .A4(new_n317), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n395), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n397), .B1(new_n400), .B2(new_n284), .ZN(new_n401));
  NAND2_X1  g200(.A1(G228gat), .A2(G233gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n394), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT29), .B1(new_n322), .B2(new_n330), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT3), .B1(new_n261), .B2(new_n395), .ZN(new_n406));
  OAI22_X1  g205(.A1(new_n405), .A2(new_n261), .B1(new_n328), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT83), .A3(new_n402), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n405), .A2(new_n261), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n343), .A2(new_n351), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n403), .B1(new_n411), .B2(new_n406), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n393), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  AOI211_X1 g214(.A(G22gat), .B(new_n413), .C1(new_n404), .C2(new_n408), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n392), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n401), .A2(new_n394), .A3(new_n403), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT83), .B1(new_n407), .B2(new_n402), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n414), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G22gat), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n409), .A2(new_n393), .A3(new_n414), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n422), .A3(new_n391), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n417), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n387), .A2(new_n425), .ZN(new_n426));
  XOR2_X1   g225(.A(KEYINPUT86), .B(KEYINPUT38), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n289), .A2(KEYINPUT37), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT37), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n282), .A2(new_n431), .A3(new_n286), .A4(new_n288), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n293), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n428), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n369), .A2(new_n371), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT6), .B1(new_n435), .B2(new_n301), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n368), .A2(new_n363), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n370), .ZN(new_n438));
  INV_X1    g237(.A(new_n371), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n301), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n436), .A2(new_n372), .B1(KEYINPUT6), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n431), .B1(new_n285), .B2(new_n276), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n442), .A2(new_n295), .A3(new_n428), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n432), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n434), .A2(new_n441), .A3(new_n296), .A4(new_n444), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n417), .A2(new_n423), .A3(KEYINPUT84), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT84), .B1(new_n417), .B2(new_n423), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n297), .A2(new_n386), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n440), .A2(KEYINPUT6), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n438), .A2(new_n301), .A3(new_n439), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n450), .B1(new_n453), .B2(new_n440), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n426), .A2(new_n445), .B1(new_n448), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT34), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n341), .B1(new_n278), .B2(new_n218), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n342), .B(new_n219), .C1(new_n247), .C2(new_n252), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G227gat), .ZN(new_n461));
  INV_X1    g260(.A(G233gat), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n457), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  AOI211_X1 g264(.A(KEYINPUT34), .B(new_n463), .C1(new_n458), .C2(new_n459), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n458), .A2(new_n463), .A3(new_n459), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT32), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT33), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  XOR2_X1   g271(.A(G15gat), .B(G43gat), .Z(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT70), .ZN(new_n474));
  XNOR2_X1  g273(.A(G71gat), .B(G99gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n470), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(KEYINPUT33), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n469), .A2(KEYINPUT32), .A3(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n477), .A2(KEYINPUT71), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT71), .B1(new_n477), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n468), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n460), .A2(new_n464), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT34), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n460), .A2(new_n457), .A3(new_n464), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n479), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n470), .A2(new_n472), .A3(new_n476), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT72), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT72), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n467), .A2(new_n477), .A3(new_n489), .A4(new_n479), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n482), .A2(new_n491), .A3(KEYINPUT36), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT73), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n479), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n468), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n484), .A2(new_n485), .A3(new_n479), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n489), .B1(new_n496), .B2(new_n477), .ZN(new_n497));
  INV_X1    g296(.A(new_n490), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n500), .B1(new_n488), .B2(new_n490), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT73), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(new_n482), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n493), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n482), .A2(new_n491), .A3(new_n423), .A4(new_n417), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT35), .B1(new_n455), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n441), .A2(new_n424), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n491), .A2(new_n495), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT35), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .A4(new_n449), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n456), .A2(new_n505), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(KEYINPUT87), .B(KEYINPUT11), .Z(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT88), .ZN(new_n514));
  XOR2_X1   g313(.A(G113gat), .B(G141gat), .Z(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G169gat), .B(G197gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT12), .ZN(new_n519));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT91), .ZN(new_n521));
  INV_X1    g320(.A(G1gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(KEYINPUT91), .A3(G1gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT16), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(G8gat), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(G29gat), .A2(G36gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT14), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT89), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n530), .B(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT89), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G43gat), .B(G50gat), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n537), .A2(KEYINPUT15), .ZN(new_n538));
  AND2_X1   g337(.A1(G29gat), .A2(G36gat), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n539), .B1(new_n537), .B2(KEYINPUT15), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n532), .A2(new_n536), .A3(new_n538), .A4(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(KEYINPUT15), .B(new_n537), .C1(new_n531), .C2(new_n539), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n541), .A2(KEYINPUT90), .A3(new_n542), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT17), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(KEYINPUT17), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n529), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n545), .A2(new_n528), .A3(new_n546), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT18), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n550), .A2(KEYINPUT18), .A3(new_n551), .A4(new_n552), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(new_n551), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n545), .A2(new_n546), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n529), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n559), .B1(new_n561), .B2(new_n552), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AND4_X1   g362(.A1(new_n519), .A2(new_n555), .A3(new_n556), .A4(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n562), .B1(new_n553), .B2(new_n554), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n519), .B1(new_n565), .B2(new_n556), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n202), .B1(new_n512), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n417), .A2(new_n423), .A3(KEYINPUT84), .ZN(new_n569));
  INV_X1    g368(.A(new_n447), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n455), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n433), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n427), .B1(new_n572), .B2(new_n429), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n372), .A2(new_n451), .A3(new_n452), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n574), .A2(new_n444), .A3(new_n450), .A4(new_n296), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n425), .B(new_n387), .C1(new_n573), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n501), .A2(new_n504), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n503), .B1(new_n502), .B2(new_n482), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n571), .B(new_n576), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n507), .A2(new_n511), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n567), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(KEYINPUT93), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT94), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G64gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n588), .A2(G57gat), .ZN(new_n589));
  INV_X1    g388(.A(G57gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(G64gat), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n587), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G71gat), .B(G78gat), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n589), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(new_n590), .B2(G64gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n588), .A2(KEYINPUT95), .A3(G57gat), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n593), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n595), .A2(KEYINPUT96), .A3(new_n597), .A4(new_n598), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n601), .A2(new_n587), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n594), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT98), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n594), .A2(new_n604), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n606), .A2(KEYINPUT21), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n529), .ZN(new_n611));
  XOR2_X1   g410(.A(G127gat), .B(G155gat), .Z(new_n612));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n611), .B(new_n614), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n605), .A2(KEYINPUT21), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT97), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT99), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n623), .A2(new_n625), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n616), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n623), .A2(new_n625), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n630), .A2(new_n615), .A3(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G190gat), .B(G218gat), .Z(new_n633));
  INV_X1    g432(.A(KEYINPUT104), .ZN(new_n634));
  XNOR2_X1  g433(.A(G99gat), .B(G106gat), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G85gat), .A2(G92gat), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT7), .B1(new_n640), .B2(KEYINPUT101), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(KEYINPUT101), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(G85gat), .A2(G92gat), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT102), .B1(G99gat), .B2(G106gat), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT8), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(KEYINPUT102), .A2(G99gat), .A3(G106gat), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n634), .B(new_n639), .C1(new_n644), .C2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n638), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n635), .A2(new_n636), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n634), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n637), .A2(KEYINPUT104), .A3(new_n638), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n655), .A2(new_n656), .A3(new_n643), .A4(new_n650), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT17), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n560), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n658), .B1(new_n660), .B2(new_n548), .ZN(new_n661));
  NAND2_X1  g460(.A1(G232gat), .A2(G233gat), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(KEYINPUT41), .ZN(new_n664));
  INV_X1    g463(.A(new_n658), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n664), .B1(new_n560), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n633), .B1(new_n661), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n666), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n665), .B1(new_n547), .B2(new_n549), .ZN(new_n669));
  INV_X1    g468(.A(new_n633), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n663), .A2(KEYINPUT41), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT100), .Z(new_n673));
  XNOR2_X1  g472(.A(G134gat), .B(G162gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT105), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n667), .A2(new_n671), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  AOI22_X1  g477(.A1(new_n667), .A2(new_n671), .B1(KEYINPUT105), .B2(new_n675), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n632), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(G120gat), .B(G148gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT106), .ZN(new_n683));
  XNOR2_X1  g482(.A(G176gat), .B(G204gat), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n683), .B(new_n684), .Z(new_n685));
  INV_X1    g484(.A(G230gat), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n462), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n658), .A2(new_n607), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n605), .A2(new_n652), .A3(new_n657), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT10), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n691), .B1(new_n652), .B2(new_n657), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n606), .A2(new_n693), .A3(new_n609), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n687), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n687), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n685), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT10), .B1(new_n688), .B2(new_n689), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n606), .A2(new_n693), .A3(new_n609), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n696), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n685), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n701), .B(new_n702), .C1(new_n696), .C2(new_n690), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n681), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n584), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n454), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(new_n522), .ZN(G1324gat));
  INV_X1    g507(.A(new_n449), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n584), .A2(new_n709), .A3(new_n705), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT108), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT16), .B(G8gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT107), .ZN(new_n714));
  MUX2_X1   g513(.A(KEYINPUT108), .B(new_n712), .S(new_n714), .Z(new_n715));
  NOR2_X1   g514(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n711), .B1(new_n710), .B2(G8gat), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n584), .A2(new_n709), .A3(new_n705), .A4(new_n714), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(G1325gat));
  OAI21_X1  g518(.A(G15gat), .B1(new_n706), .B2(new_n505), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n499), .A2(G15gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n706), .B2(new_n721), .ZN(G1326gat));
  INV_X1    g521(.A(new_n448), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n706), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT43), .B(G22gat), .Z(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1327gat));
  NOR2_X1   g525(.A1(new_n632), .A2(new_n704), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n680), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT93), .B1(new_n581), .B2(new_n582), .ZN(new_n730));
  AOI211_X1 g529(.A(new_n202), .B(new_n567), .C1(new_n579), .C2(new_n580), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n732), .A2(G29gat), .A3(new_n454), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n728), .A2(new_n567), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737));
  INV_X1    g536(.A(new_n680), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n581), .B2(new_n738), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  AOI211_X1 g540(.A(new_n680), .B(new_n741), .C1(new_n579), .C2(new_n580), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n736), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n454), .ZN(new_n746));
  OAI211_X1 g545(.A(KEYINPUT110), .B(new_n736), .C1(new_n739), .C2(new_n742), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G29gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n735), .A2(new_n749), .ZN(G1328gat));
  NOR3_X1   g549(.A1(new_n732), .A2(G36gat), .A3(new_n449), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT46), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n745), .A2(new_n709), .A3(new_n747), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G36gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1329gat));
  OAI21_X1  g554(.A(G43gat), .B1(new_n743), .B2(new_n505), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n499), .A2(G43gat), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n756), .B(KEYINPUT47), .C1(new_n732), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n732), .A2(new_n757), .ZN(new_n759));
  INV_X1    g558(.A(new_n505), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n760), .A3(new_n747), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n759), .B1(new_n761), .B2(G43gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n758), .B1(new_n762), .B2(new_n763), .ZN(G1330gat));
  NOR2_X1   g563(.A1(new_n723), .A2(G50gat), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n729), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n568), .B2(new_n583), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n732), .A2(KEYINPUT112), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G50gat), .B1(new_n743), .B2(new_n425), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(KEYINPUT48), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n745), .A2(new_n448), .A3(new_n747), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n775), .A2(G50gat), .B1(new_n771), .B2(new_n770), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n776), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g576(.A(new_n704), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n681), .A2(new_n582), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n581), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(new_n454), .ZN(new_n781));
  XNOR2_X1  g580(.A(KEYINPUT113), .B(G57gat), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1332gat));
  NOR2_X1   g582(.A1(new_n780), .A2(new_n449), .ZN(new_n784));
  NOR2_X1   g583(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n785));
  AND2_X1   g584(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n784), .B2(new_n785), .ZN(G1333gat));
  OAI21_X1  g587(.A(G71gat), .B1(new_n780), .B2(new_n505), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n499), .A2(G71gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n780), .B2(new_n790), .ZN(new_n791));
  XOR2_X1   g590(.A(new_n791), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g591(.A1(new_n780), .A2(new_n723), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g593(.A1(new_n632), .A2(new_n582), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n704), .ZN(new_n796));
  INV_X1    g595(.A(new_n739), .ZN(new_n797));
  INV_X1    g596(.A(new_n742), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n746), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G85gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n581), .A2(new_n738), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n803), .A2(KEYINPUT51), .A3(new_n795), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT51), .B1(new_n803), .B2(new_n795), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OR3_X1    g605(.A1(new_n454), .A2(new_n778), .A3(G85gat), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n801), .B1(new_n806), .B2(new_n807), .ZN(G1336gat));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809));
  INV_X1    g608(.A(new_n796), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n739), .B2(new_n742), .ZN(new_n811));
  OAI21_X1  g610(.A(G92gat), .B1(new_n811), .B2(new_n449), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n809), .B1(new_n812), .B2(KEYINPUT114), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n449), .A2(G92gat), .A3(new_n778), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n804), .B2(new_n805), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n812), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n815), .B(new_n812), .C1(KEYINPUT114), .C2(new_n809), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1337gat));
  INV_X1    g618(.A(G99gat), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n760), .B(new_n810), .C1(new_n739), .C2(new_n742), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n822), .B2(new_n821), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n509), .A2(new_n820), .A3(new_n704), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n806), .B2(new_n825), .ZN(G1338gat));
  NOR3_X1   g625(.A1(new_n425), .A2(G106gat), .A3(new_n778), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n804), .B2(new_n805), .ZN(new_n828));
  OAI21_X1  g627(.A(G106gat), .B1(new_n811), .B2(new_n723), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831));
  INV_X1    g630(.A(G106gat), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n799), .B2(new_n424), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n828), .A2(new_n831), .ZN(new_n834));
  OAI22_X1  g633(.A1(new_n830), .A2(new_n831), .B1(new_n833), .B2(new_n834), .ZN(G1339gat));
  NAND4_X1  g634(.A1(new_n632), .A2(new_n567), .A3(new_n680), .A4(new_n778), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n692), .A2(new_n687), .A3(new_n694), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n838), .A2(new_n701), .A3(KEYINPUT54), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n685), .B1(new_n701), .B2(KEYINPUT54), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n702), .B1(new_n695), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n838), .A2(new_n701), .A3(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(KEYINPUT55), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n841), .A2(new_n703), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n565), .A2(new_n519), .A3(new_n556), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n551), .B1(new_n550), .B2(new_n552), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n561), .A2(new_n552), .A3(new_n559), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n518), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n847), .B(new_n850), .C1(new_n678), .C2(new_n679), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n704), .A2(new_n847), .A3(new_n850), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n853), .B1(new_n846), .B2(new_n567), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n852), .B1(new_n854), .B2(new_n680), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n836), .B1(new_n855), .B2(new_n632), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT116), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n836), .B(new_n858), .C1(new_n855), .C2(new_n632), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n454), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n506), .A2(new_n709), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(G113gat), .B1(new_n865), .B2(new_n582), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n448), .A2(new_n499), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(new_n454), .A3(new_n709), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n567), .A2(new_n333), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(G1340gat));
  NOR3_X1   g670(.A1(new_n864), .A2(new_n337), .A3(new_n778), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n334), .B1(new_n869), .B2(new_n704), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n872), .A2(new_n873), .ZN(G1341gat));
  INV_X1    g673(.A(G127gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n865), .A2(new_n875), .A3(new_n632), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n869), .A2(new_n632), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n875), .B2(new_n877), .ZN(G1342gat));
  OR2_X1    g677(.A1(new_n680), .A2(G134gat), .ZN(new_n879));
  OR3_X1    g678(.A1(new_n864), .A2(KEYINPUT56), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT56), .B1(new_n864), .B2(new_n879), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n882));
  INV_X1    g681(.A(new_n868), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n709), .A2(new_n454), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n738), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n882), .B1(new_n885), .B2(G134gat), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n885), .A2(new_n882), .A3(G134gat), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n880), .B(new_n881), .C1(new_n886), .C2(new_n887), .ZN(G1343gat));
  AOI21_X1  g687(.A(new_n425), .B1(new_n857), .B2(new_n859), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n505), .A2(new_n884), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n892), .B(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n890), .B1(new_n856), .B2(new_n448), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G141gat), .B1(new_n897), .B2(new_n567), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT119), .B1(new_n861), .B2(new_n454), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n860), .A2(new_n900), .A3(new_n746), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n760), .A2(new_n425), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n449), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n567), .A2(G141gat), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n899), .A2(new_n901), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n898), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT58), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n898), .A2(new_n909), .A3(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1344gat));
  XNOR2_X1  g710(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n912));
  AOI211_X1 g711(.A(new_n778), .B(new_n912), .C1(new_n894), .C2(KEYINPUT121), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n889), .A2(new_n890), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n856), .A2(new_n890), .A3(new_n448), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n894), .A2(KEYINPUT121), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n913), .A2(new_n914), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n897), .A2(new_n778), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(KEYINPUT59), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n704), .A3(new_n899), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n912), .A2(G148gat), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n919), .A2(G148gat), .B1(new_n921), .B2(new_n922), .ZN(G1345gat));
  INV_X1    g722(.A(new_n632), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n318), .B1(new_n897), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n920), .A2(new_n899), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n632), .A2(new_n346), .A3(new_n347), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(G1346gat));
  NOR3_X1   g727(.A1(new_n897), .A2(new_n312), .A3(new_n680), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n920), .A2(new_n738), .A3(new_n899), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(new_n312), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n746), .A2(new_n449), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT123), .Z(new_n933));
  NOR2_X1   g732(.A1(new_n868), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(G169gat), .B1(new_n935), .B2(new_n567), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n860), .A2(new_n932), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n937), .A2(new_n506), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n237), .A3(new_n582), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(G1348gat));
  OAI21_X1  g742(.A(G176gat), .B1(new_n935), .B2(new_n778), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n938), .A2(new_n238), .A3(new_n704), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1349gat));
  AOI21_X1  g745(.A(new_n221), .B1(new_n934), .B2(new_n632), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT60), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n632), .A2(new_n216), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n938), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n948), .A2(KEYINPUT124), .A3(new_n949), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(KEYINPUT124), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT60), .B1(new_n954), .B2(new_n947), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(G1350gat));
  NAND3_X1  g755(.A1(new_n938), .A2(new_n209), .A3(new_n738), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n934), .A2(new_n738), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(G190gat), .ZN(new_n960));
  AOI211_X1 g759(.A(KEYINPUT61), .B(new_n209), .C1(new_n934), .C2(new_n738), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(G1351gat));
  NAND3_X1  g761(.A1(new_n860), .A2(new_n902), .A3(new_n932), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n963), .A2(new_n567), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n933), .A2(new_n760), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n915), .B(new_n965), .C1(new_n889), .C2(new_n890), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n582), .A2(G197gat), .ZN(new_n967));
  OAI22_X1  g766(.A1(new_n964), .A2(G197gat), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(G1352gat));
  OAI21_X1  g768(.A(G204gat), .B1(new_n966), .B2(new_n778), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n778), .A2(G204gat), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT62), .B1(new_n963), .B2(new_n972), .ZN(new_n973));
  OR3_X1    g772(.A1(new_n963), .A2(KEYINPUT62), .A3(new_n972), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n970), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT125), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n970), .A2(new_n974), .A3(new_n977), .A4(new_n973), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(G1353gat));
  OR3_X1    g778(.A1(new_n963), .A2(G211gat), .A3(new_n924), .ZN(new_n980));
  OR2_X1    g779(.A1(new_n966), .A2(new_n924), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n982));
  OAI211_X1 g781(.A(KEYINPUT63), .B(G211gat), .C1(new_n966), .C2(new_n924), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n980), .B1(new_n982), .B2(new_n984), .ZN(G1354gat));
  NOR2_X1   g784(.A1(new_n966), .A2(KEYINPUT127), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n986), .A2(new_n257), .A3(new_n680), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n966), .A2(KEYINPUT127), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n257), .B1(new_n963), .B2(new_n680), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(KEYINPUT126), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n989), .A2(KEYINPUT126), .ZN(new_n991));
  AOI22_X1  g790(.A1(new_n987), .A2(new_n988), .B1(new_n990), .B2(new_n991), .ZN(G1355gat));
endmodule


