

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U551 ( .A1(n589), .A2(n588), .ZN(G164) );
  XNOR2_X1 U552 ( .A(n650), .B(KEYINPUT30), .ZN(n652) );
  NAND2_X1 U553 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U554 ( .A1(n615), .A2(n614), .ZN(n772) );
  NOR2_X2 U555 ( .A1(G2104), .A2(n591), .ZN(n707) );
  XOR2_X1 U556 ( .A(KEYINPUT14), .B(n606), .Z(n519) );
  NOR2_X1 U557 ( .A1(n695), .A2(n685), .ZN(n520) );
  NOR2_X1 U558 ( .A1(n772), .A2(n620), .ZN(n631) );
  INV_X1 U559 ( .A(G168), .ZN(n651) );
  AND2_X1 U560 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U561 ( .A1(n645), .A2(n644), .ZN(n646) );
  INV_X1 U562 ( .A(KEYINPUT105), .ZN(n699) );
  XNOR2_X1 U563 ( .A(n700), .B(n699), .ZN(n701) );
  XOR2_X1 U564 ( .A(KEYINPUT0), .B(G543), .Z(n570) );
  XOR2_X1 U565 ( .A(KEYINPUT1), .B(n521), .Z(n796) );
  NOR2_X1 U566 ( .A1(n570), .A2(G651), .ZN(n797) );
  BUF_X1 U567 ( .A(n772), .Z(n956) );
  NOR2_X1 U568 ( .A1(G543), .A2(G651), .ZN(n802) );
  NAND2_X1 U569 ( .A1(G86), .A2(n802), .ZN(n523) );
  INV_X1 U570 ( .A(G651), .ZN(n524) );
  NOR2_X1 U571 ( .A1(G543), .A2(n524), .ZN(n521) );
  NAND2_X1 U572 ( .A1(G61), .A2(n796), .ZN(n522) );
  NAND2_X1 U573 ( .A1(n523), .A2(n522), .ZN(n528) );
  OR2_X1 U574 ( .A1(n524), .A2(n570), .ZN(n525) );
  XOR2_X2 U575 ( .A(KEYINPUT64), .B(n525), .Z(n801) );
  NAND2_X1 U576 ( .A1(n801), .A2(G73), .ZN(n526) );
  XOR2_X1 U577 ( .A(KEYINPUT2), .B(n526), .Z(n527) );
  NOR2_X1 U578 ( .A1(n528), .A2(n527), .ZN(n530) );
  NAND2_X1 U579 ( .A1(n797), .A2(G48), .ZN(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(G305) );
  NAND2_X1 U581 ( .A1(G89), .A2(n802), .ZN(n531) );
  XOR2_X1 U582 ( .A(KEYINPUT75), .B(n531), .Z(n532) );
  XNOR2_X1 U583 ( .A(n532), .B(KEYINPUT4), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G76), .A2(n801), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U586 ( .A(n535), .B(KEYINPUT5), .ZN(n540) );
  NAND2_X1 U587 ( .A1(G63), .A2(n796), .ZN(n537) );
  NAND2_X1 U588 ( .A1(G51), .A2(n797), .ZN(n536) );
  NAND2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U590 ( .A(KEYINPUT6), .B(n538), .Z(n539) );
  NAND2_X1 U591 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U592 ( .A(n541), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U593 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U594 ( .A1(n797), .A2(G53), .ZN(n542) );
  XNOR2_X1 U595 ( .A(KEYINPUT70), .B(n542), .ZN(n545) );
  NAND2_X1 U596 ( .A1(n796), .A2(G65), .ZN(n543) );
  XOR2_X1 U597 ( .A(KEYINPUT69), .B(n543), .Z(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U599 ( .A(KEYINPUT71), .B(n546), .ZN(n551) );
  NAND2_X1 U600 ( .A1(G91), .A2(n802), .ZN(n548) );
  NAND2_X1 U601 ( .A1(G78), .A2(n801), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U603 ( .A(KEYINPUT68), .B(n549), .Z(n550) );
  NAND2_X1 U604 ( .A1(n551), .A2(n550), .ZN(G299) );
  NAND2_X1 U605 ( .A1(n802), .A2(G90), .ZN(n552) );
  XNOR2_X1 U606 ( .A(n552), .B(KEYINPUT66), .ZN(n554) );
  NAND2_X1 U607 ( .A1(G77), .A2(n801), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U609 ( .A(n555), .B(KEYINPUT9), .ZN(n557) );
  NAND2_X1 U610 ( .A1(G52), .A2(n797), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U612 ( .A1(G64), .A2(n796), .ZN(n558) );
  XNOR2_X1 U613 ( .A(KEYINPUT65), .B(n558), .ZN(n559) );
  NOR2_X1 U614 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U615 ( .A(KEYINPUT67), .B(n561), .Z(G171) );
  INV_X1 U616 ( .A(G171), .ZN(G301) );
  NAND2_X1 U617 ( .A1(G88), .A2(n802), .ZN(n563) );
  NAND2_X1 U618 ( .A1(G75), .A2(n801), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U620 ( .A1(G62), .A2(n796), .ZN(n565) );
  NAND2_X1 U621 ( .A1(G50), .A2(n797), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U623 ( .A1(n567), .A2(n566), .ZN(G166) );
  INV_X1 U624 ( .A(G166), .ZN(G303) );
  NAND2_X1 U625 ( .A1(G74), .A2(G651), .ZN(n568) );
  XOR2_X1 U626 ( .A(KEYINPUT82), .B(n568), .Z(n569) );
  NOR2_X1 U627 ( .A1(n796), .A2(n569), .ZN(n572) );
  NAND2_X1 U628 ( .A1(n570), .A2(G87), .ZN(n571) );
  NAND2_X1 U629 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U630 ( .A1(G49), .A2(n797), .ZN(n573) );
  XNOR2_X1 U631 ( .A(KEYINPUT81), .B(n573), .ZN(n574) );
  NOR2_X1 U632 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U633 ( .A(KEYINPUT83), .B(n576), .ZN(G288) );
  AND2_X1 U634 ( .A1(G72), .A2(n801), .ZN(n580) );
  NAND2_X1 U635 ( .A1(G85), .A2(n802), .ZN(n578) );
  NAND2_X1 U636 ( .A1(G47), .A2(n797), .ZN(n577) );
  NAND2_X1 U637 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U638 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U639 ( .A1(n796), .A2(G60), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n582), .A2(n581), .ZN(G290) );
  NOR2_X1 U641 ( .A1(G2104), .A2(G2105), .ZN(n583) );
  XOR2_X2 U642 ( .A(KEYINPUT17), .B(n583), .Z(n883) );
  NAND2_X1 U643 ( .A1(G138), .A2(n883), .ZN(n589) );
  INV_X1 U644 ( .A(G2105), .ZN(n591) );
  AND2_X1 U645 ( .A1(n591), .A2(G2104), .ZN(n884) );
  AND2_X1 U646 ( .A1(G102), .A2(n884), .ZN(n587) );
  AND2_X1 U647 ( .A1(G2104), .A2(G2105), .ZN(n887) );
  NAND2_X1 U648 ( .A1(G114), .A2(n887), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G126), .A2(n707), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X2 U652 ( .A1(G164), .A2(G1384), .ZN(n703) );
  NAND2_X1 U653 ( .A1(n887), .A2(G113), .ZN(n594) );
  AND2_X1 U654 ( .A1(G2104), .A2(G101), .ZN(n590) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(n592), .B(KEYINPUT23), .Z(n593) );
  AND2_X1 U657 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U658 ( .A1(G125), .A2(n707), .ZN(n595) );
  AND2_X1 U659 ( .A1(n596), .A2(n595), .ZN(n766) );
  AND2_X1 U660 ( .A1(G40), .A2(n766), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n883), .A2(G137), .ZN(n767) );
  NAND2_X1 U662 ( .A1(n597), .A2(n767), .ZN(n704) );
  INV_X1 U663 ( .A(n704), .ZN(n598) );
  NAND2_X2 U664 ( .A1(n703), .A2(n598), .ZN(n661) );
  NAND2_X1 U665 ( .A1(G8), .A2(n661), .ZN(n695) );
  NOR2_X1 U666 ( .A1(G1981), .A2(G305), .ZN(n599) );
  XOR2_X1 U667 ( .A(n599), .B(KEYINPUT24), .Z(n600) );
  NOR2_X1 U668 ( .A1(n695), .A2(n600), .ZN(n702) );
  XOR2_X1 U669 ( .A(KEYINPUT32), .B(KEYINPUT103), .Z(n669) );
  INV_X1 U670 ( .A(n661), .ZN(n641) );
  NAND2_X1 U671 ( .A1(n641), .A2(G2072), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n601), .B(KEYINPUT27), .ZN(n603) );
  AND2_X1 U673 ( .A1(G1956), .A2(n661), .ZN(n602) );
  NOR2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n635) );
  INV_X1 U675 ( .A(G299), .ZN(n810) );
  NOR2_X1 U676 ( .A1(n635), .A2(n810), .ZN(n605) );
  XOR2_X1 U677 ( .A(KEYINPUT98), .B(KEYINPUT28), .Z(n604) );
  XNOR2_X1 U678 ( .A(n605), .B(n604), .ZN(n639) );
  NAND2_X1 U679 ( .A1(n796), .A2(G56), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n802), .A2(G81), .ZN(n607) );
  XNOR2_X1 U681 ( .A(n607), .B(KEYINPUT12), .ZN(n609) );
  NAND2_X1 U682 ( .A1(G68), .A2(n801), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n611) );
  INV_X1 U684 ( .A(KEYINPUT13), .ZN(n610) );
  XNOR2_X1 U685 ( .A(n611), .B(n610), .ZN(n612) );
  NOR2_X1 U686 ( .A1(n519), .A2(n612), .ZN(n613) );
  XNOR2_X1 U687 ( .A(n613), .B(KEYINPUT74), .ZN(n615) );
  NAND2_X1 U688 ( .A1(G43), .A2(n797), .ZN(n614) );
  INV_X1 U689 ( .A(G1996), .ZN(n616) );
  NOR2_X1 U690 ( .A1(n661), .A2(n616), .ZN(n617) );
  XOR2_X1 U691 ( .A(n617), .B(KEYINPUT26), .Z(n619) );
  NAND2_X1 U692 ( .A1(n661), .A2(G1341), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U694 ( .A1(G66), .A2(n796), .ZN(n622) );
  NAND2_X1 U695 ( .A1(G54), .A2(n797), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U697 ( .A1(G92), .A2(n802), .ZN(n624) );
  NAND2_X1 U698 ( .A1(G79), .A2(n801), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(KEYINPUT15), .ZN(n948) );
  NAND2_X1 U702 ( .A1(G1348), .A2(n661), .ZN(n629) );
  NAND2_X1 U703 ( .A1(G2067), .A2(n641), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n632) );
  NOR2_X1 U705 ( .A1(n948), .A2(n632), .ZN(n630) );
  OR2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n948), .A2(n632), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n635), .A2(n810), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U711 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n640), .B(KEYINPUT29), .ZN(n645) );
  NAND2_X1 U713 ( .A1(G1961), .A2(n661), .ZN(n643) );
  XOR2_X1 U714 ( .A(G2078), .B(KEYINPUT25), .Z(n924) );
  NAND2_X1 U715 ( .A1(n641), .A2(n924), .ZN(n642) );
  NAND2_X1 U716 ( .A1(n643), .A2(n642), .ZN(n655) );
  NOR2_X1 U717 ( .A1(G301), .A2(n655), .ZN(n644) );
  XNOR2_X1 U718 ( .A(n646), .B(KEYINPUT99), .ZN(n660) );
  INV_X1 U719 ( .A(KEYINPUT100), .ZN(n654) );
  NOR2_X1 U720 ( .A1(n695), .A2(G1966), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n647), .B(KEYINPUT97), .ZN(n671) );
  INV_X1 U722 ( .A(G8), .ZN(n648) );
  NOR2_X1 U723 ( .A1(G2084), .A2(n661), .ZN(n673) );
  NOR2_X1 U724 ( .A1(n648), .A2(n673), .ZN(n649) );
  AND2_X1 U725 ( .A1(n671), .A2(n649), .ZN(n650) );
  XNOR2_X1 U726 ( .A(n654), .B(n653), .ZN(n657) );
  NAND2_X1 U727 ( .A1(G301), .A2(n655), .ZN(n656) );
  NAND2_X1 U728 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U729 ( .A(n658), .B(KEYINPUT31), .ZN(n659) );
  NAND2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n670) );
  NAND2_X1 U731 ( .A1(G286), .A2(n670), .ZN(n666) );
  NOR2_X1 U732 ( .A1(G1971), .A2(n695), .ZN(n663) );
  NOR2_X1 U733 ( .A1(G2090), .A2(n661), .ZN(n662) );
  NOR2_X1 U734 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U735 ( .A1(n664), .A2(G303), .ZN(n665) );
  NAND2_X1 U736 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U737 ( .A1(G8), .A2(n667), .ZN(n668) );
  XNOR2_X1 U738 ( .A(n669), .B(n668), .ZN(n678) );
  NAND2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U740 ( .A(n672), .B(KEYINPUT101), .ZN(n675) );
  NAND2_X1 U741 ( .A1(n673), .A2(G8), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U743 ( .A(n676), .B(KEYINPUT102), .ZN(n677) );
  NAND2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n693) );
  NOR2_X1 U745 ( .A1(G1976), .A2(G288), .ZN(n943) );
  INV_X1 U746 ( .A(n943), .ZN(n681) );
  NOR2_X1 U747 ( .A1(G1971), .A2(G303), .ZN(n679) );
  XOR2_X1 U748 ( .A(n679), .B(KEYINPUT104), .Z(n680) );
  AND2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n683) );
  INV_X1 U750 ( .A(KEYINPUT33), .ZN(n682) );
  AND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U752 ( .A1(n693), .A2(n684), .ZN(n687) );
  NAND2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n944) );
  INV_X1 U754 ( .A(n944), .ZN(n685) );
  OR2_X1 U755 ( .A1(KEYINPUT33), .A2(n520), .ZN(n686) );
  NAND2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n690) );
  NAND2_X1 U757 ( .A1(n943), .A2(KEYINPUT33), .ZN(n688) );
  NOR2_X1 U758 ( .A1(n695), .A2(n688), .ZN(n689) );
  NOR2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U760 ( .A(G1981), .B(G305), .Z(n960) );
  NAND2_X1 U761 ( .A1(n691), .A2(n960), .ZN(n698) );
  NOR2_X1 U762 ( .A1(G2090), .A2(G303), .ZN(n692) );
  NAND2_X1 U763 ( .A1(G8), .A2(n692), .ZN(n694) );
  NAND2_X1 U764 ( .A1(n694), .A2(n693), .ZN(n696) );
  NAND2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n729) );
  NOR2_X1 U767 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U768 ( .A(n705), .B(KEYINPUT90), .ZN(n751) );
  NAND2_X1 U769 ( .A1(G105), .A2(n884), .ZN(n706) );
  XNOR2_X1 U770 ( .A(n706), .B(KEYINPUT38), .ZN(n714) );
  NAND2_X1 U771 ( .A1(G141), .A2(n883), .ZN(n709) );
  NAND2_X1 U772 ( .A1(G129), .A2(n707), .ZN(n708) );
  NAND2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U774 ( .A1(n887), .A2(G117), .ZN(n710) );
  XOR2_X1 U775 ( .A(KEYINPUT94), .B(n710), .Z(n711) );
  NOR2_X1 U776 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U777 ( .A1(n714), .A2(n713), .ZN(n871) );
  NAND2_X1 U778 ( .A1(G1996), .A2(n871), .ZN(n715) );
  XOR2_X1 U779 ( .A(KEYINPUT95), .B(n715), .Z(n725) );
  NAND2_X1 U780 ( .A1(G107), .A2(n887), .ZN(n717) );
  NAND2_X1 U781 ( .A1(G119), .A2(n707), .ZN(n716) );
  NAND2_X1 U782 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U783 ( .A(KEYINPUT92), .B(n718), .ZN(n721) );
  NAND2_X1 U784 ( .A1(G95), .A2(n884), .ZN(n719) );
  XNOR2_X1 U785 ( .A(KEYINPUT93), .B(n719), .ZN(n720) );
  NOR2_X1 U786 ( .A1(n721), .A2(n720), .ZN(n723) );
  NAND2_X1 U787 ( .A1(n883), .A2(G131), .ZN(n722) );
  NAND2_X1 U788 ( .A1(n723), .A2(n722), .ZN(n896) );
  NAND2_X1 U789 ( .A1(G1991), .A2(n896), .ZN(n724) );
  NAND2_X1 U790 ( .A1(n725), .A2(n724), .ZN(n1006) );
  AND2_X1 U791 ( .A1(n751), .A2(n1006), .ZN(n744) );
  XOR2_X1 U792 ( .A(n744), .B(KEYINPUT96), .Z(n727) );
  XNOR2_X1 U793 ( .A(G1986), .B(G290), .ZN(n947) );
  NAND2_X1 U794 ( .A1(n751), .A2(n947), .ZN(n726) );
  NAND2_X1 U795 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U796 ( .A1(n729), .A2(n728), .ZN(n740) );
  XNOR2_X1 U797 ( .A(KEYINPUT37), .B(G2067), .ZN(n749) );
  NAND2_X1 U798 ( .A1(G140), .A2(n883), .ZN(n731) );
  NAND2_X1 U799 ( .A1(G104), .A2(n884), .ZN(n730) );
  NAND2_X1 U800 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U801 ( .A(KEYINPUT34), .B(n732), .ZN(n738) );
  NAND2_X1 U802 ( .A1(G116), .A2(n887), .ZN(n734) );
  NAND2_X1 U803 ( .A1(G128), .A2(n707), .ZN(n733) );
  NAND2_X1 U804 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U805 ( .A(KEYINPUT91), .B(n735), .ZN(n736) );
  XNOR2_X1 U806 ( .A(KEYINPUT35), .B(n736), .ZN(n737) );
  NOR2_X1 U807 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U808 ( .A(KEYINPUT36), .B(n739), .ZN(n903) );
  NOR2_X1 U809 ( .A1(n749), .A2(n903), .ZN(n1010) );
  NAND2_X1 U810 ( .A1(n1010), .A2(n751), .ZN(n747) );
  NAND2_X1 U811 ( .A1(n740), .A2(n747), .ZN(n741) );
  XNOR2_X1 U812 ( .A(n741), .B(KEYINPUT106), .ZN(n754) );
  NOR2_X1 U813 ( .A1(G1996), .A2(n871), .ZN(n999) );
  NOR2_X1 U814 ( .A1(G1991), .A2(n896), .ZN(n1002) );
  NOR2_X1 U815 ( .A1(G1986), .A2(G290), .ZN(n742) );
  NOR2_X1 U816 ( .A1(n1002), .A2(n742), .ZN(n743) );
  NOR2_X1 U817 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U818 ( .A1(n999), .A2(n745), .ZN(n746) );
  XNOR2_X1 U819 ( .A(n746), .B(KEYINPUT39), .ZN(n748) );
  NAND2_X1 U820 ( .A1(n748), .A2(n747), .ZN(n750) );
  NAND2_X1 U821 ( .A1(n749), .A2(n903), .ZN(n1012) );
  NAND2_X1 U822 ( .A1(n750), .A2(n1012), .ZN(n752) );
  NAND2_X1 U823 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U824 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U825 ( .A(n755), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U826 ( .A(G2443), .B(G2446), .Z(n757) );
  XNOR2_X1 U827 ( .A(G2427), .B(G2451), .ZN(n756) );
  XNOR2_X1 U828 ( .A(n757), .B(n756), .ZN(n763) );
  XOR2_X1 U829 ( .A(G2430), .B(G2454), .Z(n759) );
  XNOR2_X1 U830 ( .A(G1341), .B(G1348), .ZN(n758) );
  XNOR2_X1 U831 ( .A(n759), .B(n758), .ZN(n761) );
  XOR2_X1 U832 ( .A(G2435), .B(G2438), .Z(n760) );
  XNOR2_X1 U833 ( .A(n761), .B(n760), .ZN(n762) );
  XOR2_X1 U834 ( .A(n763), .B(n762), .Z(n764) );
  AND2_X1 U835 ( .A1(G14), .A2(n764), .ZN(G401) );
  AND2_X1 U836 ( .A1(n767), .A2(n766), .ZN(G160) );
  AND2_X1 U837 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U838 ( .A(G120), .ZN(G236) );
  INV_X1 U839 ( .A(G69), .ZN(G235) );
  INV_X1 U840 ( .A(G108), .ZN(G238) );
  INV_X1 U841 ( .A(G132), .ZN(G219) );
  INV_X1 U842 ( .A(G82), .ZN(G220) );
  NAND2_X1 U843 ( .A1(G7), .A2(G661), .ZN(n768) );
  XNOR2_X1 U844 ( .A(n768), .B(KEYINPUT10), .ZN(n769) );
  XNOR2_X1 U845 ( .A(KEYINPUT72), .B(n769), .ZN(G223) );
  INV_X1 U846 ( .A(G223), .ZN(n839) );
  NAND2_X1 U847 ( .A1(n839), .A2(G567), .ZN(n770) );
  XNOR2_X1 U848 ( .A(n770), .B(KEYINPUT73), .ZN(n771) );
  XNOR2_X1 U849 ( .A(KEYINPUT11), .B(n771), .ZN(G234) );
  INV_X1 U850 ( .A(G860), .ZN(n779) );
  OR2_X1 U851 ( .A1(n956), .A2(n779), .ZN(G153) );
  NAND2_X1 U852 ( .A1(G868), .A2(G301), .ZN(n774) );
  INV_X1 U853 ( .A(G868), .ZN(n821) );
  NAND2_X1 U854 ( .A1(n948), .A2(n821), .ZN(n773) );
  NAND2_X1 U855 ( .A1(n774), .A2(n773), .ZN(G284) );
  XNOR2_X1 U856 ( .A(KEYINPUT76), .B(n821), .ZN(n775) );
  NOR2_X1 U857 ( .A1(G286), .A2(n775), .ZN(n776) );
  XOR2_X1 U858 ( .A(KEYINPUT77), .B(n776), .Z(n778) );
  NOR2_X1 U859 ( .A1(G868), .A2(G299), .ZN(n777) );
  NOR2_X1 U860 ( .A1(n778), .A2(n777), .ZN(G297) );
  NAND2_X1 U861 ( .A1(n779), .A2(G559), .ZN(n780) );
  INV_X1 U862 ( .A(n948), .ZN(n908) );
  NAND2_X1 U863 ( .A1(n780), .A2(n908), .ZN(n781) );
  XNOR2_X1 U864 ( .A(n781), .B(KEYINPUT78), .ZN(n782) );
  XNOR2_X1 U865 ( .A(KEYINPUT16), .B(n782), .ZN(G148) );
  NOR2_X1 U866 ( .A1(G868), .A2(n956), .ZN(n785) );
  NAND2_X1 U867 ( .A1(n908), .A2(G868), .ZN(n783) );
  NOR2_X1 U868 ( .A1(G559), .A2(n783), .ZN(n784) );
  NOR2_X1 U869 ( .A1(n785), .A2(n784), .ZN(G282) );
  NAND2_X1 U870 ( .A1(G135), .A2(n883), .ZN(n787) );
  NAND2_X1 U871 ( .A1(G111), .A2(n887), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U873 ( .A1(n707), .A2(G123), .ZN(n788) );
  XOR2_X1 U874 ( .A(KEYINPUT18), .B(n788), .Z(n789) );
  NOR2_X1 U875 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U876 ( .A1(n884), .A2(G99), .ZN(n791) );
  NAND2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n1003) );
  XNOR2_X1 U878 ( .A(G2096), .B(n1003), .ZN(n793) );
  NOR2_X1 U879 ( .A1(n793), .A2(G2100), .ZN(n794) );
  XNOR2_X1 U880 ( .A(n794), .B(KEYINPUT79), .ZN(G156) );
  NAND2_X1 U881 ( .A1(n908), .A2(G559), .ZN(n817) );
  XNOR2_X1 U882 ( .A(n956), .B(n817), .ZN(n795) );
  NOR2_X1 U883 ( .A1(n795), .A2(G860), .ZN(n807) );
  NAND2_X1 U884 ( .A1(G67), .A2(n796), .ZN(n799) );
  NAND2_X1 U885 ( .A1(G55), .A2(n797), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U887 ( .A(KEYINPUT80), .B(n800), .Z(n806) );
  NAND2_X1 U888 ( .A1(n801), .A2(G80), .ZN(n804) );
  NAND2_X1 U889 ( .A1(G93), .A2(n802), .ZN(n803) );
  AND2_X1 U890 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U891 ( .A1(n806), .A2(n805), .ZN(n820) );
  XOR2_X1 U892 ( .A(n807), .B(n820), .Z(G145) );
  XOR2_X1 U893 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n809) );
  XOR2_X1 U894 ( .A(n820), .B(KEYINPUT85), .Z(n808) );
  XNOR2_X1 U895 ( .A(n809), .B(n808), .ZN(n813) );
  XNOR2_X1 U896 ( .A(n810), .B(G305), .ZN(n811) );
  XNOR2_X1 U897 ( .A(n811), .B(G288), .ZN(n812) );
  XNOR2_X1 U898 ( .A(n813), .B(n812), .ZN(n815) );
  XNOR2_X1 U899 ( .A(G290), .B(G166), .ZN(n814) );
  XNOR2_X1 U900 ( .A(n815), .B(n814), .ZN(n816) );
  XNOR2_X1 U901 ( .A(n816), .B(n956), .ZN(n907) );
  XNOR2_X1 U902 ( .A(KEYINPUT86), .B(n817), .ZN(n818) );
  XNOR2_X1 U903 ( .A(n907), .B(n818), .ZN(n819) );
  NAND2_X1 U904 ( .A1(n819), .A2(G868), .ZN(n823) );
  NAND2_X1 U905 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U906 ( .A1(n823), .A2(n822), .ZN(G295) );
  NAND2_X1 U907 ( .A1(G2078), .A2(G2084), .ZN(n824) );
  XOR2_X1 U908 ( .A(KEYINPUT20), .B(n824), .Z(n825) );
  NAND2_X1 U909 ( .A1(G2090), .A2(n825), .ZN(n826) );
  XNOR2_X1 U910 ( .A(KEYINPUT21), .B(n826), .ZN(n827) );
  NAND2_X1 U911 ( .A1(n827), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U912 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U913 ( .A1(G220), .A2(G219), .ZN(n828) );
  XOR2_X1 U914 ( .A(KEYINPUT22), .B(n828), .Z(n829) );
  NOR2_X1 U915 ( .A1(G218), .A2(n829), .ZN(n830) );
  NAND2_X1 U916 ( .A1(G96), .A2(n830), .ZN(n844) );
  NAND2_X1 U917 ( .A1(n844), .A2(G2106), .ZN(n836) );
  NOR2_X1 U918 ( .A1(G235), .A2(G236), .ZN(n831) );
  XNOR2_X1 U919 ( .A(n831), .B(KEYINPUT87), .ZN(n832) );
  NOR2_X1 U920 ( .A1(G238), .A2(n832), .ZN(n833) );
  NAND2_X1 U921 ( .A1(n833), .A2(G57), .ZN(n834) );
  XNOR2_X1 U922 ( .A(n834), .B(KEYINPUT88), .ZN(n843) );
  NAND2_X1 U923 ( .A1(n843), .A2(G567), .ZN(n835) );
  NAND2_X1 U924 ( .A1(n836), .A2(n835), .ZN(n846) );
  NAND2_X1 U925 ( .A1(G483), .A2(G661), .ZN(n837) );
  NOR2_X1 U926 ( .A1(n846), .A2(n837), .ZN(n842) );
  NAND2_X1 U927 ( .A1(n842), .A2(G36), .ZN(n838) );
  XOR2_X1 U928 ( .A(KEYINPUT89), .B(n838), .Z(G176) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n839), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U931 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U933 ( .A1(n842), .A2(n841), .ZN(G188) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  NOR2_X1 U936 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U937 ( .A(n845), .B(KEYINPUT107), .ZN(G261) );
  INV_X1 U938 ( .A(G261), .ZN(G325) );
  INV_X1 U939 ( .A(n846), .ZN(G319) );
  XOR2_X1 U940 ( .A(G2100), .B(G2096), .Z(n848) );
  XNOR2_X1 U941 ( .A(KEYINPUT42), .B(G2678), .ZN(n847) );
  XNOR2_X1 U942 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U943 ( .A(KEYINPUT43), .B(G2072), .Z(n850) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2090), .ZN(n849) );
  XNOR2_X1 U945 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U946 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2084), .ZN(n853) );
  XNOR2_X1 U948 ( .A(n854), .B(n853), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1966), .B(G1956), .Z(n856) );
  XNOR2_X1 U950 ( .A(G1981), .B(G1961), .ZN(n855) );
  XNOR2_X1 U951 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U952 ( .A(n857), .B(G2474), .Z(n859) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n858) );
  XNOR2_X1 U954 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U955 ( .A(KEYINPUT41), .B(G1976), .Z(n861) );
  XNOR2_X1 U956 ( .A(G1986), .B(G1971), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U958 ( .A(n863), .B(n862), .ZN(G229) );
  NAND2_X1 U959 ( .A1(G124), .A2(n707), .ZN(n864) );
  XNOR2_X1 U960 ( .A(n864), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U961 ( .A1(n887), .A2(G112), .ZN(n865) );
  NAND2_X1 U962 ( .A1(n866), .A2(n865), .ZN(n870) );
  NAND2_X1 U963 ( .A1(G136), .A2(n883), .ZN(n868) );
  NAND2_X1 U964 ( .A1(G100), .A2(n884), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U966 ( .A1(n870), .A2(n869), .ZN(G162) );
  XNOR2_X1 U967 ( .A(G162), .B(n871), .ZN(n872) );
  XNOR2_X1 U968 ( .A(n872), .B(n1003), .ZN(n882) );
  NAND2_X1 U969 ( .A1(G118), .A2(n887), .ZN(n874) );
  NAND2_X1 U970 ( .A1(G130), .A2(n707), .ZN(n873) );
  NAND2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n880) );
  NAND2_X1 U972 ( .A1(n884), .A2(G106), .ZN(n875) );
  XNOR2_X1 U973 ( .A(n875), .B(KEYINPUT108), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G142), .A2(n883), .ZN(n876) );
  NAND2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U976 ( .A(KEYINPUT45), .B(n878), .Z(n879) );
  NOR2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U978 ( .A(n882), .B(n881), .Z(n895) );
  NAND2_X1 U979 ( .A1(G139), .A2(n883), .ZN(n886) );
  NAND2_X1 U980 ( .A1(G103), .A2(n884), .ZN(n885) );
  NAND2_X1 U981 ( .A1(n886), .A2(n885), .ZN(n893) );
  NAND2_X1 U982 ( .A1(n887), .A2(G115), .ZN(n888) );
  XNOR2_X1 U983 ( .A(n888), .B(KEYINPUT110), .ZN(n890) );
  NAND2_X1 U984 ( .A1(G127), .A2(n707), .ZN(n889) );
  NAND2_X1 U985 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U986 ( .A(KEYINPUT47), .B(n891), .Z(n892) );
  NOR2_X1 U987 ( .A1(n893), .A2(n892), .ZN(n1014) );
  XNOR2_X1 U988 ( .A(G160), .B(n1014), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n905) );
  XNOR2_X1 U990 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n898) );
  XNOR2_X1 U991 ( .A(n896), .B(KEYINPUT46), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U993 ( .A(n899), .B(KEYINPUT109), .Z(n901) );
  XNOR2_X1 U994 ( .A(G164), .B(KEYINPUT111), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U996 ( .A(n903), .B(n902), .Z(n904) );
  XNOR2_X1 U997 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U998 ( .A1(G37), .A2(n906), .ZN(G395) );
  XOR2_X1 U999 ( .A(KEYINPUT113), .B(n907), .Z(n910) );
  XNOR2_X1 U1000 ( .A(G171), .B(n908), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1002 ( .A(G286), .B(n911), .Z(n912) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n912), .ZN(G397) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n913) );
  XNOR2_X1 U1006 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1007 ( .A1(G401), .A2(n915), .ZN(n916) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n916), .ZN(n917) );
  XNOR2_X1 U1009 ( .A(KEYINPUT115), .B(n917), .ZN(n919) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1011 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1014 ( .A(KEYINPUT54), .B(G34), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(n920), .B(KEYINPUT120), .ZN(n921) );
  XNOR2_X1 U1016 ( .A(G2084), .B(n921), .ZN(n939) );
  XNOR2_X1 U1017 ( .A(G2090), .B(G35), .ZN(n936) );
  XOR2_X1 U1018 ( .A(G1991), .B(G25), .Z(n922) );
  NAND2_X1 U1019 ( .A1(G28), .A2(n922), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(n923), .B(KEYINPUT117), .ZN(n928) );
  XNOR2_X1 U1021 ( .A(G1996), .B(G32), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(n924), .B(G27), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n933) );
  XNOR2_X1 U1025 ( .A(G2067), .B(G26), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(G2072), .B(G33), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1028 ( .A(KEYINPUT118), .B(n931), .Z(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(KEYINPUT53), .B(n934), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(KEYINPUT119), .B(n937), .ZN(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1034 ( .A(KEYINPUT55), .B(n940), .Z(n941) );
  NOR2_X1 U1035 ( .A1(G29), .A2(n941), .ZN(n969) );
  XNOR2_X1 U1036 ( .A(KEYINPUT56), .B(G16), .ZN(n966) );
  XOR2_X1 U1037 ( .A(G1971), .B(G166), .Z(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n955) );
  XNOR2_X1 U1041 ( .A(G299), .B(G1956), .ZN(n953) );
  XNOR2_X1 U1042 ( .A(G301), .B(G1961), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(n948), .B(G1348), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(KEYINPUT121), .B(n951), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n958) );
  XNOR2_X1 U1048 ( .A(G1341), .B(n956), .ZN(n957) );
  NOR2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(KEYINPUT122), .B(n959), .ZN(n964) );
  XNOR2_X1 U1051 ( .A(G168), .B(G1966), .ZN(n961) );
  NAND2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(KEYINPUT57), .B(n962), .ZN(n963) );
  NAND2_X1 U1054 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1055 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1056 ( .A1(n967), .A2(G11), .ZN(n968) );
  NOR2_X1 U1057 ( .A1(n969), .A2(n968), .ZN(n996) );
  XOR2_X1 U1058 ( .A(G1966), .B(G21), .Z(n981) );
  XNOR2_X1 U1059 ( .A(KEYINPUT123), .B(G1956), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(n970), .B(G20), .ZN(n976) );
  XOR2_X1 U1061 ( .A(G4), .B(KEYINPUT124), .Z(n972) );
  XNOR2_X1 U1062 ( .A(G1348), .B(KEYINPUT59), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(n972), .B(n971), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(G1341), .B(G19), .ZN(n973) );
  NOR2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(G6), .B(G1981), .ZN(n977) );
  NOR2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(n979), .B(KEYINPUT60), .ZN(n980) );
  NAND2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(KEYINPUT125), .B(n982), .ZN(n991) );
  XNOR2_X1 U1072 ( .A(G1961), .B(G5), .ZN(n989) );
  XNOR2_X1 U1073 ( .A(G1986), .B(G24), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(G1971), .B(G22), .ZN(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n986) );
  XOR2_X1 U1076 ( .A(G1976), .B(G23), .Z(n985) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(KEYINPUT58), .B(n987), .ZN(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(KEYINPUT61), .B(n992), .ZN(n993) );
  NOR2_X1 U1082 ( .A1(n993), .A2(G16), .ZN(n994) );
  XOR2_X1 U1083 ( .A(KEYINPUT126), .B(n994), .Z(n995) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(n997), .B(KEYINPUT127), .ZN(n1025) );
  XOR2_X1 U1086 ( .A(G2090), .B(G162), .Z(n998) );
  NOR2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1088 ( .A(KEYINPUT51), .B(n1000), .Z(n1008) );
  XOR2_X1 U1089 ( .A(G160), .B(G2084), .Z(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1094 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(n1011), .B(KEYINPUT116), .ZN(n1013) );
  NAND2_X1 U1096 ( .A1(n1013), .A2(n1012), .ZN(n1019) );
  XOR2_X1 U1097 ( .A(G2072), .B(n1014), .Z(n1016) );
  XOR2_X1 U1098 ( .A(G164), .B(G2078), .Z(n1015) );
  NOR2_X1 U1099 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1100 ( .A(KEYINPUT50), .B(n1017), .Z(n1018) );
  NOR2_X1 U1101 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1102 ( .A(KEYINPUT52), .B(n1020), .ZN(n1022) );
  INV_X1 U1103 ( .A(KEYINPUT55), .ZN(n1021) );
  NAND2_X1 U1104 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1105 ( .A1(n1023), .A2(G29), .ZN(n1024) );
  NAND2_X1 U1106 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

