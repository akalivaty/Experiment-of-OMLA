//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n638, new_n639, new_n640, new_n643, new_n644, new_n646, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  OR2_X1    g035(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(KEYINPUT67), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(G125), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n463), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n463), .A2(G137), .A3(new_n464), .ZN(new_n475));
  INV_X1    g050(.A(G101), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2104), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n475), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n474), .A2(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT70), .Z(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n461), .A2(new_n462), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(new_n464), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G124), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n483), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n469), .A2(new_n470), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT68), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n464), .A2(new_n493), .A3(new_n477), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(G136), .B2(new_n495), .ZN(new_n496));
  XOR2_X1   g071(.A(new_n496), .B(KEYINPUT71), .Z(G162));
  AND2_X1   g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n464), .A2(new_n498), .ZN(new_n499));
  OR2_X1    g074(.A1(KEYINPUT72), .A2(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT72), .A2(G114), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n477), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AND3_X1   g079(.A1(new_n461), .A2(G138), .A3(new_n462), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n466), .A2(new_n505), .A3(new_n506), .A4(new_n471), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n461), .A2(G138), .A3(new_n462), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT4), .B1(new_n491), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n504), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n510), .A2(KEYINPUT73), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  AOI211_X1 g087(.A(new_n512), .B(new_n504), .C1(new_n509), .C2(new_n507), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n511), .A2(new_n513), .ZN(G164));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT74), .B(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT75), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT74), .A2(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT74), .A2(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT6), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n524), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n518), .B1(new_n527), .B2(new_n529), .ZN(new_n531));
  AOI22_X1  g106(.A1(G50), .A2(new_n530), .B1(new_n531), .B2(G88), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n523), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(G166));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT76), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n531), .A2(G89), .ZN(new_n538));
  XNOR2_X1  g113(.A(KEYINPUT5), .B(G543), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n539), .A2(G63), .A3(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n530), .A2(G51), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n537), .A2(new_n538), .A3(new_n540), .A4(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n518), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(new_n521), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT6), .ZN(new_n548));
  OR2_X1    g123(.A1(KEYINPUT74), .A2(G651), .ZN(new_n549));
  NAND2_X1  g124(.A1(KEYINPUT74), .A2(G651), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g126(.A(G90), .B(new_n539), .C1(new_n551), .C2(new_n528), .ZN(new_n552));
  XOR2_X1   g127(.A(KEYINPUT77), .B(G52), .Z(new_n553));
  OAI211_X1 g128(.A(G543), .B(new_n553), .C1(new_n551), .C2(new_n528), .ZN(new_n554));
  AND3_X1   g129(.A1(new_n552), .A2(new_n554), .A3(KEYINPUT78), .ZN(new_n555));
  AOI21_X1  g130(.A(KEYINPUT78), .B1(new_n552), .B2(new_n554), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n547), .B1(new_n555), .B2(new_n556), .ZN(G301));
  INV_X1    g132(.A(G301), .ZN(G171));
  AOI22_X1  g133(.A1(new_n539), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  INV_X1    g134(.A(new_n521), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT79), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G56), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n518), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(new_n565), .A3(new_n521), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(G43), .A2(new_n530), .B1(new_n531), .B2(G81), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(G188));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT80), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G65), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n577), .B(new_n579), .C1(new_n516), .C2(new_n517), .ZN(new_n580));
  NAND2_X1  g155(.A1(G78), .A2(G543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(G91), .A2(new_n531), .B1(new_n582), .B2(G651), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n528), .B1(new_n521), .B2(KEYINPUT6), .ZN(new_n584));
  INV_X1    g159(.A(G53), .ZN(new_n585));
  NOR4_X1   g160(.A1(new_n584), .A2(KEYINPUT9), .A3(new_n585), .A4(new_n524), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT9), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n530), .B2(G53), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n583), .B1(new_n586), .B2(new_n588), .ZN(G299));
  XOR2_X1   g164(.A(new_n533), .B(KEYINPUT81), .Z(G303));
  NAND2_X1  g165(.A1(new_n530), .A2(G49), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n531), .A2(G87), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n539), .B2(G74), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT82), .Z(G288));
  NAND2_X1  g170(.A1(G73), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n518), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(new_n521), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n531), .A2(G86), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n530), .A2(G48), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(G305));
  NAND2_X1  g181(.A1(new_n531), .A2(G85), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n530), .A2(G47), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n539), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n607), .B(new_n608), .C1(new_n560), .C2(new_n609), .ZN(G290));
  OAI211_X1 g185(.A(G92), .B(new_n539), .C1(new_n551), .C2(new_n528), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT85), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n539), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G651), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(G54), .B1(new_n530), .B2(KEYINPUT84), .ZN(new_n618));
  OAI211_X1 g193(.A(KEYINPUT84), .B(G543), .C1(new_n551), .C2(new_n528), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n614), .B(new_n617), .C1(new_n618), .C2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n584), .B2(new_n524), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n624), .A2(G54), .A3(new_n619), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n614), .B1(new_n625), .B2(new_n617), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n613), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(KEYINPUT86), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n617), .B1(new_n618), .B2(new_n620), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT85), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(new_n621), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n629), .B1(new_n632), .B2(new_n613), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G868), .ZN(new_n635));
  MUX2_X1   g210(.A(G301), .B(new_n634), .S(new_n635), .Z(G321));
  XNOR2_X1  g211(.A(G321), .B(KEYINPUT87), .ZN(G284));
  OR3_X1    g212(.A1(G168), .A2(KEYINPUT88), .A3(new_n635), .ZN(new_n638));
  OAI21_X1  g213(.A(KEYINPUT88), .B1(G168), .B2(new_n635), .ZN(new_n639));
  INV_X1    g214(.A(G299), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n638), .B(new_n639), .C1(G868), .C2(new_n640), .ZN(G297));
  OAI211_X1 g216(.A(new_n638), .B(new_n639), .C1(G868), .C2(new_n640), .ZN(G280));
  NOR2_X1   g217(.A1(new_n634), .A2(G559), .ZN(new_n643));
  INV_X1    g218(.A(new_n634), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n643), .B1(G860), .B2(new_n644), .ZN(G148));
  NAND2_X1  g220(.A1(new_n569), .A2(new_n635), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n643), .B2(new_n635), .ZN(G323));
  XNOR2_X1  g222(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g223(.A1(new_n466), .A2(new_n471), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n649), .A2(new_n478), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT12), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT13), .ZN(new_n652));
  INV_X1    g227(.A(G2100), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  OAI221_X1 g230(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n463), .C2(G111), .ZN(new_n656));
  INV_X1    g231(.A(new_n495), .ZN(new_n657));
  INV_X1    g232(.A(G135), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(G123), .B2(new_n487), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2096), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n654), .A2(new_n655), .A3(new_n661), .ZN(G156));
  XOR2_X1   g237(.A(KEYINPUT15), .B(G2435), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2438), .ZN(new_n664));
  XOR2_X1   g239(.A(G2427), .B(G2430), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT90), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT89), .B(KEYINPUT14), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n664), .A2(new_n666), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2451), .B(G2454), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT16), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1341), .B(G1348), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n670), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2443), .B(G2446), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  AND3_X1   g253(.A1(new_n677), .A2(G14), .A3(new_n678), .ZN(G401));
  INV_X1    g254(.A(KEYINPUT18), .ZN(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(KEYINPUT17), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n680), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(new_n653), .ZN(new_n687));
  XOR2_X1   g262(.A(G2072), .B(G2078), .Z(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n683), .B2(KEYINPUT18), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(G2096), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n687), .B(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT92), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1971), .B(G1976), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT19), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1956), .B(G2474), .Z(new_n698));
  XOR2_X1   g273(.A(G1961), .B(G1966), .Z(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT91), .B(KEYINPUT20), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n698), .A2(new_n699), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(new_n705), .B(new_n704), .S(new_n697), .Z(new_n706));
  NOR2_X1   g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1981), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(G1986), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(G1986), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n694), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n709), .A2(new_n694), .A3(new_n710), .ZN(new_n713));
  XNOR2_X1  g288(.A(G1991), .B(G1996), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n714), .ZN(new_n717));
  AND3_X1   g292(.A1(new_n709), .A2(new_n694), .A3(new_n710), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(new_n711), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n716), .A2(new_n720), .ZN(G229));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G22), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G166), .B2(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G1971), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n722), .A2(G6), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n599), .B(KEYINPUT83), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n728), .A2(new_n604), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n727), .B1(new_n729), .B2(new_n722), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT32), .B(G1981), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n722), .A2(G23), .ZN(new_n733));
  INV_X1    g308(.A(new_n594), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(new_n722), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT33), .B(G1976), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n726), .A2(new_n732), .A3(new_n737), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(KEYINPUT34), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(KEYINPUT34), .ZN(new_n740));
  NOR2_X1   g315(.A1(G25), .A2(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n487), .A2(G119), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n495), .A2(G131), .ZN(new_n743));
  OAI221_X1 g318(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n463), .C2(G107), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT93), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n741), .B1(new_n747), .B2(G29), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT35), .B(G1991), .Z(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n748), .A2(new_n750), .ZN(new_n752));
  MUX2_X1   g327(.A(G24), .B(G290), .S(G16), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1986), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n739), .A2(new_n740), .A3(new_n751), .A4(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n757));
  OR3_X1    g332(.A1(new_n756), .A2(KEYINPUT94), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G4), .A2(G16), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n644), .B2(G16), .ZN(new_n760));
  INV_X1    g335(.A(G1348), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G33), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n495), .A2(G139), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT95), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT25), .Z(new_n768));
  AND2_X1   g343(.A1(new_n466), .A2(new_n471), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n769), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n768), .B1(new_n770), .B2(new_n463), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(new_n764), .B(new_n772), .S(G29), .Z(new_n773));
  INV_X1    g348(.A(G2072), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT98), .ZN(new_n776));
  INV_X1    g351(.A(G29), .ZN(new_n777));
  AND2_X1   g352(.A1(KEYINPUT24), .A2(G34), .ZN(new_n778));
  NOR2_X1   g353(.A1(KEYINPUT24), .A2(G34), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT96), .Z(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G160), .B2(G29), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT97), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G2084), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n777), .A2(G32), .ZN(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT26), .Z(new_n787));
  INV_X1    g362(.A(G105), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n478), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n487), .B2(G129), .ZN(new_n790));
  INV_X1    g365(.A(G141), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n657), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n785), .B1(new_n793), .B2(new_n777), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT27), .B(G1996), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n773), .A2(new_n774), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n776), .A2(new_n784), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT99), .ZN(new_n799));
  NOR2_X1   g374(.A1(G29), .A2(G35), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G162), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT29), .ZN(new_n802));
  INV_X1    g377(.A(G2090), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G168), .A2(new_n722), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n722), .B2(G21), .ZN(new_n806));
  INV_X1    g381(.A(G1966), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT100), .ZN(new_n809));
  NOR2_X1   g384(.A1(G5), .A2(G16), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G171), .B2(G16), .ZN(new_n811));
  INV_X1    g386(.A(G1961), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n809), .B(new_n813), .C1(G2084), .C2(new_n783), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n660), .A2(G29), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT31), .B(G11), .Z(new_n816));
  INV_X1    g391(.A(KEYINPUT30), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n777), .B1(new_n817), .B2(G28), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(KEYINPUT101), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n819), .A2(KEYINPUT101), .B1(new_n817), .B2(G28), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n816), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n815), .B(new_n822), .C1(new_n795), .C2(new_n796), .ZN(new_n823));
  NOR2_X1   g398(.A1(G27), .A2(G29), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G164), .B2(G29), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n825), .A2(G2078), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n777), .A2(G26), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT28), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n487), .A2(G128), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n831));
  INV_X1    g406(.A(G116), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n831), .B1(new_n484), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n495), .B2(G140), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n829), .B1(new_n835), .B2(G29), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G2067), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n827), .B(new_n837), .C1(G2078), .C2(new_n825), .ZN(new_n838));
  NOR2_X1   g413(.A1(G16), .A2(G19), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n570), .B2(G16), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(G1341), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n722), .A2(G20), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT23), .Z(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(G299), .B2(G16), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G1956), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n806), .A2(new_n807), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n841), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n814), .A2(new_n838), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n799), .A2(new_n804), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT94), .B(KEYINPUT36), .ZN(new_n850));
  AOI211_X1 g425(.A(new_n763), .B(new_n849), .C1(new_n756), .C2(new_n850), .ZN(G311));
  AOI21_X1  g426(.A(new_n849), .B1(new_n756), .B2(new_n850), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n852), .A2(new_n758), .A3(new_n762), .ZN(G150));
  NAND2_X1  g428(.A1(new_n644), .A2(G559), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n531), .A2(G93), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  INV_X1    g432(.A(G67), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n857), .B1(new_n518), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g434(.A1(new_n530), .A2(G55), .B1(new_n859), .B2(new_n521), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n567), .A2(new_n568), .A3(new_n856), .A4(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n567), .A2(new_n568), .B1(new_n860), .B2(new_n856), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n855), .B(new_n864), .Z(new_n865));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n866));
  AOI21_X1  g441(.A(G860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n866), .B2(new_n865), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n860), .A2(new_n856), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G860), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(G145));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n660), .B(G160), .Z(new_n874));
  XNOR2_X1  g449(.A(G162), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n507), .A2(new_n509), .ZN(new_n876));
  INV_X1    g451(.A(new_n504), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n835), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n792), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n772), .ZN(new_n881));
  OAI21_X1  g456(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n882));
  INV_X1    g457(.A(G118), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n484), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n487), .B2(G130), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n495), .A2(KEYINPUT102), .A3(G142), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT102), .B1(new_n495), .B2(G142), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(new_n651), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n746), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n875), .B1(new_n881), .B2(new_n891), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n880), .A2(new_n772), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n880), .A2(new_n772), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n873), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n881), .A2(new_n897), .A3(new_n891), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n893), .B(new_n894), .C1(KEYINPUT103), .C2(new_n890), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n875), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g477(.A(new_n643), .B(new_n864), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n640), .B1(new_n632), .B2(new_n613), .ZN(new_n905));
  AOI211_X1 g480(.A(G299), .B(new_n612), .C1(new_n631), .C2(new_n621), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n627), .A2(G299), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n632), .A2(new_n640), .A3(new_n613), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(KEYINPUT41), .A3(new_n909), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n729), .B(KEYINPUT104), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(G166), .ZN(new_n916));
  XNOR2_X1  g491(.A(G290), .B(new_n594), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(G305), .B(KEYINPUT104), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n533), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n916), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n916), .A2(new_n921), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n917), .B(new_n918), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT42), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n914), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n912), .A3(new_n913), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n635), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n869), .A2(new_n635), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  OR3_X1    g507(.A1(new_n930), .A2(KEYINPUT106), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT106), .B1(new_n930), .B2(new_n932), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(G295));
  OR3_X1    g510(.A1(new_n930), .A2(KEYINPUT107), .A3(new_n932), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT107), .B1(new_n930), .B2(new_n932), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(G331));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  OAI21_X1  g514(.A(G171), .B1(new_n862), .B2(new_n863), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n569), .A2(new_n869), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n941), .A2(new_n861), .A3(G301), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(G168), .A3(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n941), .A2(new_n861), .A3(G301), .ZN(new_n944));
  AOI21_X1  g519(.A(G301), .B1(new_n941), .B2(new_n861), .ZN(new_n945));
  OAI21_X1  g520(.A(G286), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n907), .A2(new_n910), .A3(new_n943), .A4(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n905), .A2(new_n906), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n944), .A2(new_n945), .A3(G286), .ZN(new_n949));
  AOI21_X1  g524(.A(G168), .B1(new_n940), .B2(new_n942), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT108), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n924), .B1(new_n916), .B2(new_n921), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(new_n919), .B2(new_n923), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n947), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n953), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(G37), .B1(new_n925), .B2(new_n952), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n947), .A2(new_n956), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n956), .B1(new_n947), .B2(new_n951), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n925), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n958), .A2(new_n964), .A3(new_n965), .A4(new_n873), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n939), .B1(new_n961), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n958), .A2(new_n964), .A3(new_n873), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT109), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT43), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n968), .B2(KEYINPUT43), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n958), .A2(new_n959), .A3(new_n965), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n967), .B1(new_n974), .B2(new_n939), .ZN(G397));
  INV_X1    g550(.A(G40), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n474), .A2(new_n479), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n510), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n878), .A2(new_n512), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n510), .A2(KEYINPUT73), .ZN(new_n982));
  AOI21_X1  g557(.A(G1384), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT120), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n980), .B(KEYINPUT120), .C1(new_n983), .C2(new_n984), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n812), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n510), .A2(G1384), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n978), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(G2078), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n993), .B(new_n995), .C1(new_n990), .C2(new_n992), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n510), .A2(new_n990), .A3(G1384), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n978), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n983), .B2(KEYINPUT45), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n998), .B(KEYINPUT111), .C1(new_n983), .C2(KEYINPUT45), .ZN(new_n1002));
  AOI21_X1  g577(.A(G2078), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n989), .B(new_n996), .C1(new_n1003), .C2(KEYINPUT53), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(G171), .ZN(new_n1005));
  INV_X1    g580(.A(G2078), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1002), .ZN(new_n1007));
  INV_X1    g582(.A(G1384), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n511), .B2(new_n513), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n990), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT111), .B1(new_n1010), .B2(new_n998), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1006), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n994), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT118), .B1(new_n1009), .B2(new_n990), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n983), .A2(new_n1015), .A3(KEYINPUT45), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1014), .A2(new_n1016), .A3(new_n995), .A4(new_n993), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1013), .A2(G301), .A3(new_n1017), .A4(new_n989), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1005), .A2(KEYINPUT54), .A3(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT125), .B(KEYINPUT54), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1017), .B(new_n989), .C1(new_n1003), .C2(KEYINPUT53), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(G171), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1013), .A2(G301), .A3(new_n989), .A4(new_n996), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G286), .A2(G8), .ZN(new_n1026));
  XOR2_X1   g601(.A(new_n1026), .B(KEYINPUT124), .Z(new_n1027));
  NAND3_X1  g602(.A1(new_n1014), .A2(new_n1016), .A3(new_n993), .ZN(new_n1028));
  INV_X1    g603(.A(new_n985), .ZN(new_n1029));
  INV_X1    g604(.A(G2084), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1028), .A2(new_n807), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G8), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1025), .B(new_n1027), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1027), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1031), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1034), .B1(new_n1035), .B2(G8), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT51), .B1(new_n1031), .B2(new_n1027), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1033), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1019), .A2(new_n1024), .A3(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1040));
  XNOR2_X1  g615(.A(G299), .B(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1956), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n984), .B(new_n1008), .C1(new_n511), .C2(new_n513), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT50), .B1(new_n510), .B2(G1384), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(new_n977), .A3(KEYINPUT116), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT116), .B1(new_n1045), .B2(new_n977), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1043), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT56), .B(G2072), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1010), .A2(new_n998), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1042), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n987), .A2(new_n761), .A3(new_n988), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n977), .A2(new_n991), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G2067), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n634), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1049), .A2(new_n1042), .A3(new_n1051), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1052), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n644), .A2(KEYINPUT60), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT60), .B1(new_n628), .B2(new_n633), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1053), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1062), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n1067));
  INV_X1    g642(.A(G1996), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n998), .B(new_n1068), .C1(new_n983), .C2(KEYINPUT45), .ZN(new_n1069));
  XOR2_X1   g644(.A(KEYINPUT58), .B(G1341), .Z(new_n1070));
  NAND2_X1  g645(.A1(new_n1054), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n570), .ZN(new_n1073));
  NOR2_X1   g648(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1067), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n569), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1077), .A2(KEYINPUT122), .A3(new_n1074), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1066), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1041), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1081), .A2(KEYINPUT61), .A3(new_n1059), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1073), .A2(new_n1067), .A3(new_n1075), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT122), .B1(new_n1077), .B2(new_n1074), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1083), .A2(new_n1084), .A3(KEYINPUT121), .A4(KEYINPUT59), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1065), .A2(new_n1079), .A3(new_n1082), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1081), .A2(new_n1059), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT61), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT123), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1049), .A2(new_n1042), .A3(new_n1051), .ZN(new_n1090));
  OAI211_X1 g665(.A(KEYINPUT123), .B(new_n1088), .C1(new_n1090), .C2(new_n1052), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1060), .B1(new_n1086), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n605), .A2(new_n599), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G1981), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT114), .B(G1981), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1097), .B1(new_n729), .B2(new_n1098), .ZN(new_n1099));
  AND4_X1   g674(.A1(new_n1097), .A2(new_n601), .A3(new_n605), .A4(new_n1098), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT49), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1055), .A2(new_n1032), .ZN(new_n1104));
  OAI211_X1 g679(.A(KEYINPUT49), .B(new_n1096), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n734), .A2(G1976), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1054), .A2(G8), .A3(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1108), .A2(KEYINPUT52), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1108), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT113), .B(G1976), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT52), .B1(G288), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1109), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1106), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(G303), .A2(G8), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1115), .B(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1001), .A2(new_n725), .A3(new_n1002), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1029), .A2(new_n803), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1032), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1114), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n1123));
  OR3_X1    g698(.A1(new_n1047), .A2(G2090), .A3(new_n1048), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1119), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1123), .B1(new_n1119), .B2(new_n1124), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1125), .A2(new_n1126), .A3(new_n1032), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1122), .B1(new_n1127), .B2(new_n1118), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT126), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1130), .B(new_n1122), .C1(new_n1127), .C2(new_n1118), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1039), .A2(new_n1094), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(KEYINPUT62), .B(new_n1033), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1133), .A2(G171), .A3(new_n1021), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1038), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1134), .A2(new_n1129), .A3(new_n1131), .A4(new_n1136), .ZN(new_n1137));
  AOI211_X1 g712(.A(G1976), .B(G288), .C1(new_n1103), .C2(new_n1105), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1104), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n1141), .B2(new_n1114), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1035), .A2(G8), .A3(G168), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1122), .B(new_n1144), .C1(new_n1127), .C2(new_n1118), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1148), .B(new_n1122), .C1(new_n1121), .C2(new_n1118), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1142), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1132), .A2(new_n1137), .A3(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(G290), .A2(G1986), .ZN(new_n1152));
  NOR2_X1   g727(.A1(G290), .A2(G1986), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1152), .A2(new_n1153), .A3(KEYINPUT110), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n978), .A2(KEYINPUT45), .A3(new_n991), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  AOI211_X1 g731(.A(new_n1154), .B(new_n1156), .C1(KEYINPUT110), .C2(new_n1152), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n792), .B(new_n1068), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n835), .B(new_n1056), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1160), .B1(new_n746), .B2(new_n750), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n747), .A2(new_n749), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1157), .B1(new_n1163), .B2(new_n1155), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1151), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(new_n1155), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1155), .A2(new_n1153), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT48), .ZN(new_n1168));
  OAI22_X1  g743(.A1(new_n1162), .A2(new_n1160), .B1(G2067), .B2(new_n835), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1166), .A2(new_n1168), .B1(new_n1155), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1156), .B1(new_n1159), .B2(new_n793), .ZN(new_n1171));
  OR3_X1    g746(.A1(new_n1156), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1172));
  OAI21_X1  g747(.A(KEYINPUT46), .B1(new_n1156), .B2(G1996), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT47), .Z(new_n1175));
  AND2_X1   g750(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1165), .A2(new_n1176), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g752(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1179));
  INV_X1    g753(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g754(.A(new_n1180), .B1(new_n715), .B2(new_n719), .ZN(new_n1181));
  OAI21_X1  g755(.A(new_n1181), .B1(new_n896), .B2(new_n900), .ZN(new_n1182));
  NAND2_X1  g756(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n1183));
  AOI21_X1  g757(.A(new_n973), .B1(new_n1183), .B2(KEYINPUT109), .ZN(new_n1184));
  NAND3_X1  g758(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT43), .ZN(new_n1185));
  AOI211_X1 g759(.A(KEYINPUT127), .B(new_n1182), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n1183), .A2(KEYINPUT109), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n1188), .A2(new_n1185), .A3(new_n972), .ZN(new_n1189));
  INV_X1    g763(.A(new_n1182), .ZN(new_n1190));
  AOI21_X1  g764(.A(new_n1187), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g765(.A1(new_n1186), .A2(new_n1191), .ZN(G308));
  OAI21_X1  g766(.A(KEYINPUT127), .B1(new_n974), .B2(new_n1182), .ZN(new_n1193));
  NAND3_X1  g767(.A1(new_n1189), .A2(new_n1187), .A3(new_n1190), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n1193), .A2(new_n1194), .ZN(G225));
endmodule


