//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n566, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n592, new_n594, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n644,
    new_n645, new_n648, new_n649, new_n651, new_n652, new_n653, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G235), .A2(G236), .A3(G237), .A4(G238), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT68), .Z(new_n453));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT69), .Z(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n467), .A2(G2105), .B1(G137), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT71), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT70), .B1(new_n469), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(new_n477), .A3(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G101), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n474), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n475), .A2(new_n478), .A3(KEYINPUT71), .A4(G101), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n473), .A2(new_n483), .ZN(G160));
  NOR2_X1   g059(.A1(new_n465), .A2(new_n477), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  AND2_X1   g061(.A1(G112), .A2(G2105), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(G100), .B2(new_n477), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n469), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(G136), .B2(new_n472), .ZN(G162));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n470), .B2(new_n471), .ZN(new_n492));
  AND2_X1   g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  OAI21_X1  g068(.A(G2105), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n477), .C1(new_n463), .C2(new_n464), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n470), .A2(new_n471), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT4), .A2(G138), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n498), .A2(new_n500), .B1(G102), .B2(G2104), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n494), .B(new_n497), .C1(G2105), .C2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT5), .B1(new_n507), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT5), .A4(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(G88), .B1(G50), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n518), .B1(KEYINPUT72), .B2(new_n514), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n514), .A2(KEYINPUT73), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n512), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(G62), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n521), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(KEYINPUT74), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n517), .B1(new_n529), .B2(G651), .ZN(G166));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n531));
  OAI211_X1 g106(.A(G51), .B(G543), .C1(new_n504), .C2(new_n505), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n531), .B(new_n532), .C1(new_n526), .C2(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n533), .B1(new_n511), .B2(new_n512), .ZN(new_n535));
  INV_X1    g110(.A(new_n532), .ZN(new_n536));
  OAI21_X1  g111(.A(KEYINPUT75), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n504), .A2(new_n505), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n521), .A2(G89), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n534), .A2(new_n537), .A3(new_n539), .A4(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  INV_X1    g118(.A(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n521), .A2(G64), .ZN(new_n545));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n521), .A2(G90), .A3(new_n538), .ZN(new_n548));
  XOR2_X1   g123(.A(KEYINPUT76), .B(G52), .Z(new_n549));
  NAND2_X1  g124(.A1(new_n515), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n547), .A2(new_n551), .ZN(G171));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(new_n521), .B2(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n553), .B1(new_n556), .B2(new_n544), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n511), .B2(new_n512), .ZN(new_n559));
  OAI211_X1 g134(.A(KEYINPUT77), .B(G651), .C1(new_n559), .C2(new_n555), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n513), .A2(G81), .B1(G43), .B2(new_n515), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(G188));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n511), .B2(new_n512), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT78), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n514), .A2(KEYINPUT72), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(KEYINPUT5), .B1(new_n509), .B2(G543), .ZN(new_n577));
  AND4_X1   g152(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT5), .A4(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(G65), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n579), .A2(new_n580), .A3(new_n573), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n575), .A2(new_n581), .A3(G651), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n538), .A2(G53), .A3(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT9), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT9), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n515), .A2(new_n586), .A3(G53), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n585), .A2(new_n587), .B1(new_n513), .B2(G91), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n582), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n583), .B1(new_n582), .B2(new_n588), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(G299));
  AOI22_X1  g166(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n548), .B(new_n550), .C1(new_n592), .C2(new_n544), .ZN(G301));
  AND2_X1   g168(.A1(new_n525), .A2(new_n528), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n516), .B1(new_n594), .B2(new_n544), .ZN(G303));
  NAND2_X1  g170(.A1(new_n521), .A2(new_n538), .ZN(new_n596));
  INV_X1    g171(.A(G87), .ZN(new_n597));
  OAI21_X1  g172(.A(KEYINPUT80), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n513), .A2(new_n599), .A3(G87), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n602), .A2(new_n603), .B1(new_n515), .B2(G49), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n601), .A2(new_n604), .A3(new_n605), .ZN(G288));
  AND2_X1   g181(.A1(G73), .A2(G543), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(new_n521), .B2(G61), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT82), .B1(new_n608), .B2(new_n544), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n521), .A2(G86), .A3(new_n538), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT83), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n610), .A2(new_n611), .B1(new_n515), .B2(G48), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n513), .A2(KEYINPUT83), .A3(G86), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n614));
  INV_X1    g189(.A(G61), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n511), .B2(new_n512), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n614), .B(G651), .C1(new_n616), .C2(new_n607), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n609), .A2(new_n612), .A3(new_n613), .A4(new_n617), .ZN(G305));
  AOI22_X1  g193(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n619), .A2(new_n544), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n515), .A2(G47), .ZN(new_n623));
  INV_X1    g198(.A(G85), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n596), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(G290));
  XOR2_X1   g202(.A(KEYINPUT87), .B(G66), .Z(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n512), .B2(new_n511), .ZN(new_n629));
  AND2_X1   g204(.A1(G79), .A2(G543), .ZN(new_n630));
  OAI21_X1  g205(.A(G651), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(new_n538), .B2(G543), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n632), .B(G543), .C1(new_n504), .C2(new_n505), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(G54), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT85), .B(KEYINPUT10), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n513), .B2(G92), .ZN(new_n638));
  AND4_X1   g213(.A1(G92), .A2(new_n521), .A3(new_n538), .A4(new_n637), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n631), .B(new_n636), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n640), .A2(G868), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g217(.A(new_n641), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g218(.A1(G286), .A2(G868), .ZN(new_n644));
  XOR2_X1   g219(.A(G299), .B(KEYINPUT88), .Z(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n645), .B2(G868), .ZN(G297));
  OAI21_X1  g221(.A(new_n644), .B1(new_n645), .B2(G868), .ZN(G280));
  INV_X1    g222(.A(new_n640), .ZN(new_n648));
  INV_X1    g223(.A(G559), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n649), .B2(G860), .ZN(G148));
  NOR2_X1   g225(.A1(new_n563), .A2(G868), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n640), .A2(G559), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n651), .B1(G868), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT89), .ZN(G323));
  XNOR2_X1  g229(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g230(.A(new_n479), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(new_n498), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT12), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT13), .ZN(new_n659));
  INV_X1    g234(.A(G2100), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  MUX2_X1   g237(.A(G99), .B(G111), .S(G2105), .Z(new_n663));
  AOI22_X1  g238(.A1(new_n485), .A2(G123), .B1(G2104), .B2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(G135), .ZN(new_n665));
  INV_X1    g240(.A(new_n472), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(G2096), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n661), .A2(new_n662), .A3(new_n669), .ZN(G156));
  XNOR2_X1  g245(.A(G2427), .B(G2430), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT92), .Z(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT15), .B(G2435), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT91), .B(G2438), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT90), .B(KEYINPUT14), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT93), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(KEYINPUT93), .B1(new_n676), .B2(new_n677), .ZN(new_n681));
  OAI22_X1  g256(.A1(new_n680), .A2(new_n681), .B1(new_n672), .B2(new_n675), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2451), .B(G2454), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT16), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2443), .B(G2446), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1341), .B(G1348), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g264(.A(G14), .B1(new_n687), .B2(new_n688), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(G401));
  XOR2_X1   g266(.A(G2084), .B(G2090), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G2072), .B(G2078), .Z(new_n694));
  XNOR2_X1  g269(.A(G2067), .B(G2678), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT18), .ZN(new_n698));
  INV_X1    g273(.A(new_n694), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n699), .A2(KEYINPUT17), .A3(new_n692), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n692), .B1(new_n699), .B2(KEYINPUT17), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n696), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n693), .A2(new_n696), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n699), .B1(new_n703), .B2(KEYINPUT17), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n698), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(new_n668), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G2100), .ZN(G227));
  XOR2_X1   g282(.A(G1971), .B(G1976), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT19), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1956), .B(G2474), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(G1961), .B(G1966), .Z(new_n712));
  AND2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT20), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n711), .A2(new_n712), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n709), .A2(new_n713), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n709), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(G1991), .B(G1996), .ZN(new_n722));
  XNOR2_X1  g297(.A(G1981), .B(G1986), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n721), .B(new_n724), .ZN(G229));
  OR2_X1    g300(.A1(G6), .A2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(G305), .B2(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT96), .Z(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT32), .B(G1981), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT97), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(new_n731), .ZN(new_n733));
  NOR2_X1   g308(.A1(G16), .A2(G22), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G166), .B2(G16), .ZN(new_n735));
  INV_X1    g310(.A(G1971), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n732), .A2(new_n733), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G16), .A2(G23), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT98), .ZN(new_n740));
  NAND2_X1  g315(.A1(G288), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT98), .A4(new_n605), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n739), .B1(new_n744), .B2(G16), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT33), .B(G1976), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  OR3_X1    g322(.A1(new_n738), .A2(KEYINPUT34), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(KEYINPUT34), .B1(new_n738), .B2(new_n747), .ZN(new_n749));
  NOR2_X1   g324(.A1(G25), .A2(G29), .ZN(new_n750));
  MUX2_X1   g325(.A(G95), .B(G107), .S(G2105), .Z(new_n751));
  AOI22_X1  g326(.A1(new_n485), .A2(G119), .B1(G2104), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n472), .A2(G131), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(KEYINPUT94), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(KEYINPUT94), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n750), .B1(new_n758), .B2(G29), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT35), .B(G1991), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n727), .A2(G24), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT95), .Z(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n626), .B2(new_n727), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(G1986), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(G1986), .ZN(new_n766));
  AND3_X1   g341(.A1(new_n761), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n748), .A2(new_n749), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT36), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT31), .B(G11), .Z(new_n770));
  INV_X1    g345(.A(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT30), .B(G28), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n485), .A2(G129), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n656), .A2(G105), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT26), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n472), .A2(G141), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n774), .A2(new_n775), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(new_n771), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n771), .B2(G32), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT27), .B(G1996), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n773), .B1(new_n771), .B2(new_n667), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G2084), .ZN(new_n785));
  NAND2_X1  g360(.A1(G160), .A2(G29), .ZN(new_n786));
  AND2_X1   g361(.A1(KEYINPUT24), .A2(G34), .ZN(new_n787));
  NOR2_X1   g362(.A1(KEYINPUT24), .A2(G34), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n771), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n784), .B1(new_n785), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G29), .A2(G35), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G162), .B2(G29), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT29), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n791), .B1(G2090), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(G2090), .ZN(new_n796));
  INV_X1    g371(.A(G1961), .ZN(new_n797));
  NOR2_X1   g372(.A1(G171), .A2(new_n727), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G5), .B2(new_n727), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n799), .A2(new_n797), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n782), .A2(new_n783), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT103), .ZN(new_n804));
  INV_X1    g379(.A(G2072), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT100), .B(KEYINPUT25), .Z(new_n806));
  NAND3_X1  g381(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n472), .A2(G139), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n498), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n808), .B(new_n809), .C1(new_n477), .C2(new_n810), .ZN(new_n811));
  MUX2_X1   g386(.A(G33), .B(new_n811), .S(G29), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT101), .ZN(new_n813));
  AOI211_X1 g388(.A(new_n802), .B(new_n804), .C1(new_n805), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n648), .A2(G16), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G4), .B2(G16), .ZN(new_n816));
  INV_X1    g391(.A(G1348), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n771), .A2(G26), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT28), .Z(new_n820));
  MUX2_X1   g395(.A(G104), .B(G116), .S(G2105), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G2104), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT99), .Z(new_n823));
  AOI22_X1  g398(.A1(new_n485), .A2(G128), .B1(G140), .B2(new_n472), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n820), .B1(new_n825), .B2(G29), .ZN(new_n826));
  INV_X1    g401(.A(G2067), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(G27), .A2(G29), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G164), .B2(G29), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G2078), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n790), .A2(new_n785), .ZN(new_n832));
  NOR4_X1   g407(.A1(new_n818), .A2(new_n828), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n813), .A2(new_n805), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT102), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n801), .A2(new_n814), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(G299), .A2(G16), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n727), .A2(G20), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT23), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G1956), .ZN(new_n841));
  NOR2_X1   g416(.A1(G16), .A2(G19), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n564), .B2(G16), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G1341), .ZN(new_n844));
  NOR2_X1   g419(.A1(G168), .A2(new_n727), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n727), .B2(G21), .ZN(new_n846));
  INV_X1    g421(.A(G1966), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n846), .A2(new_n847), .B1(new_n816), .B2(new_n817), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  NOR4_X1   g424(.A1(new_n836), .A2(new_n841), .A3(new_n844), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n769), .A2(new_n850), .ZN(G150));
  INV_X1    g426(.A(G150), .ZN(G311));
  NAND2_X1  g427(.A1(new_n515), .A2(G55), .ZN(new_n853));
  INV_X1    g428(.A(G93), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n596), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n521), .A2(G67), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n544), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n561), .A2(new_n859), .A3(new_n562), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n859), .B1(new_n561), .B2(new_n562), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT38), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n640), .A2(new_n649), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n866));
  AOI21_X1  g441(.A(G860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n866), .B2(new_n865), .ZN(new_n868));
  INV_X1    g443(.A(new_n859), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G860), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(G145));
  XNOR2_X1  g447(.A(new_n757), .B(new_n658), .ZN(new_n873));
  MUX2_X1   g448(.A(G106), .B(G118), .S(G2105), .Z(new_n874));
  AOI22_X1  g449(.A1(new_n485), .A2(G130), .B1(G2104), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G142), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(new_n666), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n873), .B(new_n877), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n825), .B(G164), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n873), .B(new_n877), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n879), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n811), .A2(KEYINPUT104), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n779), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n881), .A2(new_n886), .A3(new_n883), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(G162), .B(G160), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n667), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n888), .A2(new_n892), .A3(new_n889), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(G395));
  NOR2_X1   g474(.A1(new_n869), .A2(G868), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n744), .A2(new_n626), .ZN(new_n901));
  NAND2_X1  g476(.A1(G290), .A2(new_n743), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G166), .B(G305), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n908), .A2(KEYINPUT42), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT108), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(KEYINPUT42), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT107), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n862), .B(new_n652), .Z(new_n914));
  OAI21_X1  g489(.A(new_n648), .B1(new_n589), .B2(new_n590), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n582), .A2(new_n588), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT79), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n582), .A2(new_n583), .A3(new_n588), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n640), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n915), .A2(new_n919), .A3(KEYINPUT41), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT41), .B1(new_n915), .B2(new_n919), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n914), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT106), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n915), .A2(new_n919), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n914), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n923), .A2(KEYINPUT106), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n913), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n910), .A2(new_n912), .A3(new_n928), .A4(new_n927), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n900), .B1(new_n932), .B2(G868), .ZN(G295));
  AOI21_X1  g508(.A(new_n900), .B1(new_n932), .B2(G868), .ZN(G331));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT41), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n589), .A2(new_n590), .A3(new_n648), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n640), .B1(new_n917), .B2(new_n918), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n563), .A2(new_n869), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n561), .A2(new_n859), .A3(new_n562), .ZN(new_n941));
  NAND2_X1  g516(.A1(G286), .A2(G301), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n535), .A2(KEYINPUT75), .A3(new_n536), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n539), .A2(new_n541), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(G171), .A2(new_n945), .A3(new_n537), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n940), .A2(new_n941), .A3(new_n942), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n942), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n860), .B2(new_n861), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n915), .A2(new_n919), .A3(KEYINPUT41), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n939), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT109), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n939), .A2(new_n950), .A3(new_n954), .A4(new_n951), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT110), .B1(new_n950), .B2(new_n925), .ZN(new_n956));
  INV_X1    g531(.A(new_n925), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n957), .A2(new_n958), .A3(new_n949), .A4(new_n947), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n953), .A2(new_n955), .A3(new_n956), .A4(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n908), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n895), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n952), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n939), .A2(new_n950), .A3(KEYINPUT111), .A4(new_n951), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n957), .A2(new_n949), .A3(new_n947), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n908), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n935), .B1(new_n962), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n960), .A2(new_n961), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n959), .A2(new_n956), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n971), .A2(new_n908), .A3(new_n955), .A4(new_n953), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n970), .A2(new_n972), .A3(KEYINPUT43), .A4(new_n895), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT44), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n962), .B2(new_n968), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT111), .B1(new_n922), .B2(new_n950), .ZN(new_n977));
  INV_X1    g552(.A(new_n965), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n967), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n961), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n980), .A2(KEYINPUT112), .A3(new_n895), .A4(new_n972), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n976), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n970), .A2(new_n972), .A3(new_n935), .A4(new_n895), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n974), .B1(new_n985), .B2(KEYINPUT44), .ZN(G397));
  XOR2_X1   g561(.A(new_n757), .B(new_n760), .Z(new_n987));
  XNOR2_X1  g562(.A(new_n825), .B(new_n827), .ZN(new_n988));
  INV_X1    g563(.A(G1996), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n779), .B(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g567(.A1(G290), .A2(G1986), .ZN(new_n993));
  NAND2_X1  g568(.A1(G290), .A2(G1986), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT113), .B(KEYINPUT45), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n502), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n473), .A2(new_n483), .A3(G40), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n995), .A2(new_n1002), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n473), .A2(G40), .A3(new_n483), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n502), .A2(KEYINPUT50), .A3(new_n998), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT50), .B1(new_n502), .B2(new_n998), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1956), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n999), .A2(new_n1001), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n998), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT56), .B(G2072), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n916), .A2(KEYINPUT57), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n582), .A2(new_n1016), .A3(new_n588), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(new_n640), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT118), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1007), .A2(new_n817), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n502), .A2(new_n998), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1023), .A2(new_n1001), .A3(G2067), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1021), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  AOI211_X1 g601(.A(KEYINPUT118), .B(new_n1024), .C1(new_n1007), .C2(new_n817), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1015), .A2(KEYINPUT119), .A3(new_n1017), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT119), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1020), .A2(new_n1028), .B1(new_n1014), .B2(new_n1031), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1026), .A2(new_n1027), .A3(KEYINPUT60), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT60), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n648), .ZN(new_n1035));
  OAI211_X1 g610(.A(KEYINPUT60), .B(new_n640), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT122), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1014), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1018), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT122), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1040), .A2(new_n1009), .A3(new_n1041), .A4(new_n1013), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1038), .A2(new_n1039), .A3(KEYINPUT61), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT61), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1040), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1044), .B1(new_n1019), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G102), .A2(G2104), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n465), .B2(new_n499), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1048), .A2(new_n477), .B1(new_n496), .B2(new_n495), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1384), .B1(new_n1049), .B2(new_n494), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1004), .B(new_n1011), .C1(new_n1050), .C2(new_n997), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1023), .A2(new_n1001), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT58), .B(G1341), .ZN(new_n1053));
  OAI22_X1  g628(.A1(new_n1051), .A2(G1996), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n564), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT59), .ZN(new_n1057));
  XOR2_X1   g632(.A(new_n1057), .B(KEYINPUT121), .Z(new_n1058));
  XNOR2_X1  g633(.A(new_n1055), .B(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1043), .A2(new_n1046), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1032), .B1(new_n1037), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n741), .A2(G1976), .A3(new_n742), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n1023), .B2(new_n1001), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT52), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n608), .A2(new_n544), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n515), .A2(G48), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n610), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(G1981), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(G305), .B2(G1981), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT49), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1063), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n612), .A2(new_n613), .ZN(new_n1075));
  INV_X1    g650(.A(G1981), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n609), .A4(new_n617), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(KEYINPUT49), .A4(new_n1070), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1073), .A2(new_n1074), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1976), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT52), .B1(G288), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1062), .A2(new_n1064), .A3(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1066), .A2(new_n1080), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n502), .A2(new_n998), .A3(new_n997), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1004), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1050), .A2(KEYINPUT45), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n847), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n785), .B(new_n1004), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(G168), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G8), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT51), .ZN(new_n1092));
  AOI21_X1  g667(.A(G168), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n1094));
  OAI211_X1 g669(.A(G8), .B(new_n1090), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1051), .A2(KEYINPUT114), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1000), .A2(new_n1098), .A3(new_n1004), .A4(new_n1011), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(new_n736), .A3(new_n1099), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1007), .A2(G2090), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G8), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT55), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(KEYINPUT115), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G8), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(KEYINPUT115), .B2(new_n1104), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(G303), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1108), .ZN(new_n1110));
  NOR3_X1   g685(.A1(G166), .A2(new_n1110), .A3(new_n1105), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1103), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1102), .A2(new_n1112), .A3(G8), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1084), .A2(new_n1096), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT45), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1023), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G2078), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n1004), .A4(new_n1085), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1001), .B1(new_n1050), .B2(new_n997), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1123), .A2(KEYINPUT123), .A3(new_n1119), .A4(new_n1118), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1122), .A2(KEYINPUT53), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1007), .A2(new_n797), .ZN(new_n1126));
  AOI21_X1  g701(.A(G2078), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1125), .B(new_n1126), .C1(new_n1127), .C2(KEYINPUT53), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G171), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1010), .A2(KEYINPUT53), .A3(new_n1119), .A4(new_n1011), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1131), .B(G301), .C1(new_n1127), .C2(KEYINPUT53), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT54), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1116), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1131), .B1(new_n1127), .B2(KEYINPUT53), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(new_n1136), .B2(G171), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1128), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT124), .B1(new_n1138), .B2(G301), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1128), .A2(new_n1140), .A3(G171), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1137), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1061), .A2(new_n1134), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1077), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G288), .A2(G1976), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(new_n1080), .B2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1063), .B(KEYINPUT117), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1066), .A2(new_n1080), .A3(new_n1083), .ZN(new_n1149));
  OAI22_X1  g724(.A1(new_n1147), .A2(new_n1148), .B1(new_n1149), .B2(new_n1115), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1091), .A2(G286), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1084), .A2(new_n1114), .A3(new_n1115), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT63), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1102), .A2(new_n1112), .A3(G8), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1112), .B1(new_n1102), .B2(G8), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1157), .A2(KEYINPUT63), .A3(new_n1084), .A4(new_n1151), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1150), .B1(new_n1154), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1143), .A2(new_n1144), .A3(new_n1159), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n1096), .A2(KEYINPUT62), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1155), .A2(new_n1149), .A3(new_n1156), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1129), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1096), .A2(KEYINPUT62), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1161), .A2(new_n1162), .A3(KEYINPUT126), .A4(new_n1163), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1160), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1144), .B1(new_n1143), .B2(new_n1159), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1003), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1002), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1173), .B1(new_n988), .B2(new_n780), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT127), .Z(new_n1175));
  NAND2_X1  g750(.A1(new_n1002), .A2(new_n989), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT46), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT47), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n758), .A2(new_n760), .ZN(new_n1180));
  OAI22_X1  g755(.A1(new_n991), .A2(new_n1180), .B1(G2067), .B2(new_n825), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1002), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n992), .A2(new_n1173), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n993), .A2(new_n1173), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1183), .B1(KEYINPUT48), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(KEYINPUT48), .B2(new_n1184), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1179), .A2(new_n1182), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1172), .A2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g763(.A1(G229), .A2(G227), .A3(new_n460), .ZN(new_n1190));
  OAI21_X1  g764(.A(new_n1190), .B1(new_n689), .B2(new_n690), .ZN(new_n1191));
  AOI21_X1  g765(.A(G37), .B1(new_n890), .B2(new_n893), .ZN(new_n1192));
  AOI21_X1  g766(.A(new_n1191), .B1(new_n1192), .B2(new_n896), .ZN(new_n1193));
  AND3_X1   g767(.A1(new_n1193), .A2(new_n969), .A3(new_n973), .ZN(G308));
  NAND3_X1  g768(.A1(new_n1193), .A2(new_n969), .A3(new_n973), .ZN(G225));
endmodule


