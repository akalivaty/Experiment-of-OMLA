//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n531, new_n532, new_n533, new_n534, new_n535, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n587, new_n588,
    new_n589, new_n592, new_n594, new_n595, new_n596, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n458), .A2(G101), .A3(G2104), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n458), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n465), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(new_n458), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n468), .A2(new_n470), .ZN(G160));
  OAI21_X1  g046(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G112), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n466), .ZN(new_n478));
  AOI211_X1 g053(.A(new_n474), .B(new_n477), .C1(G136), .C2(new_n478), .ZN(G162));
  NAND2_X1  g054(.A1(KEYINPUT4), .A2(G138), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n480), .B1(new_n463), .B2(new_n464), .ZN(new_n481));
  AND2_X1   g056(.A1(G102), .A2(G2104), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n458), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G126), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n463), .B2(new_n464), .ZN(new_n485));
  AND2_X1   g060(.A1(G114), .A2(G2104), .ZN(new_n486));
  OAI21_X1  g061(.A(G2105), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n464), .ZN(new_n488));
  NOR2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n458), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n483), .A2(new_n487), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G164));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT5), .B(G543), .ZN(new_n496));
  AOI21_X1  g071(.A(KEYINPUT68), .B1(new_n496), .B2(G62), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(G75), .B2(G543), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(KEYINPUT68), .A3(G62), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n500), .A2(KEYINPUT69), .ZN(new_n501));
  XOR2_X1   g076(.A(KEYINPUT5), .B(G543), .Z(new_n502));
  AND2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n506), .A2(G88), .B1(new_n508), .B2(G50), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n509), .B1(new_n500), .B2(KEYINPUT69), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n501), .A2(new_n510), .ZN(G303));
  INV_X1    g086(.A(G303), .ZN(G166));
  NAND3_X1  g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT7), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n503), .A2(new_n504), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G51), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(G89), .ZN(new_n519));
  NAND2_X1  g094(.A1(G63), .A2(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n502), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n518), .A2(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  INV_X1    g098(.A(G52), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n515), .A2(new_n496), .ZN(new_n525));
  INV_X1    g100(.A(G90), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n524), .A2(new_n516), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n496), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n495), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n527), .A2(new_n529), .ZN(G171));
  AOI22_X1  g105(.A1(new_n506), .A2(G81), .B1(new_n508), .B2(G43), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT70), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n496), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n495), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G860), .ZN(G153));
  NAND4_X1  g111(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g112(.A1(G1), .A2(G3), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT8), .ZN(new_n539));
  NAND4_X1  g114(.A1(G319), .A2(G483), .A3(G661), .A4(new_n539), .ZN(G188));
  NAND2_X1  g115(.A1(G78), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G65), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n502), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n543), .A2(G651), .B1(new_n506), .B2(G91), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT9), .ZN(new_n545));
  INV_X1    g120(.A(G53), .ZN(new_n546));
  OAI211_X1 g121(.A(KEYINPUT71), .B(new_n545), .C1(new_n516), .C2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n546), .B1(new_n548), .B2(KEYINPUT9), .ZN(new_n549));
  OAI211_X1 g124(.A(new_n508), .B(new_n549), .C1(new_n548), .C2(KEYINPUT9), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n544), .A2(new_n547), .A3(new_n550), .ZN(G299));
  INV_X1    g126(.A(G171), .ZN(G301));
  NAND2_X1  g127(.A1(new_n506), .A2(G87), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT72), .ZN(new_n554));
  OAI21_X1  g129(.A(G651), .B1(new_n496), .B2(G74), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n508), .A2(G49), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(G288));
  INV_X1    g132(.A(G48), .ZN(new_n558));
  INV_X1    g133(.A(G86), .ZN(new_n559));
  OAI22_X1  g134(.A1(new_n558), .A2(new_n516), .B1(new_n525), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n496), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n561), .A2(new_n495), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(G305));
  INV_X1    g139(.A(G47), .ZN(new_n565));
  XOR2_X1   g140(.A(KEYINPUT73), .B(G85), .Z(new_n566));
  OAI22_X1  g141(.A1(new_n565), .A2(new_n516), .B1(new_n525), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n496), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n495), .ZN(new_n569));
  OR3_X1    g144(.A1(new_n567), .A2(KEYINPUT74), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT74), .B1(new_n567), .B2(new_n569), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(G290));
  NAND2_X1  g147(.A1(G301), .A2(G868), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n506), .A2(G92), .ZN(new_n574));
  XOR2_X1   g149(.A(new_n574), .B(KEYINPUT10), .Z(new_n575));
  OR2_X1    g150(.A1(new_n516), .A2(KEYINPUT75), .ZN(new_n576));
  INV_X1    g151(.A(G54), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n516), .B2(KEYINPUT75), .ZN(new_n578));
  NAND2_X1  g153(.A1(G79), .A2(G543), .ZN(new_n579));
  XOR2_X1   g154(.A(KEYINPUT76), .B(G66), .Z(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n502), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n576), .A2(new_n578), .B1(G651), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n575), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n573), .B1(new_n584), .B2(G868), .ZN(G284));
  OAI21_X1  g160(.A(new_n573), .B1(new_n584), .B2(G868), .ZN(G321));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NOR2_X1   g162(.A1(G286), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g163(.A(G299), .B(KEYINPUT77), .Z(new_n589));
  AOI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(new_n587), .ZN(G297));
  AOI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n587), .ZN(G280));
  INV_X1    g166(.A(G559), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n584), .B1(new_n592), .B2(G860), .ZN(G148));
  NAND2_X1  g168(.A1(new_n532), .A2(new_n534), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(new_n587), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n583), .A2(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(new_n587), .ZN(G323));
  XNOR2_X1  g172(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g173(.A1(new_n462), .A2(G2105), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n465), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT12), .ZN(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(G2100), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(G2100), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n475), .A2(G123), .ZN(new_n606));
  OR2_X1    g181(.A1(G99), .A2(G2105), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n607), .B(G2104), .C1(G111), .C2(new_n458), .ZN(new_n608));
  INV_X1    g183(.A(G135), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n606), .B(new_n608), .C1(new_n609), .C2(new_n466), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(G2096), .Z(new_n611));
  NAND3_X1  g186(.A1(new_n604), .A2(new_n605), .A3(new_n611), .ZN(G156));
  INV_X1    g187(.A(KEYINPUT14), .ZN(new_n613));
  XNOR2_X1  g188(.A(G2427), .B(G2438), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2430), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT15), .B(G2435), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n616), .B2(new_n615), .ZN(new_n618));
  XNOR2_X1  g193(.A(G2451), .B(G2454), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT16), .ZN(new_n620));
  XNOR2_X1  g195(.A(G1341), .B(G1348), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n618), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2443), .B(G2446), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(G14), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT79), .Z(G401));
  XOR2_X1   g203(.A(G2084), .B(G2090), .Z(new_n629));
  XNOR2_X1  g204(.A(G2067), .B(G2678), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2072), .B(G2078), .Z(new_n632));
  NOR2_X1   g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT18), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n632), .B(KEYINPUT17), .ZN(new_n635));
  INV_X1    g210(.A(new_n629), .ZN(new_n636));
  INV_X1    g211(.A(new_n630), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n636), .A2(new_n632), .A3(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(new_n631), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n634), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2096), .B(G2100), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(G227));
  XOR2_X1   g218(.A(G1971), .B(G1976), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT19), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1956), .B(G2474), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1961), .B(G1966), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NOR3_X1   g224(.A1(new_n645), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n645), .A2(new_n648), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT80), .B(KEYINPUT20), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  AOI211_X1 g228(.A(new_n650), .B(new_n653), .C1(new_n645), .C2(new_n649), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT81), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1991), .B(G1996), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT82), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1981), .B(G1986), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G229));
  NOR2_X1   g239(.A1(G16), .A2(G23), .ZN(new_n665));
  XNOR2_X1  g240(.A(G288), .B(KEYINPUT83), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n665), .B1(new_n666), .B2(G16), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT33), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(G16), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(G22), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(G166), .B2(new_n670), .ZN(new_n672));
  INV_X1    g247(.A(G1971), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(G6), .A2(G16), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n563), .B2(G16), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT32), .ZN(new_n677));
  INV_X1    g252(.A(G1981), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n669), .A2(new_n674), .A3(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n680), .A2(KEYINPUT34), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(KEYINPUT34), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n475), .A2(G119), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n458), .A2(G107), .ZN(new_n684));
  OAI21_X1  g259(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n685));
  INV_X1    g260(.A(G131), .ZN(new_n686));
  OAI221_X1 g261(.A(new_n683), .B1(new_n684), .B2(new_n685), .C1(new_n686), .C2(new_n466), .ZN(new_n687));
  MUX2_X1   g262(.A(G25), .B(new_n687), .S(G29), .Z(new_n688));
  XOR2_X1   g263(.A(KEYINPUT35), .B(G1991), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n670), .A2(G24), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G290), .B2(G16), .ZN(new_n692));
  INV_X1    g267(.A(G1986), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n693), .B2(new_n692), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n681), .A2(new_n682), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT36), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G35), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G162), .B2(new_n698), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT29), .Z(new_n701));
  INV_X1    g276(.A(G2090), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n670), .A2(G20), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT23), .Z(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G299), .B2(G16), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT93), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n703), .B1(G1956), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G1956), .B2(new_n707), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT94), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n670), .A2(G19), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n535), .B2(new_n670), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(G1341), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n475), .A2(G128), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n458), .A2(G116), .ZN(new_n715));
  OAI21_X1  g290(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n716));
  INV_X1    g291(.A(G140), .ZN(new_n717));
  OAI221_X1 g292(.A(new_n714), .B1(new_n715), .B2(new_n716), .C1(new_n717), .C2(new_n466), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n698), .A2(G26), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G2067), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n701), .B2(new_n702), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n670), .A2(G4), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n584), .B2(new_n670), .ZN(new_n726));
  INV_X1    g301(.A(G1348), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  AND4_X1   g303(.A1(new_n710), .A2(new_n713), .A3(new_n724), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n670), .A2(G21), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G168), .B2(new_n670), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT86), .Z(new_n732));
  INV_X1    g307(.A(G1966), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT88), .Z(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT31), .B(G11), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT87), .B(G28), .ZN(new_n737));
  AOI21_X1  g312(.A(G29), .B1(new_n737), .B2(KEYINPUT30), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(KEYINPUT30), .B2(new_n737), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n736), .B(new_n739), .C1(new_n610), .C2(new_n698), .ZN(new_n740));
  NOR2_X1   g315(.A1(G5), .A2(G16), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT89), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G301), .B2(new_n670), .ZN(new_n743));
  INV_X1    g318(.A(G1961), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G34), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT24), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n746), .B2(KEYINPUT24), .ZN(new_n748));
  AOI22_X1  g323(.A1(G160), .A2(G29), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n745), .B1(G2084), .B2(new_n749), .ZN(new_n750));
  AOI211_X1 g325(.A(new_n740), .B(new_n750), .C1(G2084), .C2(new_n749), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n743), .A2(new_n744), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT90), .Z(new_n753));
  OAI211_X1 g328(.A(new_n751), .B(new_n753), .C1(new_n733), .C2(new_n732), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n698), .A2(G33), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT25), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(new_n458), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n757), .B(new_n759), .C1(G139), .C2(new_n478), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n755), .B1(new_n760), .B2(new_n698), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(G2072), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n698), .A2(G27), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT91), .Z(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n493), .B2(G29), .ZN(new_n765));
  INV_X1    g340(.A(G2078), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n762), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n698), .A2(G32), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n475), .A2(G129), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT84), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n478), .A2(G141), .ZN(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT26), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G105), .B2(new_n599), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n772), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT85), .Z(new_n778));
  OAI21_X1  g353(.A(new_n770), .B1(new_n778), .B2(new_n698), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT27), .B(G1996), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n735), .A2(new_n754), .A3(new_n769), .A4(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT92), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n697), .A2(new_n729), .A3(new_n783), .ZN(G150));
  INV_X1    g359(.A(G150), .ZN(G311));
  INV_X1    g360(.A(G55), .ZN(new_n786));
  INV_X1    g361(.A(G93), .ZN(new_n787));
  OAI22_X1  g362(.A1(new_n786), .A2(new_n516), .B1(new_n525), .B2(new_n787), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n496), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(new_n495), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G860), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT96), .B(KEYINPUT37), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n584), .A2(G559), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT38), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n535), .A2(new_n791), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n594), .B1(new_n790), .B2(new_n788), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n797), .B(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT39), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT95), .Z(new_n804));
  OAI21_X1  g379(.A(new_n792), .B1(new_n801), .B2(new_n802), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n795), .B1(new_n804), .B2(new_n805), .ZN(G145));
  XNOR2_X1  g381(.A(new_n718), .B(new_n493), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(new_n687), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n478), .A2(G142), .B1(G130), .B2(new_n475), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT98), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n812));
  OR3_X1    g387(.A1(new_n812), .A2(new_n458), .A3(G118), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n810), .A2(KEYINPUT98), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n812), .B1(new_n458), .B2(G118), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n811), .A2(new_n813), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n809), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(new_n601), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n808), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n777), .A2(new_n760), .ZN(new_n820));
  INV_X1    g395(.A(new_n778), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n760), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n819), .B(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(G162), .B(new_n610), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G160), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT99), .ZN(new_n827));
  AOI21_X1  g402(.A(G37), .B1(new_n823), .B2(new_n825), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g405(.A(G288), .B(KEYINPUT83), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(new_n563), .ZN(new_n832));
  XNOR2_X1  g407(.A(G290), .B(KEYINPUT101), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(G303), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n666), .A2(G305), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(G303), .ZN(new_n836));
  AND4_X1   g411(.A1(new_n832), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n834), .A2(new_n836), .B1(new_n832), .B2(new_n835), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT42), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n584), .A2(G299), .ZN(new_n841));
  INV_X1    g416(.A(G299), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n583), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT41), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n841), .A2(new_n848), .A3(new_n843), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n583), .A2(KEYINPUT100), .A3(new_n842), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT41), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n800), .B(new_n596), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n845), .B2(new_n853), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n840), .B(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G868), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(G868), .B2(new_n791), .ZN(G295));
  OAI21_X1  g433(.A(new_n857), .B1(G868), .B2(new_n791), .ZN(G331));
  INV_X1    g434(.A(new_n839), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n798), .A2(G301), .A3(new_n799), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(G301), .B1(new_n798), .B2(new_n799), .ZN(new_n863));
  OAI21_X1  g438(.A(G286), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n863), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n865), .A2(G168), .A3(new_n861), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n845), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n864), .B(new_n866), .C1(new_n847), .C2(new_n851), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(G37), .B1(new_n860), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT43), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n839), .A2(new_n868), .A3(new_n869), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n844), .B1(new_n867), .B2(new_n846), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(KEYINPUT103), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(KEYINPUT103), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n879), .A2(new_n866), .A3(new_n864), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n839), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n871), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT43), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n876), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n874), .A2(new_n875), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT44), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n872), .B1(new_n871), .B2(new_n873), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n889), .A2(KEYINPUT102), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n871), .A2(new_n883), .A3(new_n872), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n871), .A2(new_n873), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(KEYINPUT102), .A3(KEYINPUT43), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n890), .A2(new_n891), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n888), .A2(new_n895), .ZN(G397));
  INV_X1    g471(.A(G40), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n468), .A2(new_n470), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G1384), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n493), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT45), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n777), .A3(G1996), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n905), .B(KEYINPUT106), .Z(new_n906));
  XOR2_X1   g481(.A(new_n718), .B(G2067), .Z(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(new_n821), .B2(G1996), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n904), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n687), .B(new_n689), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(G290), .A2(G1986), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT105), .ZN(new_n914));
  NAND2_X1  g489(.A1(G290), .A2(G1986), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n910), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n563), .B(G1981), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT49), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n919), .B(KEYINPUT111), .Z(new_n920));
  NAND3_X1  g495(.A1(new_n898), .A2(new_n900), .A3(new_n493), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(G8), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n920), .B(new_n923), .C1(KEYINPUT49), .C2(new_n918), .ZN(new_n924));
  INV_X1    g499(.A(G1976), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n923), .B1(new_n831), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT52), .B1(G288), .B2(new_n925), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT110), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(KEYINPUT52), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G8), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n493), .A2(KEYINPUT45), .A3(new_n900), .ZN(new_n933));
  INV_X1    g508(.A(new_n903), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n933), .B1(new_n934), .B2(KEYINPUT107), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n933), .A2(KEYINPUT107), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(new_n899), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n673), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n901), .A2(KEYINPUT50), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT50), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n493), .A2(new_n941), .A3(new_n900), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(KEYINPUT108), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n941), .B1(new_n493), .B2(new_n900), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n947), .A2(new_n702), .A3(new_n898), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n932), .B1(new_n939), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(G303), .A2(G8), .ZN(new_n950));
  NAND2_X1  g525(.A1(KEYINPUT109), .A2(KEYINPUT55), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n953));
  NAND3_X1  g528(.A1(G303), .A2(G8), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n931), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n940), .A2(new_n898), .A3(new_n942), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n939), .B1(G2090), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n955), .B1(new_n959), .B2(G8), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT114), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n903), .A2(new_n933), .A3(new_n898), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n733), .ZN(new_n964));
  INV_X1    g539(.A(G2084), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n898), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n943), .B2(new_n946), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI211_X1 g544(.A(KEYINPUT115), .B(new_n966), .C1(new_n943), .C2(new_n946), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT122), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(G286), .A2(G8), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n972), .B(KEYINPUT123), .Z(new_n973));
  INV_X1    g548(.A(new_n966), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n493), .A2(new_n941), .A3(new_n900), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n975), .A2(new_n944), .A3(new_n945), .ZN(new_n976));
  INV_X1    g551(.A(new_n946), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT115), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n967), .A2(new_n968), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT122), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n979), .A2(new_n980), .A3(new_n981), .A4(new_n964), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n971), .A2(new_n973), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n973), .A2(KEYINPUT51), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(new_n980), .A3(new_n964), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT125), .B1(new_n985), .B2(G8), .ZN(new_n986));
  OAI211_X1 g561(.A(KEYINPUT125), .B(G8), .C1(new_n969), .C2(new_n970), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n984), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n971), .A2(G8), .A3(new_n982), .ZN(new_n991));
  INV_X1    g566(.A(new_n973), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n989), .B1(new_n993), .B2(KEYINPUT124), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT124), .ZN(new_n995));
  AOI211_X1 g570(.A(new_n995), .B(new_n990), .C1(new_n991), .C2(new_n992), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n983), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT62), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n999), .B(new_n983), .C1(new_n994), .C2(new_n996), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n898), .B1(new_n976), .B2(new_n977), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT118), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n947), .A2(KEYINPUT118), .A3(new_n898), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n935), .A2(new_n766), .A3(new_n937), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n1005), .A2(new_n744), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n766), .A2(KEYINPUT53), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n963), .B2(new_n1009), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1010), .A2(G171), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n998), .A2(new_n1000), .A3(new_n1011), .ZN(new_n1012));
  XOR2_X1   g587(.A(G171), .B(KEYINPUT54), .Z(new_n1013));
  INV_X1    g588(.A(new_n1007), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n1014), .B2(KEYINPUT53), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1010), .A2(new_n1013), .B1(new_n1008), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1956), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n958), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n958), .A2(KEYINPUT117), .A3(new_n1017), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(G299), .B(KEYINPUT57), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(KEYINPUT56), .B(G2072), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n935), .A2(new_n937), .A3(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1024), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT120), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT61), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT61), .ZN(new_n1032));
  OAI211_X1 g607(.A(KEYINPUT120), .B(new_n1032), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT58), .B(G1341), .Z(new_n1034));
  NAND2_X1  g609(.A1(new_n921), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n938), .B2(G1996), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n594), .B1(KEYINPUT119), .B2(KEYINPUT59), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OR2_X1    g613(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1031), .A2(new_n1033), .A3(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1003), .A2(new_n727), .A3(new_n1004), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n921), .A2(G2067), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT60), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT60), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1046), .B1(new_n1048), .B2(new_n584), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1003), .A2(new_n727), .A3(new_n1004), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1043), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT60), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1052), .A2(KEYINPUT121), .A3(new_n583), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1045), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1048), .A2(new_n1046), .A3(new_n584), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT121), .B1(new_n1052), .B2(new_n583), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1055), .A2(KEYINPUT60), .A3(new_n1056), .A4(new_n1044), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1041), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n584), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1029), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1028), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n997), .B(new_n1016), .C1(new_n1058), .C2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n962), .B1(new_n1012), .B2(new_n1062), .ZN(new_n1063));
  OR2_X1    g638(.A1(new_n949), .A2(KEYINPUT116), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n949), .A2(KEYINPUT116), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1064), .A2(new_n954), .A3(new_n952), .A4(new_n1065), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n985), .A2(G8), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G168), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n957), .A2(KEYINPUT63), .A3(new_n1066), .A4(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n962), .A2(new_n1068), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(KEYINPUT63), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n922), .B(KEYINPUT112), .ZN(new_n1073));
  NOR2_X1   g648(.A1(G288), .A2(G1976), .ZN(new_n1074));
  XOR2_X1   g649(.A(new_n1074), .B(KEYINPUT113), .Z(new_n1075));
  NAND2_X1  g650(.A1(new_n924), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n563), .A2(new_n678), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1073), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n931), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n956), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1072), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n917), .B1(new_n1063), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT46), .ZN(new_n1083));
  OR3_X1    g658(.A1(new_n910), .A2(new_n1083), .A3(G1996), .ZN(new_n1084));
  INV_X1    g659(.A(new_n907), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n904), .B1(new_n1085), .B2(new_n777), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1083), .B1(new_n910), .B2(G1996), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1088), .B(KEYINPUT47), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n718), .A2(G2067), .ZN(new_n1090));
  INV_X1    g665(.A(new_n689), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n687), .A2(new_n1091), .ZN(new_n1092));
  XOR2_X1   g667(.A(new_n1092), .B(KEYINPUT126), .Z(new_n1093));
  AOI21_X1  g668(.A(new_n1090), .B1(new_n909), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1089), .B1(new_n1094), .B2(new_n910), .ZN(new_n1095));
  XOR2_X1   g670(.A(new_n912), .B(KEYINPUT127), .Z(new_n1096));
  NOR2_X1   g671(.A1(new_n914), .A2(new_n910), .ZN(new_n1097));
  XOR2_X1   g672(.A(new_n1097), .B(KEYINPUT48), .Z(new_n1098));
  AOI21_X1  g673(.A(new_n1095), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1082), .A2(new_n1099), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g675(.A(new_n627), .ZN(new_n1102));
  INV_X1    g676(.A(G319), .ZN(new_n1103));
  NOR3_X1   g677(.A1(new_n1102), .A2(new_n1103), .A3(G227), .ZN(new_n1104));
  NAND3_X1  g678(.A1(new_n663), .A2(new_n829), .A3(new_n1104), .ZN(new_n1105));
  AND2_X1   g679(.A1(new_n890), .A2(new_n892), .ZN(new_n1106));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n1106), .B2(new_n894), .ZN(G308));
  AND2_X1   g681(.A1(new_n663), .A2(new_n1104), .ZN(new_n1108));
  INV_X1    g682(.A(new_n894), .ZN(new_n1109));
  NAND2_X1  g683(.A1(new_n890), .A2(new_n892), .ZN(new_n1110));
  OAI211_X1 g684(.A(new_n1108), .B(new_n829), .C1(new_n1109), .C2(new_n1110), .ZN(G225));
endmodule


