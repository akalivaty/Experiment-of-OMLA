//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G50), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND3_X1  g0015(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n203), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n205), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n212), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  NAND3_X1  g0043(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(G1), .A2(G13), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n247), .B1(G1), .B2(new_n210), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G50), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n204), .A2(new_n210), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n246), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT65), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n250), .B1(G50), .B2(new_n251), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n261), .A2(new_n262), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g0065(.A(new_n265), .B(KEYINPUT9), .Z(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G222), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(G1698), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n269), .B1(new_n205), .B2(new_n267), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  OAI211_X1 g0073(.A(G1), .B(G13), .C1(new_n257), .C2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G274), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n275), .A2(new_n278), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(G226), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G200), .ZN(new_n284));
  INV_X1    g0084(.A(G190), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(new_n283), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n266), .A2(new_n286), .B1(KEYINPUT67), .B2(KEYINPUT10), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT67), .A2(KEYINPUT10), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G169), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n283), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n265), .B(new_n291), .C1(G179), .C2(new_n283), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n267), .A2(G226), .A3(new_n268), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G97), .ZN(new_n295));
  INV_X1    g0095(.A(G232), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n294), .B(new_n295), .C1(new_n270), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n275), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT13), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n280), .B1(new_n281), .B2(G238), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n299), .B1(new_n298), .B2(new_n300), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT14), .B1(new_n304), .B2(new_n290), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT14), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n306), .B(G169), .C1(new_n302), .C2(new_n303), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(G179), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n209), .A2(G13), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n202), .A2(G20), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT69), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT12), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(G68), .B2(new_n249), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n252), .A2(KEYINPUT68), .A3(G50), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(new_n311), .C1(new_n259), .C2(new_n205), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT68), .B1(new_n252), .B2(G50), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n246), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT11), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n319), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n314), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n309), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n322), .B1(new_n304), .B2(G190), .ZN(new_n325));
  INV_X1    g0125(.A(G200), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n304), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n256), .A2(new_n253), .B1(new_n210), .B2(new_n205), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT15), .B(G87), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n328), .A2(KEYINPUT66), .B1(new_n258), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(KEYINPUT66), .B2(new_n328), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n246), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n249), .A2(G77), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n333), .B(new_n334), .C1(G77), .C2(new_n251), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G33), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G107), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n267), .A2(new_n268), .ZN(new_n341));
  INV_X1    g0141(.A(G238), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n340), .B1(new_n341), .B2(new_n296), .C1(new_n342), .C2(new_n270), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n275), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n280), .B1(new_n281), .B2(G244), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n290), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n344), .A2(new_n348), .A3(new_n345), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n335), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n346), .A2(new_n285), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n326), .B1(new_n344), .B2(new_n345), .ZN(new_n352));
  OR3_X1    g0152(.A1(new_n335), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n327), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n293), .A2(new_n324), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT17), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT70), .ZN(new_n357));
  INV_X1    g0157(.A(G159), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n253), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G58), .A2(G68), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n210), .B1(new_n203), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n357), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n360), .ZN(new_n363));
  NOR2_X1   g0163(.A1(G58), .A2(G68), .ZN(new_n364));
  OAI21_X1  g0164(.A(G20), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n365), .B(KEYINPUT70), .C1(new_n358), .C2(new_n253), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT7), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n267), .B2(G20), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n339), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n202), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT16), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT16), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n336), .A2(KEYINPUT71), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT71), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(new_n257), .A3(KEYINPUT3), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n338), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n368), .A2(G20), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n202), .B1(new_n380), .B2(new_n369), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n374), .B1(new_n381), .B2(new_n367), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n373), .A2(new_n382), .A3(new_n246), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n256), .A2(new_n251), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n249), .B2(new_n256), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT73), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n271), .A2(G1698), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(new_n336), .A3(new_n338), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT72), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n336), .A2(new_n338), .A3(G226), .A4(G1698), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT72), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n389), .A2(new_n336), .A3(new_n338), .A4(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n391), .A2(new_n392), .A3(new_n393), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n275), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n274), .A2(G232), .A3(new_n277), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n279), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n388), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  AOI211_X1 g0201(.A(KEYINPUT73), .B(new_n399), .C1(new_n396), .C2(new_n275), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n326), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT75), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n394), .B1(new_n267), .B2(new_n389), .ZN(new_n405));
  AND4_X1   g0205(.A1(new_n394), .A2(new_n389), .A3(new_n336), .A4(new_n338), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n393), .A2(new_n392), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n274), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n409), .A2(G190), .A3(new_n399), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n403), .A2(new_n404), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n404), .B1(new_n403), .B2(new_n411), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n387), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT76), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT73), .B1(new_n409), .B2(new_n399), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n397), .A2(new_n388), .A3(new_n400), .ZN(new_n417));
  AOI21_X1  g0217(.A(G200), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT75), .B1(new_n418), .B2(new_n410), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n403), .A2(new_n404), .A3(new_n411), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT76), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(new_n387), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n356), .B1(new_n415), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n386), .B1(new_n419), .B2(new_n420), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(KEYINPUT17), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT77), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n422), .B1(new_n421), .B2(new_n387), .ZN(new_n428));
  AOI211_X1 g0228(.A(KEYINPUT76), .B(new_n386), .C1(new_n419), .C2(new_n420), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT17), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT77), .ZN(new_n431));
  INV_X1    g0231(.A(new_n426), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n290), .B1(new_n401), .B2(new_n402), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n397), .A2(new_n348), .A3(new_n400), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n386), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT18), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n439), .A3(new_n386), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT74), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT74), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n438), .A2(new_n443), .A3(new_n440), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n427), .A2(new_n433), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n355), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT4), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n341), .B2(new_n219), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n267), .A2(KEYINPUT4), .A3(G244), .A4(new_n268), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n267), .A2(G250), .A3(G1698), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n275), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n209), .B(G45), .C1(new_n273), .C2(KEYINPUT5), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT83), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n456), .A2(new_n457), .B1(KEYINPUT5), .B2(new_n273), .ZN(new_n458));
  INV_X1    g0258(.A(G45), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(G1), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(KEYINPUT83), .C1(KEYINPUT5), .C2(new_n273), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n275), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n456), .A2(new_n457), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n273), .A2(KEYINPUT5), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G274), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n275), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g0267(.A1(G257), .A2(new_n462), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(G169), .B1(new_n455), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n455), .A2(new_n468), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n469), .B1(new_n471), .B2(new_n348), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT7), .B1(new_n339), .B2(new_n210), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n378), .B2(new_n379), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT81), .B1(new_n474), .B2(new_n220), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n380), .A2(new_n369), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT81), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(G107), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n252), .A2(G77), .ZN(new_n479));
  XOR2_X1   g0279(.A(new_n479), .B(KEYINPUT78), .Z(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT79), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT79), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G97), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n485), .A2(KEYINPUT80), .A3(KEYINPUT6), .A4(new_n220), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT80), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT79), .B(G97), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n220), .A2(KEYINPUT6), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT6), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n481), .A2(new_n220), .ZN(new_n492));
  NOR2_X1   g0292(.A1(G97), .A2(G107), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n486), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n480), .B1(new_n495), .B2(G20), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n475), .A2(new_n478), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n246), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n209), .A2(G33), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n251), .A2(new_n499), .A3(new_n245), .A4(new_n244), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT82), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G97), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n251), .A2(new_n481), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n472), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n460), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n274), .A2(G250), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n466), .B2(new_n508), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G116), .ZN(new_n511));
  OAI221_X1 g0311(.A(new_n511), .B1(new_n341), .B2(new_n342), .C1(new_n219), .C2(new_n270), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n510), .B1(new_n512), .B2(new_n275), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(G169), .ZN(new_n514));
  AOI211_X1 g0314(.A(G179), .B(new_n510), .C1(new_n512), .C2(new_n275), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT84), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n502), .B2(new_n329), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n500), .B(KEYINPUT82), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n519), .A2(KEYINPUT84), .A3(new_n330), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT85), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n330), .A2(new_n251), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT19), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n488), .B2(new_n259), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n210), .B1(new_n295), .B2(new_n524), .ZN(new_n526));
  INV_X1    g0326(.A(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n220), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n485), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n267), .A2(new_n210), .A3(G68), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n525), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n523), .B1(new_n531), .B2(new_n246), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n521), .A2(new_n522), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n522), .B1(new_n521), .B2(new_n532), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n516), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n513), .A2(new_n326), .ZN(new_n536));
  AOI211_X1 g0336(.A(new_n285), .B(new_n510), .C1(new_n512), .C2(new_n275), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n532), .B1(new_n527), .B2(new_n502), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n497), .A2(new_n246), .B1(new_n503), .B2(new_n504), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n470), .A2(G200), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n455), .A2(G190), .A3(new_n468), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n507), .A2(new_n535), .A3(new_n540), .A4(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n462), .A2(G264), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n267), .A2(G250), .A3(new_n268), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n267), .A2(G257), .A3(G1698), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G294), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n275), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n465), .A2(new_n467), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(G179), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n547), .A2(new_n554), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n551), .A2(KEYINPUT88), .A3(new_n275), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT88), .B1(new_n551), .B2(new_n275), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n555), .B1(new_n559), .B2(new_n290), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n210), .A2(G107), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT23), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT86), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n258), .A2(G116), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n562), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT86), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n566), .B(KEYINPUT23), .C1(new_n210), .C2(G107), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n563), .A2(new_n564), .A3(new_n565), .A4(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n562), .A2(new_n561), .B1(new_n258), .B2(G116), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n571), .A2(KEYINPUT87), .A3(new_n563), .A4(new_n567), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n267), .A2(new_n210), .A3(G87), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n574), .B(KEYINPUT22), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT24), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT24), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n573), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n247), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n519), .A2(G107), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n251), .A2(G107), .ZN(new_n582));
  XNOR2_X1  g0382(.A(new_n582), .B(KEYINPUT25), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n560), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n559), .A2(KEYINPUT89), .A3(new_n285), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT89), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT88), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n552), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n551), .A2(KEYINPUT88), .A3(new_n275), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n589), .A2(new_n590), .A3(new_n554), .A4(new_n547), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n587), .B1(new_n591), .B2(G190), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n553), .A2(new_n554), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n326), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n586), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n580), .A2(new_n584), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT20), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n451), .A2(new_n210), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n485), .B2(new_n257), .ZN(new_n600));
  INV_X1    g0400(.A(G116), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n244), .A2(new_n245), .B1(G20), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n598), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n488), .A2(G33), .ZN(new_n605));
  OAI211_X1 g0405(.A(KEYINPUT20), .B(new_n602), .C1(new_n605), .C2(new_n599), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  MUX2_X1   g0407(.A(new_n251), .B(new_n500), .S(G116), .Z(new_n608));
  AOI21_X1  g0408(.A(new_n290), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n267), .A2(G257), .A3(new_n268), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n339), .A2(G303), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n610), .B(new_n611), .C1(new_n270), .C2(new_n221), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n275), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n462), .A2(G270), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(new_n554), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n609), .A2(KEYINPUT21), .A3(new_n615), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n607), .A2(new_n608), .ZN(new_n620));
  AOI22_X1  g0420(.A1(G270), .A2(new_n462), .B1(new_n465), .B2(new_n467), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n620), .A2(G179), .A3(new_n613), .A4(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(G190), .A3(new_n613), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n620), .B1(new_n615), .B2(G200), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n546), .A2(new_n585), .A3(new_n597), .A4(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n448), .A2(new_n627), .ZN(G372));
  INV_X1    g0428(.A(new_n441), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n427), .A2(new_n433), .ZN(new_n630));
  INV_X1    g0430(.A(new_n350), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n324), .B1(new_n327), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n629), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n289), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(new_n292), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n472), .A2(new_n506), .A3(KEYINPUT91), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT91), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n470), .A2(new_n290), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n455), .A2(new_n348), .A3(new_n468), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n637), .B1(new_n640), .B2(new_n541), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n636), .A2(new_n641), .A3(new_n535), .A4(new_n540), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n534), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n521), .A2(new_n522), .A3(new_n532), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n539), .B1(new_n647), .B2(new_n516), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n640), .A2(new_n541), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n648), .A2(KEYINPUT92), .A3(KEYINPUT26), .A4(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n649), .A2(new_n535), .A3(new_n540), .A4(KEYINPUT26), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT92), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n644), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n648), .A2(new_n597), .A3(new_n507), .A4(new_n544), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n573), .A2(new_n575), .A3(new_n578), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n578), .B1(new_n573), .B2(new_n575), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n246), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n584), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n591), .A2(G169), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n658), .A2(new_n659), .B1(new_n660), .B2(new_n555), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT90), .B1(new_n661), .B2(new_n623), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT90), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n619), .A2(new_n622), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT21), .B1(new_n609), .B2(new_n615), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n585), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n535), .B1(new_n655), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n654), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n635), .B1(new_n448), .B2(new_n670), .ZN(G369));
  NAND3_X1  g0471(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  XOR2_X1   g0473(.A(new_n673), .B(KEYINPUT93), .Z(new_n674));
  OAI21_X1  g0474(.A(G213), .B1(new_n672), .B2(KEYINPUT27), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G343), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n623), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n585), .A2(new_n677), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT95), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n597), .B(new_n585), .C1(new_n596), .C2(new_n677), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n677), .B(KEYINPUT96), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n585), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n677), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n620), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n626), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n666), .B2(new_n688), .ZN(new_n690));
  XNOR2_X1  g0490(.A(KEYINPUT94), .B(G330), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n680), .A2(new_n681), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n686), .A2(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n213), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G1), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n488), .A2(new_n527), .A3(new_n220), .A4(new_n601), .ZN(new_n700));
  OAI22_X1  g0500(.A1(new_n699), .A2(new_n700), .B1(new_n217), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  INV_X1    g0502(.A(new_n535), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n662), .A2(new_n667), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n595), .A2(new_n596), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n545), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n703), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n644), .A2(new_n650), .A3(new_n653), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n684), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n709), .A2(KEYINPUT29), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n649), .A2(new_n535), .A3(new_n540), .A4(new_n643), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n711), .A2(new_n535), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n642), .A2(KEYINPUT26), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT98), .B1(new_n661), .B2(new_n623), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT98), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n585), .A2(new_n715), .A3(new_n666), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n712), .B(new_n713), .C1(new_n655), .C2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT29), .A3(new_n677), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n710), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n627), .A2(new_n684), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n513), .A2(G179), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(new_n593), .A3(new_n470), .A4(new_n615), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n553), .A2(new_n513), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n615), .A2(new_n348), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(new_n471), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT30), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n725), .A2(new_n471), .A3(new_n729), .A4(new_n726), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n724), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n687), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(KEYINPUT97), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n734), .B1(new_n731), .B2(new_n677), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT97), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n721), .A2(new_n735), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n691), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n720), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n702), .B1(new_n743), .B2(G1), .ZN(G364));
  INV_X1    g0544(.A(G13), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n209), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n697), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n692), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n691), .B2(new_n690), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n749), .B(KEYINPUT99), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n696), .A2(new_n339), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G355), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(G116), .B2(new_n213), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n696), .A2(new_n267), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n217), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n757), .B1(new_n459), .B2(new_n758), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n239), .A2(new_n459), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n755), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n245), .B1(G20), .B2(new_n290), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n752), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n765), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n210), .A2(new_n285), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n348), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G322), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n210), .A2(G190), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n771), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n772), .A2(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n326), .A2(G179), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n770), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n267), .B(new_n777), .C1(G303), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n778), .A2(new_n774), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G179), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n774), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G283), .A2(new_n783), .B1(new_n786), .B2(G329), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n348), .A2(new_n326), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n770), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n788), .A2(new_n774), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT33), .B(G317), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G326), .A2(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n210), .B1(new_n784), .B2(G190), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G294), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n781), .A2(new_n787), .A3(new_n794), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n785), .A2(new_n358), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT32), .ZN(new_n800));
  INV_X1    g0600(.A(G50), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n789), .A2(new_n801), .B1(new_n775), .B2(new_n205), .ZN(new_n802));
  INV_X1    g0602(.A(new_n772), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(G58), .B2(new_n803), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n202), .A2(new_n791), .B1(new_n779), .B2(new_n527), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n782), .A2(new_n220), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n805), .A2(new_n339), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n796), .A2(G97), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n800), .A2(new_n804), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n769), .B1(new_n798), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n768), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n764), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n690), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n751), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  INV_X1    g0615(.A(new_n752), .ZN(new_n816));
  INV_X1    g0616(.A(new_n775), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G143), .A2(new_n803), .B1(new_n817), .B2(G159), .ZN(new_n818));
  INV_X1    g0618(.A(G137), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n818), .B1(new_n819), .B2(new_n789), .C1(new_n254), .C2(new_n791), .ZN(new_n820));
  XOR2_X1   g0620(.A(KEYINPUT100), .B(KEYINPUT34), .Z(new_n821));
  XNOR2_X1  g0621(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n796), .A2(G58), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n339), .B1(new_n780), .B2(G50), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n782), .A2(new_n202), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G132), .B2(new_n786), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n791), .A2(new_n828), .B1(new_n775), .B2(new_n601), .ZN(new_n829));
  INV_X1    g0629(.A(G294), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n772), .A2(new_n830), .B1(new_n782), .B2(new_n527), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n267), .B1(new_n780), .B2(G107), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n790), .A2(G303), .B1(new_n786), .B2(G311), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n832), .A2(new_n808), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n769), .B1(new_n827), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n765), .A2(new_n762), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n816), .B(new_n836), .C1(new_n205), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n335), .A2(new_n687), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n353), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n350), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n631), .A2(new_n677), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n838), .B1(new_n844), .B2(new_n763), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT101), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n709), .B(new_n844), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n847), .A2(new_n741), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n749), .B1(new_n847), .B2(new_n741), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G384));
  NAND2_X1  g0651(.A1(new_n360), .A2(G77), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n217), .A2(new_n852), .B1(G50), .B2(new_n202), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(G1), .A3(new_n745), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT102), .Z(new_n855));
  AOI211_X1 g0655(.A(new_n601), .B(new_n216), .C1(new_n495), .C2(KEYINPUT35), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(KEYINPUT35), .B2(new_n495), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT36), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n858), .B2(new_n857), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n676), .B(KEYINPUT105), .Z(new_n861));
  NOR2_X1   g0661(.A1(new_n629), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n428), .A2(new_n429), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n861), .A2(new_n386), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n437), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n373), .A2(new_n246), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n372), .A2(KEYINPUT16), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n385), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n436), .B2(new_n676), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n415), .A2(new_n423), .A3(new_n873), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n864), .A2(new_n869), .B1(new_n874), .B2(KEYINPUT37), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n872), .A2(new_n676), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(new_n446), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n877), .A2(KEYINPUT38), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n879), .B(new_n875), .C1(new_n446), .C2(new_n876), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n842), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n709), .B2(new_n844), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n309), .A2(KEYINPUT103), .A3(new_n322), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT103), .B1(new_n309), .B2(new_n322), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n687), .A2(new_n322), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n327), .A2(new_n886), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n309), .A2(new_n322), .A3(new_n687), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT104), .B1(new_n883), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n683), .B(new_n844), .C1(new_n654), .C2(new_n669), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n842), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT104), .ZN(new_n894));
  INV_X1    g0694(.A(new_n890), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n863), .B1(new_n881), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n878), .A2(new_n880), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT107), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n430), .A2(new_n432), .A3(new_n629), .ZN(new_n902));
  INV_X1    g0702(.A(new_n865), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n864), .A2(new_n869), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n868), .B1(new_n866), .B2(new_n425), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n902), .A2(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n901), .B1(new_n906), .B2(KEYINPUT38), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n415), .A2(new_n423), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n426), .B1(new_n908), .B2(KEYINPUT17), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n865), .B1(new_n909), .B2(new_n629), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n904), .A2(new_n905), .ZN(new_n911));
  OAI211_X1 g0711(.A(KEYINPUT107), .B(new_n879), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n446), .A2(new_n876), .ZN(new_n914));
  INV_X1    g0714(.A(new_n875), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT39), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n900), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n884), .A2(new_n885), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n919), .A2(new_n687), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n898), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT108), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n355), .A2(new_n447), .A3(new_n710), .A4(new_n719), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n635), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n721), .A2(new_n736), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n890), .A2(new_n843), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n878), .B2(new_n880), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n902), .A2(new_n903), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n904), .A2(new_n905), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT107), .B1(new_n935), .B2(new_n879), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n906), .A2(new_n901), .A3(KEYINPUT38), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n916), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n929), .A2(new_n932), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n931), .A2(new_n932), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n448), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n941), .A2(new_n927), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n940), .A2(new_n941), .A3(new_n927), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(new_n691), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n925), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n209), .B2(new_n746), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n925), .A2(new_n945), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n860), .B1(new_n947), .B2(new_n948), .ZN(G367));
  INV_X1    g0749(.A(new_n678), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n693), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n507), .A2(new_n544), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n683), .A2(new_n541), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n952), .A2(KEYINPUT109), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(KEYINPUT109), .B1(new_n952), .B2(new_n953), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n649), .A2(new_n684), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT42), .B1(new_n951), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT42), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n682), .A2(new_n960), .A3(new_n957), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n585), .B1(new_n954), .B2(new_n955), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n683), .B1(new_n962), .B2(new_n649), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n959), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n687), .A2(new_n538), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n648), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n535), .B2(new_n965), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT43), .Z(new_n968));
  NAND2_X1  g0768(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n959), .A2(new_n970), .A3(new_n961), .A4(new_n963), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT110), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n969), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT111), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n971), .B(new_n972), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(KEYINPUT111), .A3(new_n969), .ZN(new_n979));
  INV_X1    g0779(.A(new_n694), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n977), .A2(new_n979), .A3(new_n980), .A4(new_n957), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n975), .A2(new_n976), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT111), .B1(new_n978), .B2(new_n969), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n982), .A2(new_n983), .B1(new_n694), .B2(new_n958), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n697), .B(KEYINPUT41), .Z(new_n985));
  INV_X1    g0785(.A(KEYINPUT45), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT112), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n686), .B2(new_n957), .ZN(new_n988));
  NOR4_X1   g0788(.A1(new_n682), .A2(new_n958), .A3(KEYINPUT112), .A4(new_n685), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n685), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n951), .A2(new_n991), .A3(new_n957), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT112), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n686), .A2(new_n987), .A3(new_n957), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n993), .A2(KEYINPUT45), .A3(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT44), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n686), .B2(new_n957), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n958), .B(KEYINPUT44), .C1(new_n682), .C2(new_n685), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n990), .A2(new_n995), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n980), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT113), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n680), .A2(new_n681), .A3(new_n678), .ZN(new_n1003));
  AND3_X1   g0803(.A1(new_n951), .A2(new_n692), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n692), .B1(new_n951), .B2(new_n1003), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1002), .B1(new_n742), .B2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1006), .A2(new_n720), .A3(KEYINPUT113), .A4(new_n741), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n990), .A2(new_n995), .A3(new_n694), .A4(new_n999), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1001), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n985), .B1(new_n1011), .B2(new_n743), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n981), .B(new_n984), .C1(new_n1012), .C2(new_n748), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n766), .B1(new_n213), .B2(new_n329), .C1(new_n757), .C2(new_n235), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n752), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n267), .B1(new_n790), .B2(G311), .ZN(new_n1016));
  INV_X1    g0816(.A(G317), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1016), .B1(new_n1017), .B2(new_n785), .C1(new_n488), .C2(new_n782), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G294), .A2(new_n792), .B1(new_n803), .B2(G303), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n828), .B2(new_n775), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n780), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT46), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n779), .B2(new_n601), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1021), .B(new_n1023), .C1(new_n220), .C2(new_n795), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1018), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n796), .A2(G68), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n201), .B2(new_n779), .C1(new_n254), .C2(new_n772), .ZN(new_n1027));
  INV_X1    g0827(.A(G143), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n789), .A2(new_n1028), .B1(new_n785), .B2(new_n819), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n791), .A2(new_n358), .B1(new_n775), .B2(new_n801), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n782), .A2(new_n205), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1032), .A2(new_n339), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT114), .Z(new_n1034));
  AOI21_X1  g0834(.A(new_n1025), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT47), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1015), .B1(new_n769), .B2(new_n1036), .C1(new_n967), .C2(new_n812), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1013), .A2(new_n1037), .ZN(G387));
  NAND2_X1  g0838(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1039), .B(new_n697), .C1(new_n743), .C2(new_n1006), .ZN(new_n1040));
  AOI211_X1 g0840(.A(G45), .B(new_n700), .C1(G68), .C2(G77), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n256), .A2(G50), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT50), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n757), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n459), .B2(new_n232), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n753), .A2(new_n700), .B1(new_n220), .B2(new_n696), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(KEYINPUT115), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n766), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT115), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n752), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n202), .A2(new_n775), .B1(new_n782), .B2(new_n481), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n339), .B(new_n1051), .C1(G159), .C2(new_n790), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n256), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G50), .A2(new_n803), .B1(new_n792), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G77), .A2(new_n780), .B1(new_n786), .B2(G150), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n795), .A2(new_n329), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .A4(new_n1057), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n779), .A2(new_n830), .B1(new_n795), .B2(new_n828), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n772), .A2(new_n1017), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n789), .A2(new_n773), .B1(new_n791), .B2(new_n776), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(G303), .C2(new_n817), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1059), .B1(new_n1062), .B2(KEYINPUT48), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(KEYINPUT48), .B2(new_n1062), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT49), .Z(new_n1065));
  AOI21_X1  g0865(.A(new_n267), .B1(new_n786), .B2(G326), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n601), .B2(new_n782), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1058), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1050), .B1(new_n1068), .B2(new_n765), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n693), .B2(new_n812), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1007), .B2(new_n747), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1040), .A2(new_n1072), .ZN(G393));
  NAND2_X1  g0873(.A1(new_n1001), .A2(new_n1010), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n1039), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n1011), .A3(new_n697), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1001), .A2(new_n748), .A3(new_n1010), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n766), .B1(new_n213), .B2(new_n488), .C1(new_n757), .C2(new_n242), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n752), .A2(new_n1078), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n267), .B(new_n806), .C1(G116), .C2(new_n796), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G303), .A2(new_n792), .B1(new_n817), .B2(G294), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G283), .A2(new_n780), .B1(new_n786), .B2(G322), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n789), .A2(new_n1017), .B1(new_n772), .B2(new_n776), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n795), .A2(new_n205), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n339), .B(new_n1087), .C1(G87), .C2(new_n783), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n792), .A2(G50), .B1(new_n817), .B2(new_n1053), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G68), .A2(new_n780), .B1(new_n786), .B2(G143), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n789), .A2(new_n254), .B1(new_n772), .B2(new_n358), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT51), .Z(new_n1093));
  OAI22_X1  g0893(.A1(new_n1083), .A2(new_n1086), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1079), .B1(new_n1094), .B2(new_n765), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n957), .B2(new_n812), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1077), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1076), .A2(new_n1097), .ZN(G390));
  INV_X1    g0898(.A(new_n920), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n883), .B2(new_n890), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n900), .B2(new_n917), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n718), .A2(new_n677), .A3(new_n841), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n842), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT117), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1102), .A2(KEYINPUT117), .A3(new_n842), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n890), .A2(KEYINPUT118), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT118), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n888), .B2(new_n889), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1105), .A2(new_n1106), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n938), .A2(new_n1099), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n735), .A2(new_n738), .A3(new_n739), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n627), .A2(new_n684), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n691), .B(new_n844), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n895), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1101), .A2(new_n1112), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n927), .A2(new_n928), .A3(G330), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n1101), .B2(new_n1112), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n938), .A2(new_n899), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n914), .A2(new_n915), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n879), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1124), .A2(KEYINPUT39), .A3(new_n916), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n762), .ZN(new_n1127));
  INV_X1    g0927(.A(G125), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n791), .A2(new_n819), .B1(new_n785), .B2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT54), .B(G143), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n339), .B(new_n1129), .C1(new_n817), .C2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n796), .A2(G159), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n779), .A2(new_n254), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT53), .ZN(new_n1135));
  INV_X1    g0935(.A(G132), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n772), .A2(new_n1136), .B1(new_n782), .B2(new_n801), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G128), .B2(new_n790), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1132), .A2(new_n1133), .A3(new_n1135), .A4(new_n1138), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1087), .B(new_n825), .C1(G294), .C2(new_n786), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n339), .B1(new_n779), .B2(new_n527), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT120), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n792), .A2(G107), .B1(new_n817), .B2(new_n485), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G283), .A2(new_n790), .B1(new_n803), .B2(G116), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1140), .A2(new_n1142), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n769), .B1(new_n1139), .B2(new_n1145), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n816), .B(new_n1146), .C1(new_n256), .C2(new_n837), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1121), .A2(new_n748), .B1(new_n1127), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1101), .A2(new_n1112), .A3(new_n1117), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1111), .A2(new_n1099), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n907), .A2(new_n912), .B1(new_n877), .B2(KEYINPUT38), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n1126), .B2(new_n1100), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1149), .B1(new_n1153), .B2(new_n1119), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n927), .A2(G330), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n635), .B(new_n923), .C1(new_n448), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1115), .A2(new_n890), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n883), .B1(new_n1157), .B2(new_n1119), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1110), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n927), .A2(G330), .A3(new_n844), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1116), .A2(new_n895), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1158), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1156), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n698), .B1(new_n1154), .B2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1149), .B(new_n1164), .C1(new_n1153), .C2(new_n1119), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT119), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1165), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1169));
  AND4_X1   g0969(.A1(KEYINPUT119), .A2(new_n1169), .A3(new_n697), .A4(new_n1167), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1148), .B1(new_n1168), .B2(new_n1170), .ZN(G378));
  NAND2_X1  g0971(.A1(new_n938), .A2(new_n939), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n929), .B1(new_n1124), .B2(new_n916), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1172), .B(G330), .C1(new_n1173), .C2(KEYINPUT40), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n265), .A2(new_n676), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT121), .Z(new_n1176));
  XNOR2_X1  g0976(.A(new_n293), .B(new_n1176), .ZN(new_n1177));
  XOR2_X1   g0977(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1178));
  XNOR2_X1  g0978(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1174), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n940), .A2(G330), .A3(new_n1179), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT122), .ZN(new_n1184));
  OAI21_X1  g0984(.A(KEYINPUT123), .B1(new_n921), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1122), .A2(new_n920), .A3(new_n1125), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1124), .A2(new_n916), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n894), .B1(new_n893), .B2(new_n895), .ZN(new_n1188));
  AOI211_X1 g0988(.A(KEYINPUT104), .B(new_n890), .C1(new_n892), .C2(new_n842), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n862), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1186), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT123), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1192), .A2(KEYINPUT122), .A3(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1183), .A2(new_n1185), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1193), .B1(new_n1192), .B2(KEYINPUT122), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1184), .B(KEYINPUT123), .C1(new_n1186), .C2(new_n1191), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1196), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1156), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1167), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1195), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT57), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1196), .A2(new_n921), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1192), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1203), .B1(new_n1167), .B2(new_n1200), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n698), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1204), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1195), .A2(new_n1199), .A3(new_n748), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n748), .B(new_n697), .C1(new_n801), .C2(new_n837), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n789), .A2(new_n1128), .B1(new_n791), .B2(new_n1136), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n780), .A2(new_n1131), .B1(new_n817), .B2(G137), .ZN(new_n1214));
  INV_X1    g1014(.A(G128), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1214), .B1(new_n1215), .B2(new_n772), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1213), .B(new_n1216), .C1(G150), .C2(new_n796), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT59), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n783), .A2(G159), .ZN(new_n1221));
  AOI211_X1 g1021(.A(G33), .B(G41), .C1(new_n786), .C2(G124), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G41), .B(new_n267), .C1(new_n780), .C2(G77), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n783), .A2(G58), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n786), .A2(G283), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1224), .A2(new_n1026), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n789), .A2(new_n601), .B1(new_n775), .B2(new_n329), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n481), .A2(new_n791), .B1(new_n772), .B2(new_n220), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(KEYINPUT58), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1230), .A2(KEYINPUT58), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n273), .B1(new_n337), .B2(new_n257), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n801), .ZN(new_n1234));
  AND4_X1   g1034(.A1(new_n1223), .A2(new_n1231), .A3(new_n1232), .A4(new_n1234), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1212), .B1(new_n769), .B2(new_n1235), .C1(new_n1179), .C2(new_n763), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1211), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1210), .A2(new_n1238), .ZN(G375));
  NAND2_X1  g1039(.A1(new_n1156), .A2(new_n1163), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1241), .A2(new_n985), .A3(new_n1164), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n816), .B1(new_n202), .B2(new_n837), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(G116), .A2(new_n792), .B1(new_n817), .B2(G107), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n830), .B2(new_n789), .ZN(new_n1245));
  XOR2_X1   g1045(.A(new_n1245), .B(KEYINPUT124), .Z(new_n1246));
  AOI22_X1  g1046(.A1(G283), .A2(new_n803), .B1(new_n786), .B2(G303), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n481), .B2(new_n779), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1248), .A2(new_n267), .A3(new_n1032), .A4(new_n1056), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n779), .A2(new_n358), .B1(new_n785), .B2(new_n1215), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT125), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1225), .B(new_n267), .C1(new_n801), .C2(new_n795), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n789), .A2(new_n1136), .B1(new_n791), .B2(new_n1130), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n772), .A2(new_n819), .B1(new_n775), .B2(new_n254), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1246), .A2(new_n1249), .B1(new_n1251), .B2(new_n1255), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1243), .B1(new_n769), .B2(new_n1256), .C1(new_n1110), .C2(new_n763), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n1163), .B2(new_n747), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1242), .A2(new_n1258), .ZN(G381));
  AOI21_X1  g1059(.A(new_n1237), .B1(new_n1204), .B2(new_n1209), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1169), .A2(new_n697), .A3(new_n1167), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1148), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT126), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1148), .A2(new_n1261), .A3(KEYINPUT126), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1260), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(G390), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1242), .A2(new_n1258), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(G393), .A2(G396), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n850), .A4(new_n1270), .ZN(new_n1271));
  OR3_X1    g1071(.A1(new_n1267), .A2(G387), .A3(new_n1271), .ZN(G407));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G343), .C2(new_n1267), .ZN(G409));
  AOI21_X1  g1073(.A(new_n814), .B1(new_n1040), .B2(new_n1072), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1270), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1012), .A2(new_n748), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n984), .A2(new_n981), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G390), .B(new_n1037), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(G390), .B1(new_n1013), .B2(new_n1037), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1276), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G387), .A2(new_n1268), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(new_n1275), .A3(new_n1279), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1156), .A2(new_n1163), .A3(KEYINPUT60), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1286), .A2(new_n697), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT60), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1240), .B1(new_n1164), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1258), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1290), .A2(G384), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(G384), .ZN(new_n1293));
  INV_X1    g1093(.A(G213), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1294), .A2(G343), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(G2897), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1292), .A2(new_n1293), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1183), .A2(new_n1192), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1206), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n748), .A3(new_n1301), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1236), .B(new_n1302), .C1(new_n1202), .C2(new_n985), .ZN(new_n1303));
  AOI22_X1  g1103(.A1(new_n1260), .A2(G378), .B1(new_n1266), .B2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1299), .B1(new_n1304), .B2(new_n1295), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1210), .A2(G378), .A3(new_n1238), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT126), .B1(new_n1148), .B2(new_n1261), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1265), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1303), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1295), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .A4(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1305), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  AOI211_X1 g1117(.A(new_n1295), .B(new_n1313), .C1(new_n1306), .C2(new_n1309), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1318), .A2(new_n1311), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1285), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1295), .B1(new_n1306), .B2(new_n1309), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1314), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1299), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT63), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1322), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1282), .A2(new_n1316), .A3(new_n1284), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(KEYINPUT127), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT127), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1282), .A2(new_n1284), .A3(new_n1329), .A4(new_n1316), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1331), .B1(new_n1318), .B2(KEYINPUT63), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1326), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1320), .A2(new_n1333), .ZN(G405));
  NAND2_X1  g1134(.A1(G375), .A2(new_n1266), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1306), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1314), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1335), .A2(new_n1306), .A3(new_n1313), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(new_n1339), .B(new_n1285), .ZN(G402));
endmodule


