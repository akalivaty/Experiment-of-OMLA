

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U551 ( .A(n521), .B(KEYINPUT17), .ZN(n539) );
  NOR2_X2 U552 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U553 ( .A(n690), .B(KEYINPUT32), .ZN(n711) );
  BUF_X1 U554 ( .A(n661), .Z(n677) );
  AND2_X1 U555 ( .A1(n539), .A2(G137), .ZN(n522) );
  BUF_X1 U556 ( .A(n539), .Z(n540) );
  AND2_X1 U557 ( .A1(n711), .A2(n692), .ZN(n693) );
  XNOR2_X1 U558 ( .A(n608), .B(n607), .ZN(n610) );
  NOR2_X1 U559 ( .A1(n666), .A2(n665), .ZN(n668) );
  XNOR2_X1 U560 ( .A(n701), .B(n700), .ZN(n706) );
  NAND2_X1 U561 ( .A1(n699), .A2(n519), .ZN(n701) );
  NAND2_X1 U562 ( .A1(n529), .A2(n520), .ZN(n521) );
  XNOR2_X1 U563 ( .A(n526), .B(KEYINPUT23), .ZN(n527) );
  INV_X1 U564 ( .A(KEYINPUT66), .ZN(n526) );
  XOR2_X1 U565 ( .A(n620), .B(KEYINPUT26), .Z(n516) );
  AND2_X1 U566 ( .A1(n998), .A2(n769), .ZN(n517) );
  AND2_X1 U567 ( .A1(n516), .A2(n632), .ZN(n518) );
  AND2_X1 U568 ( .A1(n698), .A2(n697), .ZN(n519) );
  AND2_X1 U569 ( .A1(n653), .A2(G1996), .ZN(n620) );
  INV_X1 U570 ( .A(n981), .ZN(n630) );
  AND2_X1 U571 ( .A1(n631), .A2(n630), .ZN(n632) );
  INV_X1 U572 ( .A(KEYINPUT29), .ZN(n648) );
  NOR2_X1 U573 ( .A1(G2084), .A2(n677), .ZN(n670) );
  NAND2_X1 U574 ( .A1(n673), .A2(n672), .ZN(n674) );
  INV_X1 U575 ( .A(KEYINPUT107), .ZN(n700) );
  INV_X1 U576 ( .A(KEYINPUT108), .ZN(n707) );
  INV_X1 U577 ( .A(G2105), .ZN(n520) );
  NOR2_X1 U578 ( .A1(n756), .A2(n517), .ZN(n757) );
  NOR2_X1 U579 ( .A1(G651), .A2(G543), .ZN(n800) );
  NOR2_X2 U580 ( .A1(n529), .A2(G2105), .ZN(n898) );
  NOR2_X1 U581 ( .A1(G651), .A2(n584), .ZN(n803) );
  BUF_X1 U582 ( .A(n604), .Z(G160) );
  XNOR2_X1 U583 ( .A(n522), .B(KEYINPUT67), .ZN(n524) );
  AND2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n893) );
  NAND2_X1 U585 ( .A1(n893), .A2(G113), .ZN(n523) );
  NAND2_X1 U586 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U587 ( .A(n525), .B(KEYINPUT68), .ZN(n534) );
  INV_X2 U588 ( .A(G2104), .ZN(n529) );
  NAND2_X1 U589 ( .A1(G101), .A2(n898), .ZN(n528) );
  XNOR2_X1 U590 ( .A(n528), .B(n527), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n529), .A2(G2105), .ZN(n530) );
  XNOR2_X2 U592 ( .A(n530), .B(KEYINPUT65), .ZN(n894) );
  NAND2_X1 U593 ( .A1(G125), .A2(n894), .ZN(n531) );
  NAND2_X1 U594 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U595 ( .A(n535), .B(KEYINPUT64), .ZN(n604) );
  NAND2_X1 U596 ( .A1(n893), .A2(G114), .ZN(n538) );
  NAND2_X1 U597 ( .A1(G102), .A2(n898), .ZN(n536) );
  XOR2_X1 U598 ( .A(KEYINPUT87), .B(n536), .Z(n537) );
  NAND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n544) );
  NAND2_X1 U600 ( .A1(G138), .A2(n540), .ZN(n542) );
  NAND2_X1 U601 ( .A1(G126), .A2(n894), .ZN(n541) );
  NAND2_X1 U602 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U603 ( .A1(n544), .A2(n543), .ZN(G164) );
  XOR2_X1 U604 ( .A(G543), .B(KEYINPUT0), .Z(n584) );
  NAND2_X1 U605 ( .A1(G53), .A2(n803), .ZN(n545) );
  XNOR2_X1 U606 ( .A(n545), .B(KEYINPUT72), .ZN(n554) );
  INV_X1 U607 ( .A(G651), .ZN(n549) );
  NOR2_X1 U608 ( .A1(G543), .A2(n549), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT1), .B(n546), .Z(n799) );
  NAND2_X1 U610 ( .A1(G65), .A2(n799), .ZN(n548) );
  NAND2_X1 U611 ( .A1(G91), .A2(n800), .ZN(n547) );
  NAND2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n552) );
  NOR2_X1 U613 ( .A1(n584), .A2(n549), .ZN(n804) );
  NAND2_X1 U614 ( .A1(G78), .A2(n804), .ZN(n550) );
  XNOR2_X1 U615 ( .A(KEYINPUT71), .B(n550), .ZN(n551) );
  NOR2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(G299) );
  NAND2_X1 U618 ( .A1(G90), .A2(n800), .ZN(n556) );
  NAND2_X1 U619 ( .A1(G77), .A2(n804), .ZN(n555) );
  NAND2_X1 U620 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U621 ( .A(KEYINPUT9), .B(n557), .ZN(n561) );
  NAND2_X1 U622 ( .A1(n803), .A2(G52), .ZN(n559) );
  NAND2_X1 U623 ( .A1(G64), .A2(n799), .ZN(n558) );
  AND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(G301) );
  NAND2_X1 U626 ( .A1(n800), .A2(G89), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U628 ( .A1(G76), .A2(n804), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(KEYINPUT5), .B(n565), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n803), .A2(G51), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT75), .B(n566), .Z(n568) );
  NAND2_X1 U633 ( .A1(n799), .A2(G63), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT6), .B(n569), .Z(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(KEYINPUT7), .B(n572), .ZN(G168) );
  NAND2_X1 U638 ( .A1(G88), .A2(n800), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G75), .A2(n804), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n579) );
  NAND2_X1 U641 ( .A1(G62), .A2(n799), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n575), .B(KEYINPUT82), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n803), .A2(G50), .ZN(n576) );
  NAND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(G166) );
  INV_X1 U646 ( .A(G166), .ZN(G303) );
  XOR2_X1 U647 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U648 ( .A1(G651), .A2(G74), .ZN(n580) );
  XOR2_X1 U649 ( .A(KEYINPUT79), .B(n580), .Z(n582) );
  NAND2_X1 U650 ( .A1(n803), .A2(G49), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U652 ( .A(KEYINPUT80), .B(n583), .Z(n586) );
  NAND2_X1 U653 ( .A1(n584), .A2(G87), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U655 ( .A1(n799), .A2(n587), .ZN(n588) );
  XNOR2_X1 U656 ( .A(KEYINPUT81), .B(n588), .ZN(G288) );
  NAND2_X1 U657 ( .A1(G61), .A2(n799), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G86), .A2(n800), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U660 ( .A1(n804), .A2(G73), .ZN(n591) );
  XOR2_X1 U661 ( .A(KEYINPUT2), .B(n591), .Z(n592) );
  NOR2_X1 U662 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n803), .A2(G48), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(G305) );
  NAND2_X1 U665 ( .A1(n803), .A2(G47), .ZN(n596) );
  XOR2_X1 U666 ( .A(KEYINPUT69), .B(n596), .Z(n598) );
  NAND2_X1 U667 ( .A1(n799), .A2(G60), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U669 ( .A(KEYINPUT70), .B(n599), .Z(n603) );
  NAND2_X1 U670 ( .A1(G85), .A2(n800), .ZN(n601) );
  NAND2_X1 U671 ( .A1(G72), .A2(n804), .ZN(n600) );
  AND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n603), .A2(n602), .ZN(G290) );
  NAND2_X1 U674 ( .A1(n604), .A2(G40), .ZN(n735) );
  INV_X1 U675 ( .A(n735), .ZN(n605) );
  NOR2_X1 U676 ( .A1(G164), .A2(G1384), .ZN(n736) );
  NAND2_X2 U677 ( .A1(n605), .A2(n736), .ZN(n661) );
  INV_X1 U678 ( .A(KEYINPUT94), .ZN(n606) );
  XNOR2_X2 U679 ( .A(n661), .B(n606), .ZN(n651) );
  NAND2_X1 U680 ( .A1(n651), .A2(G2067), .ZN(n608) );
  INV_X1 U681 ( .A(KEYINPUT99), .ZN(n607) );
  NAND2_X1 U682 ( .A1(G1348), .A2(n677), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U684 ( .A(n611), .B(KEYINPUT100), .ZN(n634) );
  NAND2_X1 U685 ( .A1(G79), .A2(n804), .ZN(n618) );
  NAND2_X1 U686 ( .A1(G66), .A2(n799), .ZN(n613) );
  NAND2_X1 U687 ( .A1(G92), .A2(n800), .ZN(n612) );
  NAND2_X1 U688 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n803), .A2(G54), .ZN(n614) );
  XOR2_X1 U690 ( .A(KEYINPUT74), .B(n614), .Z(n615) );
  NOR2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n619), .B(KEYINPUT15), .ZN(n918) );
  INV_X1 U694 ( .A(n661), .ZN(n653) );
  NAND2_X1 U695 ( .A1(n677), .A2(G1341), .ZN(n631) );
  NAND2_X1 U696 ( .A1(G56), .A2(n799), .ZN(n621) );
  XOR2_X1 U697 ( .A(KEYINPUT14), .B(n621), .Z(n627) );
  NAND2_X1 U698 ( .A1(n800), .A2(G81), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n622), .B(KEYINPUT12), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G68), .A2(n804), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U702 ( .A(KEYINPUT13), .B(n625), .Z(n626) );
  NOR2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n803), .A2(G43), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n981) );
  NAND2_X1 U706 ( .A1(n918), .A2(n518), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n634), .A2(n633), .ZN(n636) );
  OR2_X1 U708 ( .A1(n918), .A2(n518), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n642) );
  XOR2_X1 U710 ( .A(KEYINPUT97), .B(KEYINPUT27), .Z(n638) );
  NAND2_X1 U711 ( .A1(G2072), .A2(n651), .ZN(n637) );
  XNOR2_X1 U712 ( .A(n638), .B(n637), .ZN(n640) );
  INV_X1 U713 ( .A(G1956), .ZN(n1013) );
  NOR2_X1 U714 ( .A1(n651), .A2(n1013), .ZN(n639) );
  NOR2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n643) );
  INV_X1 U716 ( .A(G299), .ZN(n812) );
  NAND2_X1 U717 ( .A1(n643), .A2(n812), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n642), .A2(n641), .ZN(n647) );
  NOR2_X1 U719 ( .A1(n643), .A2(n812), .ZN(n645) );
  XOR2_X1 U720 ( .A(KEYINPUT28), .B(KEYINPUT98), .Z(n644) );
  XNOR2_X1 U721 ( .A(n645), .B(n644), .ZN(n646) );
  NAND2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n649), .B(n648), .ZN(n658) );
  XNOR2_X1 U724 ( .A(G2078), .B(KEYINPUT25), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n650), .B(KEYINPUT95), .ZN(n960) );
  INV_X1 U726 ( .A(n651), .ZN(n652) );
  NOR2_X1 U727 ( .A1(n960), .A2(n652), .ZN(n655) );
  NOR2_X1 U728 ( .A1(n653), .A2(G1961), .ZN(n654) );
  NOR2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n659) );
  NOR2_X1 U730 ( .A1(n659), .A2(G301), .ZN(n656) );
  XOR2_X1 U731 ( .A(KEYINPUT96), .B(n656), .Z(n657) );
  NAND2_X1 U732 ( .A1(n658), .A2(n657), .ZN(n684) );
  NAND2_X1 U733 ( .A1(n659), .A2(G301), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n660), .B(KEYINPUT101), .ZN(n666) );
  NAND2_X1 U735 ( .A1(G8), .A2(n661), .ZN(n721) );
  NOR2_X1 U736 ( .A1(G1966), .A2(n721), .ZN(n671) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n662) );
  NAND2_X1 U738 ( .A1(G8), .A2(n662), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(KEYINPUT30), .ZN(n664) );
  NOR2_X1 U740 ( .A1(n664), .A2(G168), .ZN(n665) );
  XOR2_X1 U741 ( .A(KEYINPUT102), .B(KEYINPUT31), .Z(n667) );
  XNOR2_X1 U742 ( .A(n668), .B(n667), .ZN(n682) );
  NAND2_X1 U743 ( .A1(n684), .A2(n682), .ZN(n669) );
  XNOR2_X1 U744 ( .A(n669), .B(KEYINPUT103), .ZN(n675) );
  NAND2_X1 U745 ( .A1(G8), .A2(n670), .ZN(n673) );
  INV_X1 U746 ( .A(n671), .ZN(n672) );
  OR2_X2 U747 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U748 ( .A(n676), .B(KEYINPUT104), .ZN(n710) );
  NOR2_X1 U749 ( .A1(G1971), .A2(n721), .ZN(n679) );
  NOR2_X1 U750 ( .A1(G2090), .A2(n677), .ZN(n678) );
  NOR2_X1 U751 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U752 ( .A(KEYINPUT105), .B(n680), .Z(n681) );
  NAND2_X1 U753 ( .A1(n681), .A2(G303), .ZN(n685) );
  AND2_X1 U754 ( .A1(n682), .A2(n685), .ZN(n683) );
  NAND2_X1 U755 ( .A1(n684), .A2(n683), .ZN(n688) );
  INV_X1 U756 ( .A(n685), .ZN(n686) );
  OR2_X1 U757 ( .A1(n686), .A2(G286), .ZN(n687) );
  AND2_X1 U758 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U759 ( .A1(n689), .A2(G8), .ZN(n690) );
  NAND2_X1 U760 ( .A1(G1976), .A2(G288), .ZN(n992) );
  INV_X1 U761 ( .A(n721), .ZN(n691) );
  NAND2_X1 U762 ( .A1(n992), .A2(n691), .ZN(n696) );
  INV_X1 U763 ( .A(n696), .ZN(n692) );
  NAND2_X1 U764 ( .A1(n710), .A2(n693), .ZN(n699) );
  NOR2_X1 U765 ( .A1(G288), .A2(G1976), .ZN(n694) );
  XNOR2_X1 U766 ( .A(n694), .B(KEYINPUT106), .ZN(n702) );
  NOR2_X1 U767 ( .A1(G1971), .A2(G303), .ZN(n695) );
  NOR2_X1 U768 ( .A1(n702), .A2(n695), .ZN(n993) );
  OR2_X1 U769 ( .A1(n696), .A2(n993), .ZN(n698) );
  INV_X1 U770 ( .A(KEYINPUT33), .ZN(n697) );
  INV_X1 U771 ( .A(n702), .ZN(n703) );
  NOR2_X1 U772 ( .A1(n721), .A2(n703), .ZN(n704) );
  NAND2_X1 U773 ( .A1(KEYINPUT33), .A2(n704), .ZN(n705) );
  NAND2_X1 U774 ( .A1(n706), .A2(n705), .ZN(n708) );
  XNOR2_X1 U775 ( .A(n708), .B(n707), .ZN(n709) );
  XOR2_X1 U776 ( .A(G1981), .B(G305), .Z(n986) );
  NAND2_X1 U777 ( .A1(n709), .A2(n986), .ZN(n717) );
  NAND2_X1 U778 ( .A1(n710), .A2(n711), .ZN(n714) );
  NOR2_X1 U779 ( .A1(G2090), .A2(G303), .ZN(n712) );
  NAND2_X1 U780 ( .A1(G8), .A2(n712), .ZN(n713) );
  NAND2_X1 U781 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U782 ( .A1(n715), .A2(n721), .ZN(n716) );
  NAND2_X1 U783 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U784 ( .A(n718), .B(KEYINPUT109), .ZN(n723) );
  NOR2_X1 U785 ( .A1(G1981), .A2(G305), .ZN(n719) );
  XOR2_X1 U786 ( .A(n719), .B(KEYINPUT24), .Z(n720) );
  OR2_X1 U787 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U788 ( .A1(n723), .A2(n722), .ZN(n758) );
  XNOR2_X1 U789 ( .A(G2067), .B(KEYINPUT37), .ZN(n724) );
  XNOR2_X1 U790 ( .A(n724), .B(KEYINPUT88), .ZN(n767) );
  NAND2_X1 U791 ( .A1(G104), .A2(n898), .ZN(n726) );
  NAND2_X1 U792 ( .A1(G140), .A2(n540), .ZN(n725) );
  NAND2_X1 U793 ( .A1(n726), .A2(n725), .ZN(n728) );
  XOR2_X1 U794 ( .A(KEYINPUT89), .B(KEYINPUT34), .Z(n727) );
  XNOR2_X1 U795 ( .A(n728), .B(n727), .ZN(n733) );
  NAND2_X1 U796 ( .A1(G116), .A2(n893), .ZN(n730) );
  NAND2_X1 U797 ( .A1(G128), .A2(n894), .ZN(n729) );
  NAND2_X1 U798 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U799 ( .A(KEYINPUT35), .B(n731), .Z(n732) );
  NOR2_X1 U800 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U801 ( .A(KEYINPUT36), .B(n734), .ZN(n906) );
  NOR2_X1 U802 ( .A1(n767), .A2(n906), .ZN(n939) );
  NOR2_X1 U803 ( .A1(n736), .A2(n735), .ZN(n769) );
  NAND2_X1 U804 ( .A1(n939), .A2(n769), .ZN(n737) );
  XNOR2_X1 U805 ( .A(n737), .B(KEYINPUT90), .ZN(n765) );
  XOR2_X1 U806 ( .A(KEYINPUT92), .B(KEYINPUT38), .Z(n739) );
  NAND2_X1 U807 ( .A1(G105), .A2(n898), .ZN(n738) );
  XNOR2_X1 U808 ( .A(n739), .B(n738), .ZN(n743) );
  NAND2_X1 U809 ( .A1(G117), .A2(n893), .ZN(n741) );
  NAND2_X1 U810 ( .A1(G129), .A2(n894), .ZN(n740) );
  NAND2_X1 U811 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U812 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U813 ( .A(KEYINPUT93), .B(n744), .Z(n746) );
  NAND2_X1 U814 ( .A1(n540), .A2(G141), .ZN(n745) );
  NAND2_X1 U815 ( .A1(n746), .A2(n745), .ZN(n908) );
  NAND2_X1 U816 ( .A1(n908), .A2(G1996), .ZN(n755) );
  NAND2_X1 U817 ( .A1(G107), .A2(n893), .ZN(n748) );
  NAND2_X1 U818 ( .A1(G119), .A2(n894), .ZN(n747) );
  NAND2_X1 U819 ( .A1(n748), .A2(n747), .ZN(n751) );
  NAND2_X1 U820 ( .A1(G95), .A2(n898), .ZN(n749) );
  XNOR2_X1 U821 ( .A(KEYINPUT91), .B(n749), .ZN(n750) );
  NOR2_X1 U822 ( .A1(n751), .A2(n750), .ZN(n753) );
  NAND2_X1 U823 ( .A1(n540), .A2(G131), .ZN(n752) );
  NAND2_X1 U824 ( .A1(n753), .A2(n752), .ZN(n890) );
  NAND2_X1 U825 ( .A1(n890), .A2(G1991), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n755), .A2(n754), .ZN(n933) );
  NAND2_X1 U827 ( .A1(n933), .A2(n769), .ZN(n759) );
  NAND2_X1 U828 ( .A1(n765), .A2(n759), .ZN(n756) );
  XNOR2_X1 U829 ( .A(G1986), .B(G290), .ZN(n998) );
  NAND2_X1 U830 ( .A1(n758), .A2(n757), .ZN(n772) );
  NOR2_X1 U831 ( .A1(G1996), .A2(n908), .ZN(n931) );
  INV_X1 U832 ( .A(n759), .ZN(n762) );
  NOR2_X1 U833 ( .A1(G1991), .A2(n890), .ZN(n935) );
  NOR2_X1 U834 ( .A1(G1986), .A2(G290), .ZN(n760) );
  NOR2_X1 U835 ( .A1(n935), .A2(n760), .ZN(n761) );
  NOR2_X1 U836 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U837 ( .A1(n931), .A2(n763), .ZN(n764) );
  XNOR2_X1 U838 ( .A(KEYINPUT39), .B(n764), .ZN(n766) );
  NAND2_X1 U839 ( .A1(n766), .A2(n765), .ZN(n768) );
  NAND2_X1 U840 ( .A1(n767), .A2(n906), .ZN(n940) );
  NAND2_X1 U841 ( .A1(n768), .A2(n940), .ZN(n770) );
  NAND2_X1 U842 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U843 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U844 ( .A(n773), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U845 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U846 ( .A(G132), .ZN(G219) );
  INV_X1 U847 ( .A(G82), .ZN(G220) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n774) );
  XNOR2_X1 U849 ( .A(n774), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U850 ( .A(G223), .ZN(n851) );
  NAND2_X1 U851 ( .A1(n851), .A2(G567), .ZN(n775) );
  XOR2_X1 U852 ( .A(KEYINPUT11), .B(n775), .Z(G234) );
  INV_X1 U853 ( .A(G860), .ZN(n780) );
  OR2_X1 U854 ( .A1(n981), .A2(n780), .ZN(G153) );
  NAND2_X1 U855 ( .A1(G868), .A2(G301), .ZN(n777) );
  INV_X1 U856 ( .A(n918), .ZN(n978) );
  INV_X1 U857 ( .A(G868), .ZN(n820) );
  NAND2_X1 U858 ( .A1(n978), .A2(n820), .ZN(n776) );
  NAND2_X1 U859 ( .A1(n777), .A2(n776), .ZN(G284) );
  NOR2_X1 U860 ( .A1(G286), .A2(n820), .ZN(n779) );
  NOR2_X1 U861 ( .A1(G868), .A2(G299), .ZN(n778) );
  NOR2_X1 U862 ( .A1(n779), .A2(n778), .ZN(G297) );
  NAND2_X1 U863 ( .A1(n780), .A2(G559), .ZN(n781) );
  NAND2_X1 U864 ( .A1(n781), .A2(n918), .ZN(n782) );
  XNOR2_X1 U865 ( .A(n782), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U866 ( .A1(G868), .A2(n981), .ZN(n785) );
  NAND2_X1 U867 ( .A1(G868), .A2(n918), .ZN(n783) );
  NOR2_X1 U868 ( .A1(G559), .A2(n783), .ZN(n784) );
  NOR2_X1 U869 ( .A1(n785), .A2(n784), .ZN(G282) );
  NAND2_X1 U870 ( .A1(G99), .A2(n898), .ZN(n787) );
  NAND2_X1 U871 ( .A1(G111), .A2(n893), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n793) );
  NAND2_X1 U873 ( .A1(G123), .A2(n894), .ZN(n788) );
  XNOR2_X1 U874 ( .A(n788), .B(KEYINPUT76), .ZN(n789) );
  XNOR2_X1 U875 ( .A(n789), .B(KEYINPUT18), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G135), .A2(n540), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U878 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U879 ( .A(KEYINPUT77), .B(n794), .Z(n934) );
  XNOR2_X1 U880 ( .A(n934), .B(G2096), .ZN(n795) );
  XNOR2_X1 U881 ( .A(n795), .B(KEYINPUT78), .ZN(n797) );
  INV_X1 U882 ( .A(G2100), .ZN(n796) );
  NAND2_X1 U883 ( .A1(n797), .A2(n796), .ZN(G156) );
  NAND2_X1 U884 ( .A1(n918), .A2(G559), .ZN(n818) );
  XNOR2_X1 U885 ( .A(n981), .B(n818), .ZN(n798) );
  NOR2_X1 U886 ( .A1(n798), .A2(G860), .ZN(n809) );
  NAND2_X1 U887 ( .A1(G67), .A2(n799), .ZN(n802) );
  NAND2_X1 U888 ( .A1(G93), .A2(n800), .ZN(n801) );
  NAND2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n808) );
  NAND2_X1 U890 ( .A1(G55), .A2(n803), .ZN(n806) );
  NAND2_X1 U891 ( .A1(G80), .A2(n804), .ZN(n805) );
  NAND2_X1 U892 ( .A1(n806), .A2(n805), .ZN(n807) );
  OR2_X1 U893 ( .A1(n808), .A2(n807), .ZN(n821) );
  XOR2_X1 U894 ( .A(n809), .B(n821), .Z(G145) );
  XNOR2_X1 U895 ( .A(KEYINPUT19), .B(KEYINPUT83), .ZN(n810) );
  XOR2_X1 U896 ( .A(n810), .B(n821), .Z(n811) );
  XNOR2_X1 U897 ( .A(n812), .B(n811), .ZN(n815) );
  XNOR2_X1 U898 ( .A(G166), .B(G305), .ZN(n813) );
  XNOR2_X1 U899 ( .A(n813), .B(n981), .ZN(n814) );
  XNOR2_X1 U900 ( .A(n815), .B(n814), .ZN(n816) );
  XNOR2_X1 U901 ( .A(n816), .B(G290), .ZN(n817) );
  XNOR2_X1 U902 ( .A(n817), .B(G288), .ZN(n915) );
  XOR2_X1 U903 ( .A(n915), .B(n818), .Z(n819) );
  NAND2_X1 U904 ( .A1(G868), .A2(n819), .ZN(n823) );
  NAND2_X1 U905 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U906 ( .A1(n823), .A2(n822), .ZN(G295) );
  NAND2_X1 U907 ( .A1(G2084), .A2(G2078), .ZN(n825) );
  XOR2_X1 U908 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n824) );
  XNOR2_X1 U909 ( .A(n825), .B(n824), .ZN(n826) );
  NAND2_X1 U910 ( .A1(G2090), .A2(n826), .ZN(n827) );
  XNOR2_X1 U911 ( .A(KEYINPUT21), .B(n827), .ZN(n828) );
  NAND2_X1 U912 ( .A1(n828), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U913 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U914 ( .A(KEYINPUT73), .B(G57), .ZN(G237) );
  NOR2_X1 U915 ( .A1(G220), .A2(G219), .ZN(n829) );
  XOR2_X1 U916 ( .A(KEYINPUT22), .B(n829), .Z(n830) );
  NOR2_X1 U917 ( .A1(G218), .A2(n830), .ZN(n831) );
  XOR2_X1 U918 ( .A(KEYINPUT85), .B(n831), .Z(n832) );
  NAND2_X1 U919 ( .A1(G96), .A2(n832), .ZN(n857) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n857), .ZN(n837) );
  NAND2_X1 U921 ( .A1(G69), .A2(G120), .ZN(n833) );
  XNOR2_X1 U922 ( .A(KEYINPUT86), .B(n833), .ZN(n834) );
  NOR2_X1 U923 ( .A1(G237), .A2(n834), .ZN(n835) );
  NAND2_X1 U924 ( .A1(G108), .A2(n835), .ZN(n856) );
  NAND2_X1 U925 ( .A1(G567), .A2(n856), .ZN(n836) );
  NAND2_X1 U926 ( .A1(n837), .A2(n836), .ZN(n858) );
  NAND2_X1 U927 ( .A1(G483), .A2(G661), .ZN(n838) );
  NOR2_X1 U928 ( .A1(n858), .A2(n838), .ZN(n854) );
  NAND2_X1 U929 ( .A1(n854), .A2(G36), .ZN(G176) );
  XNOR2_X1 U930 ( .A(G1341), .B(G1348), .ZN(n839) );
  XNOR2_X1 U931 ( .A(n839), .B(G2443), .ZN(n849) );
  XOR2_X1 U932 ( .A(KEYINPUT112), .B(G2430), .Z(n841) );
  XNOR2_X1 U933 ( .A(G2454), .B(G2438), .ZN(n840) );
  XNOR2_X1 U934 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U935 ( .A(G2446), .B(KEYINPUT111), .Z(n843) );
  XNOR2_X1 U936 ( .A(G2451), .B(G2427), .ZN(n842) );
  XNOR2_X1 U937 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U938 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U939 ( .A(G2435), .B(KEYINPUT110), .ZN(n846) );
  XNOR2_X1 U940 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U941 ( .A(n849), .B(n848), .ZN(n850) );
  NAND2_X1 U942 ( .A1(n850), .A2(G14), .ZN(n921) );
  XNOR2_X1 U943 ( .A(KEYINPUT113), .B(n921), .ZN(G401) );
  NAND2_X1 U944 ( .A1(G2106), .A2(n851), .ZN(G217) );
  AND2_X1 U945 ( .A1(G15), .A2(G2), .ZN(n852) );
  NAND2_X1 U946 ( .A1(G661), .A2(n852), .ZN(G259) );
  NAND2_X1 U947 ( .A1(G3), .A2(G1), .ZN(n853) );
  XNOR2_X1 U948 ( .A(KEYINPUT114), .B(n853), .ZN(n855) );
  NAND2_X1 U949 ( .A1(n855), .A2(n854), .ZN(G188) );
  XNOR2_X1 U950 ( .A(G120), .B(KEYINPUT115), .ZN(G236) );
  INV_X1 U952 ( .A(G108), .ZN(G238) );
  INV_X1 U953 ( .A(G96), .ZN(G221) );
  INV_X1 U954 ( .A(G69), .ZN(G235) );
  NOR2_X1 U955 ( .A1(n857), .A2(n856), .ZN(G325) );
  INV_X1 U956 ( .A(G325), .ZN(G261) );
  INV_X1 U957 ( .A(n858), .ZN(G319) );
  XOR2_X1 U958 ( .A(G2100), .B(G2096), .Z(n860) );
  XNOR2_X1 U959 ( .A(KEYINPUT42), .B(G2678), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U961 ( .A(KEYINPUT43), .B(G2090), .Z(n862) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2072), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U964 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U965 ( .A(G2084), .B(G2078), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(G227) );
  XOR2_X1 U967 ( .A(G1956), .B(G1971), .Z(n868) );
  XNOR2_X1 U968 ( .A(G1986), .B(G1976), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U970 ( .A(n869), .B(KEYINPUT41), .Z(n871) );
  XNOR2_X1 U971 ( .A(G1996), .B(G1991), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U973 ( .A(G2474), .B(G1961), .Z(n873) );
  XNOR2_X1 U974 ( .A(G1981), .B(G1966), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(G229) );
  NAND2_X1 U977 ( .A1(G100), .A2(n898), .ZN(n877) );
  NAND2_X1 U978 ( .A1(G112), .A2(n893), .ZN(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G124), .A2(n894), .ZN(n878) );
  XNOR2_X1 U981 ( .A(n878), .B(KEYINPUT44), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n540), .A2(G136), .ZN(n879) );
  NAND2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U984 ( .A1(n882), .A2(n881), .ZN(G162) );
  XNOR2_X1 U985 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n892) );
  NAND2_X1 U986 ( .A1(G103), .A2(n898), .ZN(n884) );
  NAND2_X1 U987 ( .A1(G139), .A2(n540), .ZN(n883) );
  NAND2_X1 U988 ( .A1(n884), .A2(n883), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G115), .A2(n893), .ZN(n886) );
  NAND2_X1 U990 ( .A1(G127), .A2(n894), .ZN(n885) );
  NAND2_X1 U991 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n887), .Z(n888) );
  NOR2_X1 U993 ( .A1(n889), .A2(n888), .ZN(n946) );
  XNOR2_X1 U994 ( .A(n890), .B(n946), .ZN(n891) );
  XNOR2_X1 U995 ( .A(n892), .B(n891), .ZN(n905) );
  NAND2_X1 U996 ( .A1(G118), .A2(n893), .ZN(n896) );
  NAND2_X1 U997 ( .A1(G130), .A2(n894), .ZN(n895) );
  NAND2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n903) );
  NAND2_X1 U999 ( .A1(n540), .A2(G142), .ZN(n897) );
  XNOR2_X1 U1000 ( .A(n897), .B(KEYINPUT116), .ZN(n900) );
  NAND2_X1 U1001 ( .A1(G106), .A2(n898), .ZN(n899) );
  NAND2_X1 U1002 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1003 ( .A(n901), .B(KEYINPUT45), .Z(n902) );
  NOR2_X1 U1004 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1005 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U1006 ( .A(n907), .B(n906), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1008 ( .A(n910), .B(n934), .Z(n912) );
  XNOR2_X1 U1009 ( .A(G164), .B(G162), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(G160), .B(n913), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n914), .ZN(G395) );
  INV_X1 U1013 ( .A(G301), .ZN(G171) );
  XOR2_X1 U1014 ( .A(KEYINPUT117), .B(n915), .Z(n917) );
  XNOR2_X1 U1015 ( .A(G171), .B(G286), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(n917), .B(n916), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n920), .ZN(G397) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n921), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(KEYINPUT118), .B(n922), .ZN(n926) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n923) );
  XOR2_X1 U1022 ( .A(KEYINPUT119), .B(n923), .Z(n924) );
  XNOR2_X1 U1023 ( .A(n924), .B(KEYINPUT49), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(KEYINPUT120), .B(n927), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(G395), .A2(G397), .ZN(n928) );
  NAND2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1028 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1031 ( .A(KEYINPUT51), .B(n932), .Z(n945) );
  INV_X1 U1032 ( .A(n933), .ZN(n937) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n943) );
  XOR2_X1 U1037 ( .A(G160), .B(G2084), .Z(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n952) );
  XOR2_X1 U1040 ( .A(G2072), .B(n946), .Z(n948) );
  XOR2_X1 U1041 ( .A(G164), .B(G2078), .Z(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(n949), .B(KEYINPUT121), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(n950), .B(KEYINPUT50), .ZN(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(KEYINPUT52), .B(n953), .ZN(n954) );
  XOR2_X1 U1047 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n974) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n974), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n955), .A2(G29), .ZN(n956) );
  XOR2_X1 U1050 ( .A(KEYINPUT123), .B(n956), .Z(n1033) );
  XOR2_X1 U1051 ( .A(G1991), .B(G25), .Z(n957) );
  NAND2_X1 U1052 ( .A1(n957), .A2(G28), .ZN(n966) );
  XNOR2_X1 U1053 ( .A(G2067), .B(G26), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(G33), .B(G2072), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(G1996), .B(G32), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(G27), .B(n960), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1061 ( .A(KEYINPUT53), .B(n967), .Z(n970) );
  XOR2_X1 U1062 ( .A(G34), .B(KEYINPUT54), .Z(n968) );
  XNOR2_X1 U1063 ( .A(G2084), .B(n968), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(G35), .B(G2090), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1067 ( .A(n974), .B(n973), .Z(n976) );
  INV_X1 U1068 ( .A(G29), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n977), .A2(G11), .ZN(n1031) );
  XNOR2_X1 U1071 ( .A(G16), .B(KEYINPUT56), .ZN(n1002) );
  XNOR2_X1 U1072 ( .A(G301), .B(G1961), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(n978), .B(G1348), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(G299), .B(G1956), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(n981), .B(G1341), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G168), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(n988), .B(KEYINPUT124), .ZN(n989) );
  XOR2_X1 U1082 ( .A(KEYINPUT57), .B(n989), .Z(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n1000) );
  AND2_X1 U1084 ( .A1(G303), .A2(G1971), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(KEYINPUT125), .B(n996), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1029) );
  INV_X1 U1091 ( .A(G16), .ZN(n1027) );
  XNOR2_X1 U1092 ( .A(G1986), .B(G24), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(G1976), .B(G23), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G22), .B(G1971), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(KEYINPUT127), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(KEYINPUT58), .B(n1008), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G1966), .B(G21), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(G5), .B(G1961), .ZN(n1009) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1024) );
  XNOR2_X1 U1103 ( .A(G20), .B(n1013), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(G1981), .B(G6), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(G19), .B(G1341), .ZN(n1014) );
  NOR2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  XOR2_X1 U1108 ( .A(KEYINPUT59), .B(G1348), .Z(n1018) );
  XNOR2_X1 U1109 ( .A(G4), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1111 ( .A(KEYINPUT126), .B(n1021), .Z(n1022) );
  XNOR2_X1 U1112 ( .A(KEYINPUT60), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1114 ( .A(KEYINPUT61), .B(n1025), .ZN(n1026) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1034), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

