

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735;

  XNOR2_X1 U363 ( .A(n512), .B(G134), .ZN(n519) );
  XNOR2_X1 U364 ( .A(n519), .B(n398), .ZN(n717) );
  INV_X1 U365 ( .A(G953), .ZN(n719) );
  XOR2_X1 U366 ( .A(KEYINPUT31), .B(n613), .Z(n688) );
  XNOR2_X2 U367 ( .A(G128), .B(KEYINPUT82), .ZN(n481) );
  XNOR2_X2 U368 ( .A(n463), .B(n352), .ZN(n571) );
  OR2_X2 U369 ( .A1(n693), .A2(n532), .ZN(n463) );
  AND2_X1 U370 ( .A1(n614), .A2(n648), .ZN(n613) );
  XNOR2_X1 U371 ( .A(n595), .B(KEYINPUT0), .ZN(n614) );
  NOR2_X1 U372 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U373 ( .A(n646), .B(n424), .ZN(n608) );
  NAND2_X1 U374 ( .A1(n456), .A2(n457), .ZN(n646) );
  XNOR2_X1 U375 ( .A(n534), .B(KEYINPUT25), .ZN(n535) );
  XNOR2_X1 U376 ( .A(n477), .B(KEYINPUT65), .ZN(n518) );
  XNOR2_X1 U377 ( .A(G146), .B(KEYINPUT4), .ZN(n477) );
  XNOR2_X1 U378 ( .A(G119), .B(G110), .ZN(n523) );
  BUF_X1 U379 ( .A(n658), .Z(n340) );
  XNOR2_X1 U380 ( .A(n442), .B(n455), .ZN(n341) );
  XNOR2_X1 U381 ( .A(n604), .B(KEYINPUT33), .ZN(n658) );
  XNOR2_X1 U382 ( .A(n442), .B(n455), .ZN(n707) );
  XOR2_X1 U383 ( .A(KEYINPUT68), .B(G101), .Z(n520) );
  XNOR2_X1 U384 ( .A(n717), .B(n520), .ZN(n429) );
  NOR2_X1 U385 ( .A1(n618), .A2(n682), .ZN(n585) );
  XNOR2_X1 U386 ( .A(n518), .B(G131), .ZN(n398) );
  INV_X1 U387 ( .A(n443), .ZN(n600) );
  XNOR2_X1 U388 ( .A(n646), .B(KEYINPUT105), .ZN(n564) );
  NOR2_X1 U389 ( .A1(G902), .A2(n696), .ZN(n549) );
  XNOR2_X1 U390 ( .A(n535), .B(n531), .ZN(n440) );
  XNOR2_X1 U391 ( .A(n489), .B(n397), .ZN(n547) );
  INV_X1 U392 ( .A(G107), .ZN(n397) );
  INV_X1 U393 ( .A(KEYINPUT45), .ZN(n455) );
  NAND2_X1 U394 ( .A1(n372), .A2(n453), .ZN(n718) );
  AND2_X1 U395 ( .A1(n727), .A2(n454), .ZN(n453) );
  XNOR2_X1 U396 ( .A(n373), .B(n363), .ZN(n372) );
  INV_X1 U397 ( .A(n691), .ZN(n454) );
  INV_X1 U398 ( .A(n707), .ZN(n412) );
  XNOR2_X1 U399 ( .A(n438), .B(n480), .ZN(n484) );
  NOR2_X1 U400 ( .A1(n571), .A2(n629), .ZN(n422) );
  OR2_X1 U401 ( .A1(n564), .A2(n343), .ZN(n378) );
  XNOR2_X1 U402 ( .A(G137), .B(KEYINPUT5), .ZN(n513) );
  NOR2_X1 U403 ( .A1(G953), .A2(G237), .ZN(n515) );
  XNOR2_X1 U404 ( .A(n625), .B(KEYINPUT69), .ZN(n627) );
  NOR2_X1 U405 ( .A1(n731), .A2(KEYINPUT44), .ZN(n625) );
  NAND2_X1 U406 ( .A1(n353), .A2(n374), .ZN(n373) );
  XNOR2_X1 U407 ( .A(n419), .B(n358), .ZN(n374) );
  AND2_X1 U408 ( .A1(n345), .A2(n608), .ZN(n572) );
  XNOR2_X1 U409 ( .A(n404), .B(n464), .ZN(n371) );
  XNOR2_X1 U410 ( .A(n465), .B(KEYINPUT91), .ZN(n464) );
  XNOR2_X1 U411 ( .A(n485), .B(n466), .ZN(n404) );
  INV_X1 U412 ( .A(G113), .ZN(n465) );
  XOR2_X1 U413 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n487) );
  XNOR2_X1 U414 ( .A(n429), .B(n394), .ZN(n696) );
  XNOR2_X1 U415 ( .A(n548), .B(n395), .ZN(n394) );
  XNOR2_X1 U416 ( .A(n547), .B(n396), .ZN(n395) );
  NAND2_X1 U417 ( .A1(n391), .A2(n388), .ZN(n562) );
  AND2_X1 U418 ( .A1(n393), .A2(n392), .ZN(n391) );
  NAND2_X1 U419 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U420 ( .A1(n562), .A2(KEYINPUT40), .ZN(n387) );
  XNOR2_X1 U421 ( .A(n572), .B(KEYINPUT110), .ZN(n423) );
  AND2_X1 U422 ( .A1(n596), .A2(n408), .ZN(n407) );
  INV_X1 U423 ( .A(n608), .ZN(n408) );
  XNOR2_X1 U424 ( .A(n422), .B(KEYINPUT19), .ZN(n594) );
  AND2_X1 U425 ( .A1(n458), .A2(n461), .ZN(n457) );
  NAND2_X1 U426 ( .A1(n521), .A2(n460), .ZN(n459) );
  BUF_X1 U427 ( .A(n637), .Z(n443) );
  XNOR2_X1 U428 ( .A(n467), .B(n356), .ZN(n607) );
  NAND2_X1 U429 ( .A1(n614), .A2(n468), .ZN(n467) );
  AND2_X1 U430 ( .A1(n630), .A2(n346), .ZN(n468) );
  NAND2_X1 U431 ( .A1(n412), .A2(n411), .ZN(n410) );
  AND2_X1 U432 ( .A1(n415), .A2(n414), .ZN(n413) );
  NOR2_X1 U433 ( .A1(n718), .A2(KEYINPUT2), .ZN(n411) );
  XNOR2_X1 U434 ( .A(n451), .B(n510), .ZN(n698) );
  XOR2_X1 U435 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n509) );
  INV_X1 U436 ( .A(KEYINPUT123), .ZN(n474) );
  NOR2_X1 U437 ( .A1(n476), .A2(n659), .ZN(n660) );
  XNOR2_X1 U438 ( .A(n447), .B(n446), .ZN(n420) );
  INV_X1 U439 ( .A(KEYINPUT84), .ZN(n446) );
  NAND2_X1 U440 ( .A1(n584), .A2(n681), .ZN(n447) );
  XNOR2_X1 U441 ( .A(n450), .B(KEYINPUT104), .ZN(n632) );
  XNOR2_X1 U442 ( .A(G116), .B(KEYINPUT73), .ZN(n466) );
  XNOR2_X1 U443 ( .A(G119), .B(KEYINPUT3), .ZN(n485) );
  INV_X1 U444 ( .A(KEYINPUT86), .ZN(n587) );
  XOR2_X1 U445 ( .A(G122), .B(G104), .Z(n500) );
  XNOR2_X1 U446 ( .A(G113), .B(G146), .ZN(n499) );
  XOR2_X1 U447 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n493) );
  XNOR2_X1 U448 ( .A(G131), .B(G143), .ZN(n494) );
  XOR2_X1 U449 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n495) );
  INV_X1 U450 ( .A(G140), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n518), .B(n439), .ZN(n438) );
  INV_X1 U452 ( .A(KEYINPUT17), .ZN(n439) );
  INV_X1 U453 ( .A(KEYINPUT18), .ZN(n478) );
  NOR2_X1 U454 ( .A1(n376), .A2(n375), .ZN(n560) );
  AND2_X1 U455 ( .A1(n564), .A2(KEYINPUT30), .ZN(n375) );
  NAND2_X1 U456 ( .A1(n378), .A2(n351), .ZN(n376) );
  NOR2_X1 U457 ( .A1(G902), .A2(G237), .ZN(n491) );
  INV_X1 U458 ( .A(n561), .ZN(n581) );
  INV_X1 U459 ( .A(G902), .ZN(n460) );
  NAND2_X1 U460 ( .A1(n462), .A2(G902), .ZN(n461) );
  XNOR2_X1 U461 ( .A(n371), .B(n514), .ZN(n517) );
  XNOR2_X1 U462 ( .A(n449), .B(n448), .ZN(n522) );
  INV_X1 U463 ( .A(KEYINPUT8), .ZN(n448) );
  NAND2_X1 U464 ( .A1(n719), .A2(G234), .ZN(n449) );
  XNOR2_X1 U465 ( .A(G116), .B(G107), .ZN(n506) );
  XOR2_X1 U466 ( .A(KEYINPUT102), .B(G122), .Z(n507) );
  INV_X1 U467 ( .A(KEYINPUT83), .ZN(n416) );
  XNOR2_X1 U468 ( .A(n426), .B(n425), .ZN(n561) );
  INV_X1 U469 ( .A(G478), .ZN(n425) );
  OR2_X1 U470 ( .A1(n698), .A2(G902), .ZN(n426) );
  INV_X1 U471 ( .A(KEYINPUT6), .ZN(n424) );
  XNOR2_X1 U472 ( .A(n488), .B(n547), .ZN(n405) );
  XNOR2_X1 U473 ( .A(G122), .B(KEYINPUT16), .ZN(n486) );
  NAND2_X1 U474 ( .A1(n385), .A2(n384), .ZN(n383) );
  AND2_X1 U475 ( .A1(n441), .A2(n563), .ZN(n384) );
  AND2_X1 U476 ( .A1(n423), .A2(n422), .ZN(n573) );
  XNOR2_X1 U477 ( .A(n599), .B(n598), .ZN(n733) );
  NOR2_X1 U478 ( .A1(n582), .A2(n561), .ZN(n687) );
  NAND2_X1 U479 ( .A1(n578), .A2(n577), .ZN(n682) );
  NAND2_X1 U480 ( .A1(n607), .A2(n609), .ZN(n601) );
  XNOR2_X1 U481 ( .A(n379), .B(n368), .ZN(G57) );
  XNOR2_X1 U482 ( .A(n382), .B(n357), .ZN(n381) );
  XNOR2_X1 U483 ( .A(n475), .B(n473), .ZN(n699) );
  XNOR2_X1 U484 ( .A(n698), .B(n474), .ZN(n473) );
  INV_X1 U485 ( .A(KEYINPUT122), .ZN(n435) );
  INV_X1 U486 ( .A(KEYINPUT56), .ZN(n433) );
  INV_X1 U487 ( .A(KEYINPUT53), .ZN(n399) );
  OR2_X1 U488 ( .A1(n701), .A2(G902), .ZN(n342) );
  OR2_X1 U489 ( .A1(n629), .A2(KEYINPUT30), .ZN(n343) );
  AND2_X1 U490 ( .A1(n387), .A2(n386), .ZN(n344) );
  INV_X1 U491 ( .A(n683), .ZN(n441) );
  AND2_X1 U492 ( .A1(n565), .A2(n441), .ZN(n345) );
  XOR2_X1 U493 ( .A(KEYINPUT21), .B(n537), .Z(n346) );
  XOR2_X1 U494 ( .A(n517), .B(n516), .Z(n347) );
  XOR2_X1 U495 ( .A(n523), .B(KEYINPUT96), .Z(n348) );
  XOR2_X1 U496 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n349) );
  OR2_X2 U497 ( .A1(n627), .A2(n626), .ZN(n350) );
  AND2_X1 U498 ( .A1(n377), .A2(n557), .ZN(n351) );
  NAND2_X1 U499 ( .A1(G210), .A2(n550), .ZN(n352) );
  AND2_X1 U500 ( .A1(n420), .A2(n421), .ZN(n353) );
  AND2_X1 U501 ( .A1(n586), .A2(n585), .ZN(n354) );
  XOR2_X1 U502 ( .A(KEYINPUT74), .B(KEYINPUT39), .Z(n355) );
  XOR2_X1 U503 ( .A(KEYINPUT22), .B(KEYINPUT76), .Z(n356) );
  XOR2_X1 U504 ( .A(n667), .B(n666), .Z(n357) );
  INV_X1 U505 ( .A(n532), .ZN(n661) );
  XOR2_X1 U506 ( .A(KEYINPUT46), .B(KEYINPUT64), .Z(n358) );
  XOR2_X1 U507 ( .A(KEYINPUT85), .B(KEYINPUT35), .Z(n359) );
  XOR2_X1 U508 ( .A(n693), .B(n692), .Z(n360) );
  XNOR2_X1 U509 ( .A(n662), .B(KEYINPUT59), .ZN(n361) );
  XOR2_X1 U510 ( .A(n696), .B(n695), .Z(n362) );
  XNOR2_X1 U511 ( .A(n587), .B(KEYINPUT48), .ZN(n363) );
  AND2_X1 U512 ( .A1(n532), .A2(G472), .ZN(n364) );
  AND2_X1 U513 ( .A1(n532), .A2(G475), .ZN(n365) );
  AND2_X1 U514 ( .A1(n532), .A2(G210), .ZN(n366) );
  AND2_X1 U515 ( .A1(n532), .A2(G469), .ZN(n367) );
  INV_X1 U516 ( .A(n703), .ZN(n380) );
  XNOR2_X1 U517 ( .A(KEYINPUT90), .B(KEYINPUT63), .ZN(n368) );
  XOR2_X1 U518 ( .A(n664), .B(KEYINPUT60), .Z(n369) );
  AND2_X1 U519 ( .A1(n532), .A2(G217), .ZN(n370) );
  NAND2_X1 U520 ( .A1(n629), .A2(KEYINPUT30), .ZN(n377) );
  XNOR2_X1 U521 ( .A(n405), .B(n371), .ZN(n710) );
  NAND2_X1 U522 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U523 ( .A1(n430), .A2(n364), .ZN(n382) );
  NAND2_X1 U524 ( .A1(n344), .A2(n383), .ZN(n734) );
  INV_X1 U525 ( .A(n562), .ZN(n385) );
  NAND2_X1 U526 ( .A1(n683), .A2(KEYINPUT40), .ZN(n386) );
  NOR2_X1 U527 ( .A1(n628), .A2(n355), .ZN(n389) );
  INV_X1 U528 ( .A(n580), .ZN(n390) );
  NAND2_X1 U529 ( .A1(n628), .A2(n355), .ZN(n392) );
  NAND2_X1 U530 ( .A1(n580), .A2(n355), .ZN(n393) );
  XNOR2_X1 U531 ( .A(n400), .B(n399), .ZN(G75) );
  NAND2_X1 U532 ( .A1(n401), .A2(n719), .ZN(n400) );
  XNOR2_X1 U533 ( .A(n402), .B(KEYINPUT121), .ZN(n401) );
  NAND2_X1 U534 ( .A1(n427), .A2(n660), .ZN(n402) );
  NAND2_X1 U535 ( .A1(n430), .A2(n365), .ZN(n663) );
  AND2_X1 U536 ( .A1(n430), .A2(n532), .ZN(n403) );
  NAND2_X1 U537 ( .A1(n430), .A2(n370), .ZN(n700) );
  NAND2_X1 U538 ( .A1(n430), .A2(n366), .ZN(n694) );
  NAND2_X1 U539 ( .A1(n430), .A2(n367), .ZN(n697) );
  NAND2_X1 U540 ( .A1(n403), .A2(G478), .ZN(n475) );
  NAND2_X2 U541 ( .A1(n413), .A2(n410), .ZN(n430) );
  XNOR2_X1 U542 ( .A(n428), .B(KEYINPUT2), .ZN(n427) );
  INV_X1 U543 ( .A(n640), .ZN(n609) );
  NAND2_X1 U544 ( .A1(n640), .A2(n346), .ZN(n558) );
  XNOR2_X2 U545 ( .A(n440), .B(n342), .ZN(n640) );
  NAND2_X1 U546 ( .A1(n607), .A2(n406), .ZN(n599) );
  AND2_X1 U547 ( .A1(n407), .A2(n609), .ZN(n406) );
  NAND2_X1 U548 ( .A1(n412), .A2(n409), .ZN(n417) );
  INV_X1 U549 ( .A(n718), .ZN(n409) );
  NAND2_X1 U550 ( .A1(n718), .A2(KEYINPUT2), .ZN(n414) );
  NAND2_X1 U551 ( .A1(n341), .A2(KEYINPUT2), .ZN(n415) );
  NAND2_X1 U552 ( .A1(n417), .A2(n416), .ZN(n428) );
  NOR2_X1 U553 ( .A1(n638), .A2(n418), .ZN(n559) );
  XNOR2_X1 U554 ( .A(n418), .B(KEYINPUT1), .ZN(n637) );
  NOR2_X1 U555 ( .A1(n567), .A2(n418), .ZN(n578) );
  XNOR2_X2 U556 ( .A(n549), .B(G469), .ZN(n418) );
  NAND2_X1 U557 ( .A1(n734), .A2(n735), .ZN(n419) );
  NOR2_X1 U558 ( .A1(n729), .A2(n354), .ZN(n421) );
  XNOR2_X1 U559 ( .A(n429), .B(n347), .ZN(n665) );
  NAND2_X1 U560 ( .A1(n431), .A2(n608), .ZN(n604) );
  XNOR2_X1 U561 ( .A(n612), .B(KEYINPUT106), .ZN(n431) );
  NOR2_X1 U562 ( .A1(n637), .A2(n638), .ZN(n612) );
  INV_X1 U563 ( .A(n606), .ZN(n470) );
  XNOR2_X1 U564 ( .A(n432), .B(n369), .ZN(G60) );
  NAND2_X1 U565 ( .A1(n437), .A2(n380), .ZN(n432) );
  XNOR2_X1 U566 ( .A(n434), .B(n433), .ZN(G51) );
  NAND2_X1 U567 ( .A1(n445), .A2(n380), .ZN(n434) );
  XNOR2_X1 U568 ( .A(n436), .B(n435), .ZN(G54) );
  NAND2_X1 U569 ( .A1(n444), .A2(n380), .ZN(n436) );
  XNOR2_X1 U570 ( .A(n663), .B(n361), .ZN(n437) );
  AND2_X1 U571 ( .A1(n623), .A2(n624), .ZN(n452) );
  XNOR2_X1 U572 ( .A(n573), .B(KEYINPUT36), .ZN(n574) );
  XNOR2_X1 U573 ( .A(n348), .B(n525), .ZN(n526) );
  NAND2_X1 U574 ( .A1(n452), .A2(n350), .ZN(n442) );
  XNOR2_X1 U575 ( .A(n697), .B(n362), .ZN(n444) );
  XNOR2_X1 U576 ( .A(n694), .B(n360), .ZN(n445) );
  NAND2_X1 U577 ( .A1(n522), .A2(G217), .ZN(n508) );
  INV_X1 U578 ( .A(n687), .ZN(n678) );
  NAND2_X1 U579 ( .A1(n576), .A2(n683), .ZN(n450) );
  XNOR2_X1 U580 ( .A(n687), .B(KEYINPUT103), .ZN(n576) );
  XNOR2_X1 U581 ( .A(n519), .B(n511), .ZN(n451) );
  XNOR2_X2 U582 ( .A(n481), .B(G143), .ZN(n512) );
  OR2_X1 U583 ( .A1(n665), .A2(n459), .ZN(n456) );
  NAND2_X1 U584 ( .A1(n665), .A2(n462), .ZN(n458) );
  INV_X1 U585 ( .A(n521), .ZN(n462) );
  XNOR2_X2 U586 ( .A(n469), .B(n359), .ZN(n731) );
  NAND2_X1 U587 ( .A1(n471), .A2(n470), .ZN(n469) );
  XNOR2_X1 U588 ( .A(n605), .B(n472), .ZN(n471) );
  INV_X1 U589 ( .A(KEYINPUT34), .ZN(n472) );
  AND2_X1 U590 ( .A1(n656), .A2(n655), .ZN(n476) );
  XNOR2_X1 U591 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U592 ( .A(n512), .B(n482), .ZN(n483) );
  XNOR2_X1 U593 ( .A(n484), .B(n483), .ZN(n490) );
  XNOR2_X1 U594 ( .A(n526), .B(n527), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n597), .B(KEYINPUT81), .ZN(n598) );
  NOR2_X1 U596 ( .A1(G952), .A2(n719), .ZN(n703) );
  NAND2_X1 U597 ( .A1(G224), .A2(n719), .ZN(n479) );
  XNOR2_X1 U598 ( .A(n520), .B(G125), .ZN(n482) );
  XNOR2_X1 U599 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U600 ( .A(G110), .B(G104), .ZN(n489) );
  XNOR2_X1 U601 ( .A(n490), .B(n710), .ZN(n693) );
  XOR2_X2 U602 ( .A(G902), .B(KEYINPUT15), .Z(n532) );
  XNOR2_X1 U603 ( .A(n491), .B(KEYINPUT79), .ZN(n550) );
  XNOR2_X1 U604 ( .A(KEYINPUT13), .B(G475), .ZN(n505) );
  NAND2_X1 U605 ( .A1(G214), .A2(n515), .ZN(n492) );
  XNOR2_X1 U606 ( .A(n493), .B(n492), .ZN(n497) );
  XNOR2_X1 U607 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U608 ( .A(n497), .B(n496), .Z(n503) );
  XNOR2_X1 U609 ( .A(G125), .B(G140), .ZN(n498) );
  XNOR2_X1 U610 ( .A(n498), .B(KEYINPUT10), .ZN(n529) );
  XNOR2_X1 U611 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U612 ( .A(n529), .B(n501), .ZN(n502) );
  XNOR2_X1 U613 ( .A(n503), .B(n502), .ZN(n662) );
  NOR2_X1 U614 ( .A1(G902), .A2(n662), .ZN(n504) );
  XNOR2_X1 U615 ( .A(n505), .B(n504), .ZN(n582) );
  XNOR2_X1 U616 ( .A(n507), .B(n506), .ZN(n511) );
  XNOR2_X1 U617 ( .A(n509), .B(n508), .ZN(n510) );
  NAND2_X1 U618 ( .A1(n582), .A2(n561), .ZN(n683) );
  XNOR2_X1 U619 ( .A(KEYINPUT75), .B(G472), .ZN(n521) );
  XOR2_X1 U620 ( .A(n513), .B(KEYINPUT99), .Z(n514) );
  NAND2_X1 U621 ( .A1(n515), .A2(G210), .ZN(n516) );
  NAND2_X1 U622 ( .A1(G221), .A2(n522), .ZN(n527) );
  XNOR2_X1 U623 ( .A(G146), .B(G128), .ZN(n524) );
  XNOR2_X1 U624 ( .A(n349), .B(n524), .ZN(n525) );
  XNOR2_X1 U625 ( .A(G137), .B(KEYINPUT72), .ZN(n544) );
  INV_X1 U626 ( .A(n544), .ZN(n528) );
  XOR2_X1 U627 ( .A(n529), .B(n528), .Z(n715) );
  XNOR2_X1 U628 ( .A(n530), .B(n715), .ZN(n701) );
  XNOR2_X1 U629 ( .A(KEYINPUT97), .B(KEYINPUT80), .ZN(n531) );
  NAND2_X1 U630 ( .A1(G234), .A2(n661), .ZN(n533) );
  XNOR2_X1 U631 ( .A(KEYINPUT20), .B(n533), .ZN(n536) );
  NAND2_X1 U632 ( .A1(n536), .A2(G217), .ZN(n534) );
  NAND2_X1 U633 ( .A1(n536), .A2(G221), .ZN(n537) );
  NAND2_X1 U634 ( .A1(G234), .A2(G237), .ZN(n538) );
  XNOR2_X1 U635 ( .A(n538), .B(KEYINPUT14), .ZN(n540) );
  NAND2_X1 U636 ( .A1(n540), .A2(G902), .ZN(n588) );
  NOR2_X1 U637 ( .A1(G900), .A2(n588), .ZN(n539) );
  NAND2_X1 U638 ( .A1(G953), .A2(n539), .ZN(n542) );
  NAND2_X1 U639 ( .A1(n540), .A2(G952), .ZN(n541) );
  XNOR2_X1 U640 ( .A(KEYINPUT93), .B(n541), .ZN(n655) );
  NAND2_X1 U641 ( .A1(n655), .A2(n719), .ZN(n591) );
  NAND2_X1 U642 ( .A1(n542), .A2(n591), .ZN(n557) );
  NAND2_X1 U643 ( .A1(n346), .A2(n557), .ZN(n543) );
  NOR2_X1 U644 ( .A1(n640), .A2(n543), .ZN(n565) );
  NAND2_X1 U645 ( .A1(n719), .A2(G227), .ZN(n545) );
  XOR2_X1 U646 ( .A(n545), .B(n544), .Z(n546) );
  XOR2_X1 U647 ( .A(n546), .B(KEYINPUT95), .Z(n548) );
  NAND2_X1 U648 ( .A1(n550), .A2(G214), .ZN(n551) );
  XOR2_X1 U649 ( .A(KEYINPUT92), .B(n551), .Z(n629) );
  NOR2_X1 U650 ( .A1(n600), .A2(n629), .ZN(n552) );
  NAND2_X1 U651 ( .A1(n572), .A2(n552), .ZN(n553) );
  XNOR2_X1 U652 ( .A(KEYINPUT107), .B(n553), .ZN(n554) );
  XOR2_X1 U653 ( .A(KEYINPUT43), .B(n554), .Z(n555) );
  NAND2_X1 U654 ( .A1(n571), .A2(n555), .ZN(n556) );
  XNOR2_X1 U655 ( .A(n556), .B(KEYINPUT108), .ZN(n727) );
  XNOR2_X1 U656 ( .A(n558), .B(KEYINPUT70), .ZN(n638) );
  XNOR2_X1 U657 ( .A(n559), .B(KEYINPUT98), .ZN(n615) );
  NAND2_X1 U658 ( .A1(n560), .A2(n615), .ZN(n580) );
  XOR2_X1 U659 ( .A(KEYINPUT38), .B(n571), .Z(n628) );
  NOR2_X1 U660 ( .A1(n562), .A2(n576), .ZN(n691) );
  INV_X1 U661 ( .A(KEYINPUT40), .ZN(n563) );
  INV_X1 U662 ( .A(n564), .ZN(n602) );
  NAND2_X1 U663 ( .A1(n602), .A2(n565), .ZN(n566) );
  XNOR2_X1 U664 ( .A(n566), .B(KEYINPUT28), .ZN(n567) );
  XOR2_X1 U665 ( .A(KEYINPUT109), .B(KEYINPUT41), .Z(n569) );
  NOR2_X1 U666 ( .A1(n628), .A2(n629), .ZN(n633) );
  NOR2_X1 U667 ( .A1(n582), .A2(n581), .ZN(n630) );
  NAND2_X1 U668 ( .A1(n633), .A2(n630), .ZN(n568) );
  XNOR2_X1 U669 ( .A(n569), .B(n568), .ZN(n657) );
  NAND2_X1 U670 ( .A1(n578), .A2(n657), .ZN(n570) );
  XNOR2_X1 U671 ( .A(n570), .B(KEYINPUT42), .ZN(n735) );
  XOR2_X1 U672 ( .A(n600), .B(KEYINPUT89), .Z(n596) );
  NAND2_X1 U673 ( .A1(n574), .A2(n596), .ZN(n575) );
  XNOR2_X1 U674 ( .A(n575), .B(KEYINPUT111), .ZN(n729) );
  INV_X1 U675 ( .A(n632), .ZN(n618) );
  INV_X1 U676 ( .A(n594), .ZN(n577) );
  INV_X1 U677 ( .A(n585), .ZN(n579) );
  NAND2_X1 U678 ( .A1(KEYINPUT47), .A2(n579), .ZN(n584) );
  NAND2_X1 U679 ( .A1(n582), .A2(n581), .ZN(n606) );
  NOR2_X1 U680 ( .A1(n571), .A2(n606), .ZN(n583) );
  NAND2_X1 U681 ( .A1(n390), .A2(n583), .ZN(n681) );
  XNOR2_X1 U682 ( .A(KEYINPUT47), .B(KEYINPUT71), .ZN(n586) );
  INV_X1 U683 ( .A(n588), .ZN(n589) );
  NOR2_X1 U684 ( .A1(G898), .A2(n719), .ZN(n712) );
  NAND2_X1 U685 ( .A1(n589), .A2(n712), .ZN(n590) );
  NAND2_X1 U686 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U687 ( .A(KEYINPUT94), .B(n592), .Z(n593) );
  XOR2_X1 U688 ( .A(KEYINPUT66), .B(KEYINPUT32), .Z(n597) );
  NOR2_X1 U689 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U690 ( .A1(n443), .A2(n603), .ZN(n677) );
  NAND2_X1 U691 ( .A1(n733), .A2(n677), .ZN(n626) );
  NAND2_X1 U692 ( .A1(n626), .A2(KEYINPUT44), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n658), .A2(n614), .ZN(n605) );
  NAND2_X1 U694 ( .A1(n731), .A2(KEYINPUT44), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n443), .A2(n607), .ZN(n611) );
  OR2_X1 U696 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U697 ( .A1(n611), .A2(n610), .ZN(n668) );
  AND2_X1 U698 ( .A1(n612), .A2(n646), .ZN(n648) );
  NAND2_X1 U699 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U700 ( .A1(n646), .A2(n616), .ZN(n671) );
  NOR2_X1 U701 ( .A1(n688), .A2(n671), .ZN(n617) );
  NOR2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U703 ( .A1(n668), .A2(n619), .ZN(n620) );
  NAND2_X1 U704 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U705 ( .A(n622), .B(KEYINPUT87), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n636), .A2(n340), .ZN(n652) );
  AND2_X1 U711 ( .A1(n638), .A2(n443), .ZN(n639) );
  XOR2_X1 U712 ( .A(KEYINPUT50), .B(n639), .Z(n644) );
  NOR2_X1 U713 ( .A1(n346), .A2(n640), .ZN(n641) );
  XOR2_X1 U714 ( .A(KEYINPUT49), .B(n641), .Z(n642) );
  XNOR2_X1 U715 ( .A(KEYINPUT119), .B(n642), .ZN(n643) );
  NAND2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U717 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U718 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U719 ( .A(KEYINPUT51), .B(n649), .ZN(n650) );
  NAND2_X1 U720 ( .A1(n650), .A2(n657), .ZN(n651) );
  NAND2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n653), .B(KEYINPUT52), .ZN(n654) );
  XNOR2_X1 U723 ( .A(KEYINPUT120), .B(n654), .ZN(n656) );
  AND2_X1 U724 ( .A1(n340), .A2(n657), .ZN(n659) );
  INV_X1 U725 ( .A(KEYINPUT67), .ZN(n664) );
  XOR2_X1 U726 ( .A(n665), .B(KEYINPUT112), .Z(n667) );
  XOR2_X1 U727 ( .A(KEYINPUT88), .B(KEYINPUT62), .Z(n666) );
  XOR2_X1 U728 ( .A(G101), .B(n668), .Z(G3) );
  XOR2_X1 U729 ( .A(G104), .B(KEYINPUT113), .Z(n670) );
  NAND2_X1 U730 ( .A1(n671), .A2(n441), .ZN(n669) );
  XNOR2_X1 U731 ( .A(n670), .B(n669), .ZN(G6) );
  XNOR2_X1 U732 ( .A(G107), .B(KEYINPUT114), .ZN(n675) );
  XOR2_X1 U733 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n673) );
  NAND2_X1 U734 ( .A1(n671), .A2(n687), .ZN(n672) );
  XNOR2_X1 U735 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U736 ( .A(n675), .B(n674), .ZN(G9) );
  XOR2_X1 U737 ( .A(G110), .B(KEYINPUT115), .Z(n676) );
  XNOR2_X1 U738 ( .A(n677), .B(n676), .ZN(G12) );
  NOR2_X1 U739 ( .A1(n678), .A2(n682), .ZN(n680) );
  XNOR2_X1 U740 ( .A(G128), .B(KEYINPUT29), .ZN(n679) );
  XNOR2_X1 U741 ( .A(n680), .B(n679), .ZN(G30) );
  XNOR2_X1 U742 ( .A(G143), .B(n681), .ZN(G45) );
  NOR2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U744 ( .A(KEYINPUT116), .B(n684), .Z(n685) );
  XNOR2_X1 U745 ( .A(G146), .B(n685), .ZN(G48) );
  NAND2_X1 U746 ( .A1(n441), .A2(n688), .ZN(n686) );
  XNOR2_X1 U747 ( .A(G113), .B(n686), .ZN(G15) );
  XOR2_X1 U748 ( .A(G116), .B(KEYINPUT117), .Z(n690) );
  NAND2_X1 U749 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U750 ( .A(n690), .B(n689), .ZN(G18) );
  XOR2_X1 U751 ( .A(G134), .B(n691), .Z(G36) );
  XOR2_X1 U752 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n692) );
  XOR2_X1 U753 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n695) );
  NOR2_X1 U754 ( .A1(n703), .A2(n699), .ZN(G63) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U756 ( .A1(n703), .A2(n702), .ZN(G66) );
  NAND2_X1 U757 ( .A1(G953), .A2(G224), .ZN(n704) );
  XNOR2_X1 U758 ( .A(KEYINPUT61), .B(n704), .ZN(n705) );
  NAND2_X1 U759 ( .A1(n705), .A2(G898), .ZN(n706) );
  XOR2_X1 U760 ( .A(KEYINPUT124), .B(n706), .Z(n709) );
  NOR2_X1 U761 ( .A1(G953), .A2(n341), .ZN(n708) );
  NOR2_X1 U762 ( .A1(n709), .A2(n708), .ZN(n714) );
  XNOR2_X1 U763 ( .A(G101), .B(n710), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U765 ( .A(n714), .B(n713), .Z(G69) );
  XOR2_X1 U766 ( .A(n715), .B(KEYINPUT125), .Z(n716) );
  XNOR2_X1 U767 ( .A(n717), .B(n716), .ZN(n721) );
  XNOR2_X1 U768 ( .A(n718), .B(n721), .ZN(n720) );
  NAND2_X1 U769 ( .A1(n720), .A2(n719), .ZN(n726) );
  XNOR2_X1 U770 ( .A(G227), .B(n721), .ZN(n722) );
  NAND2_X1 U771 ( .A1(n722), .A2(G900), .ZN(n723) );
  XNOR2_X1 U772 ( .A(KEYINPUT126), .B(n723), .ZN(n724) );
  NAND2_X1 U773 ( .A1(n724), .A2(G953), .ZN(n725) );
  NAND2_X1 U774 ( .A1(n726), .A2(n725), .ZN(G72) );
  XNOR2_X1 U775 ( .A(G140), .B(n727), .ZN(n728) );
  XNOR2_X1 U776 ( .A(n728), .B(KEYINPUT118), .ZN(G42) );
  XNOR2_X1 U777 ( .A(G125), .B(n729), .ZN(n730) );
  XNOR2_X1 U778 ( .A(n730), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U779 ( .A(n731), .B(G122), .Z(G24) );
  XOR2_X1 U780 ( .A(G119), .B(KEYINPUT127), .Z(n732) );
  XNOR2_X1 U781 ( .A(n733), .B(n732), .ZN(G21) );
  XNOR2_X1 U782 ( .A(G131), .B(n734), .ZN(G33) );
  XNOR2_X1 U783 ( .A(G137), .B(n735), .ZN(G39) );
endmodule

