

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586;

  OR2_X1 U321 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U322 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U323 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n428) );
  XNOR2_X1 U324 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n471) );
  XOR2_X1 U325 ( .A(n384), .B(n383), .Z(n550) );
  NOR2_X1 U326 ( .A1(n549), .A2(n548), .ZN(n562) );
  XNOR2_X1 U327 ( .A(n345), .B(n289), .ZN(n346) );
  XOR2_X1 U328 ( .A(n344), .B(n343), .Z(n289) );
  XNOR2_X1 U329 ( .A(n347), .B(n346), .ZN(n407) );
  XOR2_X1 U330 ( .A(G50GAT), .B(n369), .Z(n290) );
  XNOR2_X1 U331 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U332 ( .A(n418), .B(n334), .ZN(n335) );
  INV_X1 U333 ( .A(G176GAT), .ZN(n440) );
  INV_X1 U334 ( .A(KEYINPUT74), .ZN(n389) );
  INV_X1 U335 ( .A(G36GAT), .ZN(n377) );
  XNOR2_X1 U336 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U337 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U338 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U339 ( .A(n392), .B(n391), .ZN(n396) );
  XNOR2_X1 U340 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U341 ( .A(n469), .B(KEYINPUT97), .ZN(n484) );
  NOR2_X1 U342 ( .A1(n498), .A2(n430), .ZN(n568) );
  NOR2_X1 U343 ( .A1(n450), .A2(n534), .ZN(n451) );
  XNOR2_X1 U344 ( .A(n472), .B(n471), .ZN(n519) );
  XNOR2_X1 U345 ( .A(n451), .B(KEYINPUT121), .ZN(n565) );
  XOR2_X1 U346 ( .A(n449), .B(n448), .Z(n534) );
  XNOR2_X1 U347 ( .A(n452), .B(G190GAT), .ZN(n453) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n474) );
  XNOR2_X1 U349 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XNOR2_X1 U350 ( .A(n475), .B(n474), .ZN(G1330GAT) );
  XOR2_X1 U351 ( .A(G204GAT), .B(KEYINPUT22), .Z(n292) );
  XNOR2_X1 U352 ( .A(G218GAT), .B(KEYINPUT90), .ZN(n291) );
  XNOR2_X1 U353 ( .A(n292), .B(n291), .ZN(n308) );
  XOR2_X1 U354 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n294) );
  NAND2_X1 U355 ( .A1(G228GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U356 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U357 ( .A(n295), .B(KEYINPUT23), .Z(n301) );
  XOR2_X1 U358 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n297) );
  XNOR2_X1 U359 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n296) );
  XNOR2_X1 U360 ( .A(n297), .B(n296), .ZN(n315) );
  XOR2_X1 U361 ( .A(G78GAT), .B(G148GAT), .Z(n299) );
  XNOR2_X1 U362 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n298) );
  XNOR2_X1 U363 ( .A(n299), .B(n298), .ZN(n385) );
  XNOR2_X1 U364 ( .A(n315), .B(n385), .ZN(n300) );
  XNOR2_X1 U365 ( .A(n301), .B(n300), .ZN(n304) );
  XOR2_X1 U366 ( .A(G211GAT), .B(KEYINPUT21), .Z(n303) );
  XNOR2_X1 U367 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n302) );
  XNOR2_X1 U368 ( .A(n303), .B(n302), .ZN(n419) );
  XOR2_X1 U369 ( .A(n304), .B(n419), .Z(n306) );
  XOR2_X1 U370 ( .A(G50GAT), .B(G162GAT), .Z(n342) );
  XOR2_X1 U371 ( .A(G22GAT), .B(G155GAT), .Z(n358) );
  XNOR2_X1 U372 ( .A(n342), .B(n358), .ZN(n305) );
  XNOR2_X1 U373 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U374 ( .A(n308), .B(n307), .Z(n464) );
  XOR2_X1 U375 ( .A(G134GAT), .B(KEYINPUT75), .Z(n338) );
  XOR2_X1 U376 ( .A(G85GAT), .B(G162GAT), .Z(n310) );
  XNOR2_X1 U377 ( .A(G29GAT), .B(G148GAT), .ZN(n309) );
  XNOR2_X1 U378 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U379 ( .A(n338), .B(n311), .Z(n313) );
  NAND2_X1 U380 ( .A1(G225GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U381 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U382 ( .A(n314), .B(G57GAT), .Z(n317) );
  XNOR2_X1 U383 ( .A(n315), .B(KEYINPUT92), .ZN(n316) );
  XNOR2_X1 U384 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U385 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n319) );
  XNOR2_X1 U386 ( .A(G1GAT), .B(G155GAT), .ZN(n318) );
  XNOR2_X1 U387 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U388 ( .A(n321), .B(n320), .Z(n330) );
  XNOR2_X1 U389 ( .A(G127GAT), .B(KEYINPUT81), .ZN(n322) );
  XNOR2_X1 U390 ( .A(n322), .B(KEYINPUT0), .ZN(n323) );
  XOR2_X1 U391 ( .A(n323), .B(KEYINPUT80), .Z(n325) );
  XNOR2_X1 U392 ( .A(G113GAT), .B(G120GAT), .ZN(n324) );
  XNOR2_X1 U393 ( .A(n325), .B(n324), .ZN(n445) );
  XOR2_X1 U394 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n327) );
  XNOR2_X1 U395 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n326) );
  XNOR2_X1 U396 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U397 ( .A(n445), .B(n328), .ZN(n329) );
  XOR2_X1 U398 ( .A(n330), .B(n329), .Z(n520) );
  INV_X1 U399 ( .A(n520), .ZN(n498) );
  XOR2_X1 U400 ( .A(G99GAT), .B(G85GAT), .Z(n388) );
  XNOR2_X1 U401 ( .A(G36GAT), .B(G190GAT), .ZN(n331) );
  XNOR2_X1 U402 ( .A(n331), .B(G218GAT), .ZN(n418) );
  NAND2_X1 U403 ( .A1(G232GAT), .A2(G233GAT), .ZN(n333) );
  INV_X1 U404 ( .A(KEYINPUT65), .ZN(n332) );
  XOR2_X1 U405 ( .A(n388), .B(n335), .Z(n340) );
  XOR2_X1 U406 ( .A(G29GAT), .B(G43GAT), .Z(n337) );
  XNOR2_X1 U407 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n336) );
  XNOR2_X1 U408 ( .A(n337), .B(n336), .ZN(n382) );
  XNOR2_X1 U409 ( .A(n382), .B(n338), .ZN(n339) );
  XNOR2_X1 U410 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U411 ( .A(n341), .B(KEYINPUT9), .Z(n347) );
  XNOR2_X1 U412 ( .A(n342), .B(G92GAT), .ZN(n345) );
  XOR2_X1 U413 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n344) );
  XNOR2_X1 U414 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n343) );
  XOR2_X1 U415 ( .A(KEYINPUT36), .B(n407), .Z(n583) );
  XOR2_X1 U416 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n349) );
  XNOR2_X1 U417 ( .A(KEYINPUT77), .B(KEYINPUT15), .ZN(n348) );
  XNOR2_X1 U418 ( .A(n349), .B(n348), .ZN(n366) );
  XOR2_X1 U419 ( .A(KEYINPUT76), .B(KEYINPUT78), .Z(n351) );
  NAND2_X1 U420 ( .A1(G231GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U421 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U422 ( .A(n352), .B(KEYINPUT14), .Z(n357) );
  XNOR2_X1 U423 ( .A(G15GAT), .B(G1GAT), .ZN(n353) );
  XNOR2_X1 U424 ( .A(n353), .B(KEYINPUT69), .ZN(n369) );
  XOR2_X1 U425 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n355) );
  XNOR2_X1 U426 ( .A(G71GAT), .B(G57GAT), .ZN(n354) );
  XNOR2_X1 U427 ( .A(n355), .B(n354), .ZN(n399) );
  XNOR2_X1 U428 ( .A(n369), .B(n399), .ZN(n356) );
  XNOR2_X1 U429 ( .A(n357), .B(n356), .ZN(n362) );
  XOR2_X1 U430 ( .A(G8GAT), .B(G183GAT), .Z(n420) );
  XOR2_X1 U431 ( .A(n420), .B(G211GAT), .Z(n360) );
  XNOR2_X1 U432 ( .A(G78GAT), .B(n358), .ZN(n359) );
  XNOR2_X1 U433 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U434 ( .A(n362), .B(n361), .Z(n364) );
  XNOR2_X1 U435 ( .A(G127GAT), .B(G64GAT), .ZN(n363) );
  XNOR2_X1 U436 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U437 ( .A(n366), .B(n365), .Z(n581) );
  INV_X1 U438 ( .A(n581), .ZN(n559) );
  NAND2_X1 U439 ( .A1(n583), .A2(n559), .ZN(n368) );
  XOR2_X1 U440 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n367) );
  XNOR2_X1 U441 ( .A(n368), .B(n367), .ZN(n403) );
  NAND2_X1 U442 ( .A1(G229GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U443 ( .A(n290), .B(n370), .ZN(n380) );
  XOR2_X1 U444 ( .A(G197GAT), .B(G22GAT), .Z(n372) );
  XNOR2_X1 U445 ( .A(G169GAT), .B(G141GAT), .ZN(n371) );
  XNOR2_X1 U446 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U447 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n374) );
  XNOR2_X1 U448 ( .A(G113GAT), .B(G8GAT), .ZN(n373) );
  XNOR2_X1 U449 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U450 ( .A(n376), .B(n375), .ZN(n378) );
  XOR2_X1 U451 ( .A(n381), .B(KEYINPUT67), .Z(n384) );
  XNOR2_X1 U452 ( .A(n382), .B(KEYINPUT68), .ZN(n383) );
  XOR2_X1 U453 ( .A(n385), .B(KEYINPUT72), .Z(n387) );
  NAND2_X1 U454 ( .A1(G230GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U455 ( .A(n387), .B(n386), .ZN(n392) );
  XNOR2_X1 U456 ( .A(G120GAT), .B(n388), .ZN(n390) );
  XOR2_X1 U457 ( .A(KEYINPUT32), .B(KEYINPUT71), .Z(n394) );
  XNOR2_X1 U458 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U460 ( .A(n396), .B(n395), .Z(n401) );
  XOR2_X1 U461 ( .A(G64GAT), .B(G92GAT), .Z(n398) );
  XNOR2_X1 U462 ( .A(G176GAT), .B(G204GAT), .ZN(n397) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n421) );
  XNOR2_X1 U464 ( .A(n421), .B(n399), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n575) );
  NOR2_X1 U466 ( .A1(n550), .A2(n575), .ZN(n402) );
  AND2_X1 U467 ( .A1(n403), .A2(n402), .ZN(n404) );
  XNOR2_X1 U468 ( .A(n404), .B(KEYINPUT113), .ZN(n413) );
  INV_X1 U469 ( .A(n550), .ZN(n569) );
  XNOR2_X1 U470 ( .A(n575), .B(KEYINPUT41), .ZN(n555) );
  NOR2_X1 U471 ( .A1(n569), .A2(n555), .ZN(n405) );
  XNOR2_X1 U472 ( .A(n405), .B(KEYINPUT46), .ZN(n406) );
  NOR2_X1 U473 ( .A1(n559), .A2(n406), .ZN(n408) );
  INV_X1 U474 ( .A(n407), .ZN(n563) );
  NAND2_X1 U475 ( .A1(n408), .A2(n407), .ZN(n411) );
  XNOR2_X1 U476 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n409), .B(KEYINPUT47), .ZN(n410) );
  XNOR2_X1 U478 ( .A(n411), .B(n410), .ZN(n412) );
  NAND2_X1 U479 ( .A1(n413), .A2(n412), .ZN(n414) );
  XNOR2_X1 U480 ( .A(n414), .B(KEYINPUT48), .ZN(n533) );
  XOR2_X1 U481 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n416) );
  XNOR2_X1 U482 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n415) );
  XNOR2_X1 U483 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U484 ( .A(G169GAT), .B(n417), .Z(n448) );
  INV_X1 U485 ( .A(n448), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n425) );
  XOR2_X1 U487 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U488 ( .A1(G226GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U489 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U491 ( .A(n427), .B(n426), .Z(n501) );
  NAND2_X1 U492 ( .A1(n533), .A2(n501), .ZN(n429) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n430) );
  NAND2_X1 U494 ( .A1(n464), .A2(n568), .ZN(n431) );
  XOR2_X1 U495 ( .A(n431), .B(KEYINPUT55), .Z(n450) );
  XOR2_X1 U496 ( .A(G71GAT), .B(KEYINPUT82), .Z(n433) );
  XNOR2_X1 U497 ( .A(G15GAT), .B(G183GAT), .ZN(n432) );
  XNOR2_X1 U498 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U499 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n435) );
  XNOR2_X1 U500 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n434) );
  XNOR2_X1 U501 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U502 ( .A(n437), .B(n436), .Z(n447) );
  XOR2_X1 U503 ( .A(G190GAT), .B(G99GAT), .Z(n439) );
  XNOR2_X1 U504 ( .A(G43GAT), .B(G134GAT), .ZN(n438) );
  XNOR2_X1 U505 ( .A(n439), .B(n438), .ZN(n443) );
  NAND2_X1 U506 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U507 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U508 ( .A(n447), .B(n446), .ZN(n449) );
  NOR2_X1 U509 ( .A1(n565), .A2(n407), .ZN(n454) );
  XNOR2_X1 U510 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n452) );
  INV_X1 U511 ( .A(n534), .ZN(n492) );
  NAND2_X1 U512 ( .A1(n492), .A2(n501), .ZN(n455) );
  NAND2_X1 U513 ( .A1(n455), .A2(n464), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n456), .B(KEYINPUT25), .ZN(n457) );
  XNOR2_X1 U515 ( .A(n457), .B(KEYINPUT96), .ZN(n461) );
  INV_X1 U516 ( .A(n501), .ZN(n522) );
  XOR2_X1 U517 ( .A(KEYINPUT27), .B(KEYINPUT94), .Z(n458) );
  XOR2_X1 U518 ( .A(n522), .B(n458), .Z(n463) );
  NOR2_X1 U519 ( .A1(n492), .A2(n464), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n459), .B(KEYINPUT26), .ZN(n567) );
  INV_X1 U521 ( .A(n567), .ZN(n549) );
  NOR2_X1 U522 ( .A1(n463), .A2(n549), .ZN(n460) );
  NOR2_X1 U523 ( .A1(n461), .A2(n460), .ZN(n462) );
  NOR2_X1 U524 ( .A1(n498), .A2(n462), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n463), .A2(n520), .ZN(n532) );
  XOR2_X1 U526 ( .A(n464), .B(KEYINPUT28), .Z(n505) );
  INV_X1 U527 ( .A(n505), .ZN(n536) );
  NAND2_X1 U528 ( .A1(n532), .A2(n536), .ZN(n465) );
  NOR2_X1 U529 ( .A1(n492), .A2(n465), .ZN(n466) );
  XOR2_X1 U530 ( .A(KEYINPUT95), .B(n466), .Z(n467) );
  NOR2_X1 U531 ( .A1(n559), .A2(n484), .ZN(n470) );
  NAND2_X1 U532 ( .A1(n583), .A2(n470), .ZN(n472) );
  NOR2_X1 U533 ( .A1(n569), .A2(n575), .ZN(n485) );
  NAND2_X1 U534 ( .A1(n519), .A2(n485), .ZN(n473) );
  XOR2_X1 U535 ( .A(KEYINPUT38), .B(n473), .Z(n504) );
  NAND2_X1 U536 ( .A1(n504), .A2(n492), .ZN(n475) );
  NOR2_X1 U537 ( .A1(n565), .A2(n555), .ZN(n478) );
  XNOR2_X1 U538 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n476), .B(G176GAT), .ZN(n477) );
  XNOR2_X1 U540 ( .A(n478), .B(n477), .ZN(G1349GAT) );
  NOR2_X1 U541 ( .A1(n569), .A2(n565), .ZN(n481) );
  INV_X1 U542 ( .A(G169GAT), .ZN(n479) );
  XNOR2_X1 U543 ( .A(n479), .B(KEYINPUT122), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n481), .B(n480), .ZN(G1348GAT) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n488) );
  NAND2_X1 U546 ( .A1(n559), .A2(n407), .ZN(n482) );
  XNOR2_X1 U547 ( .A(n482), .B(KEYINPUT16), .ZN(n483) );
  NOR2_X1 U548 ( .A1(n484), .A2(n483), .ZN(n509) );
  NAND2_X1 U549 ( .A1(n509), .A2(n485), .ZN(n486) );
  XOR2_X1 U550 ( .A(KEYINPUT98), .B(n486), .Z(n496) );
  NAND2_X1 U551 ( .A1(n498), .A2(n496), .ZN(n487) );
  XNOR2_X1 U552 ( .A(n488), .B(n487), .ZN(G1324GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n490) );
  NAND2_X1 U554 ( .A1(n496), .A2(n501), .ZN(n489) );
  XNOR2_X1 U555 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U556 ( .A(G8GAT), .B(n491), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n494) );
  NAND2_X1 U558 ( .A1(n496), .A2(n492), .ZN(n493) );
  XNOR2_X1 U559 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U560 ( .A(G15GAT), .B(n495), .Z(G1326GAT) );
  NAND2_X1 U561 ( .A1(n496), .A2(n505), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n497), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT39), .Z(n500) );
  NAND2_X1 U564 ( .A1(n498), .A2(n504), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  XOR2_X1 U566 ( .A(G36GAT), .B(KEYINPUT103), .Z(n503) );
  NAND2_X1 U567 ( .A1(n504), .A2(n501), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(G1329GAT) );
  XNOR2_X1 U569 ( .A(G50GAT), .B(KEYINPUT104), .ZN(n507) );
  NAND2_X1 U570 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(G1331GAT) );
  NOR2_X1 U572 ( .A1(n555), .A2(n550), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n508), .B(KEYINPUT106), .ZN(n518) );
  NAND2_X1 U574 ( .A1(n509), .A2(n518), .ZN(n515) );
  NOR2_X1 U575 ( .A1(n520), .A2(n515), .ZN(n511) );
  XNOR2_X1 U576 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U579 ( .A1(n522), .A2(n515), .ZN(n513) );
  XOR2_X1 U580 ( .A(G64GAT), .B(n513), .Z(G1333GAT) );
  NOR2_X1 U581 ( .A1(n534), .A2(n515), .ZN(n514) );
  XOR2_X1 U582 ( .A(G71GAT), .B(n514), .Z(G1334GAT) );
  NOR2_X1 U583 ( .A1(n536), .A2(n515), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n529) );
  NOR2_X1 U587 ( .A1(n520), .A2(n529), .ZN(n521) );
  XOR2_X1 U588 ( .A(G85GAT), .B(n521), .Z(G1336GAT) );
  NOR2_X1 U589 ( .A1(n522), .A2(n529), .ZN(n524) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(KEYINPUT107), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n524), .B(n523), .ZN(G1337GAT) );
  NOR2_X1 U592 ( .A1(n534), .A2(n529), .ZN(n525) );
  XOR2_X1 U593 ( .A(KEYINPUT108), .B(n525), .Z(n526) );
  XNOR2_X1 U594 ( .A(G99GAT), .B(n526), .ZN(G1338GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n528) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U597 ( .A(n528), .B(n527), .ZN(n531) );
  NOR2_X1 U598 ( .A1(n536), .A2(n529), .ZN(n530) );
  XOR2_X1 U599 ( .A(n531), .B(n530), .Z(G1339GAT) );
  NAND2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n548) );
  NOR2_X1 U601 ( .A1(n534), .A2(n548), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n535), .B(KEYINPUT114), .ZN(n537) );
  NAND2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n544) );
  NOR2_X1 U604 ( .A1(n569), .A2(n544), .ZN(n538) );
  XOR2_X1 U605 ( .A(G113GAT), .B(n538), .Z(G1340GAT) );
  NOR2_X1 U606 ( .A1(n555), .A2(n544), .ZN(n540) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NOR2_X1 U609 ( .A1(n581), .A2(n544), .ZN(n542) );
  XNOR2_X1 U610 ( .A(KEYINPUT115), .B(KEYINPUT50), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  NOR2_X1 U613 ( .A1(n407), .A2(n544), .ZN(n546) );
  XNOR2_X1 U614 ( .A(KEYINPUT51), .B(KEYINPUT116), .ZN(n545) );
  XNOR2_X1 U615 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U616 ( .A(G134GAT), .B(n547), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n562), .A2(n550), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n553) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U622 ( .A(KEYINPUT52), .B(n554), .Z(n558) );
  INV_X1 U623 ( .A(n555), .ZN(n556) );
  NAND2_X1 U624 ( .A1(n562), .A2(n556), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  XOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT119), .Z(n561) );
  NAND2_X1 U627 ( .A1(n562), .A2(n559), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U631 ( .A1(n581), .A2(n565), .ZN(n566) );
  XOR2_X1 U632 ( .A(G183GAT), .B(n566), .Z(G1350GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n580) );
  NOR2_X1 U634 ( .A1(n569), .A2(n580), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT124), .B(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  INV_X1 U640 ( .A(n580), .ZN(n584) );
  AND2_X1 U641 ( .A1(n584), .A2(n575), .ZN(n579) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n577) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(G211GAT), .B(n582), .Z(G1354GAT) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(KEYINPUT62), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

