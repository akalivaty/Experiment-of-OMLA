//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n201), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(new_n204), .A2(G50), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT0), .ZN(new_n213));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n210), .ZN(new_n215));
  INV_X1    g0015(.A(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n212), .B1(new_n213), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G116), .ZN(new_n222));
  INV_X1    g0022(.A(G270), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G68), .A2(G238), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n225), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n224), .B(new_n229), .C1(G58), .C2(G232), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n215), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT1), .Z(new_n232));
  AOI211_X1 g0032(.A(new_n220), .B(new_n232), .C1(new_n213), .C2(new_n219), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT2), .ZN(new_n237));
  INV_X1    g0037(.A(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n223), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G97), .B(G107), .Z(new_n244));
  INV_X1    g0044(.A(G87), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  INV_X1    g0048(.A(G50), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n202), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G351));
  OAI21_X1  g0052(.A(G20), .B1(new_n201), .B2(new_n204), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G150), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n253), .B(new_n255), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n209), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n214), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n260), .A2(new_n262), .B1(new_n249), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n261), .A2(new_n209), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n214), .A2(G20), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n265), .B1(new_n249), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT66), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT3), .B(G33), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G223), .A3(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(G222), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G77), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n274), .B(new_n276), .C1(new_n277), .C2(new_n273), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n214), .B1(G41), .B2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n279), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n281), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G226), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n280), .A2(new_n284), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G190), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n269), .A2(new_n270), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(G200), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n272), .A2(new_n291), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(new_n269), .C1(G169), .C2(new_n290), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n273), .A2(G232), .A3(G1698), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT67), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n300), .A2(new_n301), .B1(G33), .B2(G97), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n273), .A2(G226), .A3(new_n275), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n302), .B(new_n303), .C1(new_n301), .C2(new_n300), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n279), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n287), .A2(G238), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n305), .A2(KEYINPUT69), .A3(new_n306), .A4(new_n284), .ZN(new_n307));
  NAND2_X1  g0107(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT13), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n305), .A2(new_n311), .A3(new_n306), .A4(new_n284), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT69), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n283), .B1(new_n304), .B2(new_n279), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n315), .A2(KEYINPUT69), .A3(new_n306), .A4(new_n308), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n310), .A2(new_n314), .A3(G190), .A4(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT70), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n313), .A2(new_n312), .B1(new_n307), .B2(new_n309), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n320), .A2(KEYINPUT70), .A3(G190), .A4(new_n316), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n257), .A2(G77), .B1(new_n254), .B2(G50), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n210), .B2(G68), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(KEYINPUT11), .A3(new_n262), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n203), .B2(new_n268), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n263), .A2(G68), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT12), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT11), .B1(new_n324), .B2(new_n262), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n326), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G200), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n315), .A2(new_n306), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT13), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(new_n333), .B2(new_n312), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n322), .A2(new_n330), .A3(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n310), .A2(new_n314), .A3(G179), .A4(new_n316), .ZN(new_n337));
  NAND2_X1  g0137(.A1(KEYINPUT71), .A2(KEYINPUT14), .ZN(new_n338));
  INV_X1    g0138(.A(new_n312), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n311), .B1(new_n315), .B2(new_n306), .ZN(new_n340));
  OAI211_X1 g0140(.A(G169), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G169), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n333), .B2(new_n312), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT71), .B(KEYINPUT14), .Z(new_n344));
  OAI211_X1 g0144(.A(new_n337), .B(new_n341), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n330), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n259), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(new_n254), .B1(G20), .B2(G77), .ZN(new_n349));
  XOR2_X1   g0149(.A(KEYINPUT15), .B(G87), .Z(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n258), .B2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n262), .B1(new_n277), .B2(new_n264), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n277), .B2(new_n268), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n287), .A2(G244), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G238), .A2(G1698), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n273), .B(new_n356), .C1(new_n235), .C2(G1698), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(new_n279), .C1(G107), .C2(new_n273), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(new_n284), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n354), .B1(G200), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G190), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(new_n359), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n336), .A2(new_n347), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT3), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT72), .B1(new_n364), .B2(G33), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT72), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(new_n256), .A3(KEYINPUT3), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT73), .B1(new_n256), .B2(KEYINPUT3), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(new_n364), .A3(G33), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n238), .A2(G1698), .ZN(new_n373));
  OR2_X1    g0173(.A1(G223), .A2(G1698), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n368), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n256), .B2(new_n245), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n279), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n286), .A2(new_n235), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n284), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G200), .ZN(new_n381));
  XNOR2_X1  g0181(.A(G58), .B(G68), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(G20), .B1(G159), .B2(new_n254), .ZN(new_n383));
  AOI21_X1  g0183(.A(G20), .B1(new_n368), .B2(new_n372), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  OAI21_X1  g0185(.A(G68), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n365), .A2(new_n367), .B1(new_n369), .B2(new_n371), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n387), .A2(KEYINPUT7), .A3(G20), .ZN(new_n388));
  OAI211_X1 g0188(.A(KEYINPUT16), .B(new_n383), .C1(new_n386), .C2(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(KEYINPUT74), .B(KEYINPUT7), .C1(new_n273), .C2(G20), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n364), .A2(G33), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n394));
  OR2_X1    g0194(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n393), .A2(new_n210), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n383), .B1(new_n397), .B2(new_n203), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n389), .A2(new_n400), .A3(new_n262), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n348), .A2(new_n267), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT75), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n264), .A2(new_n262), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n403), .A2(new_n404), .B1(new_n264), .B2(new_n259), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n377), .A2(G190), .A3(new_n284), .A4(new_n379), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n381), .A2(new_n401), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT17), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n401), .A2(new_n405), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n377), .A2(G179), .A3(new_n284), .A4(new_n379), .ZN(new_n410));
  AOI211_X1 g0210(.A(new_n283), .B(new_n378), .C1(new_n376), .C2(new_n279), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n410), .B1(new_n411), .B2(new_n342), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n409), .A2(new_n412), .A3(KEYINPUT18), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n408), .A2(new_n417), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n359), .A2(G179), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n359), .A2(new_n342), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n354), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NOR4_X1   g0222(.A1(new_n299), .A2(new_n363), .A3(new_n418), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT81), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT21), .ZN(new_n425));
  INV_X1    g0225(.A(G45), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(G1), .ZN(new_n427));
  AND2_X1   g0227(.A1(KEYINPUT5), .A2(G41), .ZN(new_n428));
  NOR2_X1   g0228(.A1(KEYINPUT5), .A2(G41), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n430), .A2(new_n282), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n285), .A2(new_n430), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n431), .B1(new_n223), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G264), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(new_n275), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n368), .A2(new_n372), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n393), .A2(G303), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n368), .A2(new_n372), .A3(G257), .A4(new_n275), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT78), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT78), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n387), .A2(new_n441), .A3(G257), .A4(new_n275), .ZN(new_n442));
  AOI211_X1 g0242(.A(KEYINPUT79), .B(new_n438), .C1(new_n440), .C2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT79), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n440), .A2(new_n442), .ZN(new_n445));
  INV_X1    g0245(.A(new_n438), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n433), .B1(new_n448), .B2(new_n279), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n264), .A2(new_n222), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n214), .A2(G33), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n266), .A2(new_n263), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G116), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n222), .A2(G20), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n262), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT80), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G283), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n458), .B(new_n210), .C1(G33), .C2(new_n227), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT20), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n456), .A2(KEYINPUT80), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n462), .B1(new_n262), .B2(new_n455), .ZN(new_n463));
  OAI211_X1 g0263(.A(KEYINPUT20), .B(new_n459), .C1(new_n461), .C2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n450), .B(new_n454), .C1(new_n460), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G169), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n425), .B1(new_n449), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n449), .A2(G179), .A3(new_n466), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n445), .A2(new_n446), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT79), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n445), .A2(new_n444), .A3(new_n446), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n279), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n433), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n467), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT21), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n468), .A2(new_n469), .A3(new_n477), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n473), .A2(G190), .A3(new_n474), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n331), .B1(new_n473), .B2(new_n474), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n479), .A2(new_n480), .A3(new_n466), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n424), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n468), .A2(new_n469), .A3(new_n477), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n485), .A2(new_n481), .A3(KEYINPUT81), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G294), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n387), .B1(G250), .B2(G1698), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n275), .A2(G257), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n279), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n432), .A2(new_n434), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n493), .A2(G179), .A3(new_n431), .A4(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n431), .ZN(new_n497));
  AOI211_X1 g0297(.A(new_n497), .B(new_n494), .C1(new_n492), .C2(new_n279), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n496), .B1(new_n498), .B2(new_n342), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n245), .A2(G20), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n368), .A2(new_n372), .A3(KEYINPUT22), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n391), .A3(new_n392), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT22), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT23), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n210), .B2(G107), .ZN(new_n506));
  INV_X1    g0306(.A(G107), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n507), .A2(KEYINPUT23), .A3(G20), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n503), .A2(new_n504), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n257), .A2(G116), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n502), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT82), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT82), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n502), .A2(new_n509), .A3(new_n513), .A4(new_n510), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT24), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n512), .A2(KEYINPUT24), .A3(new_n514), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n262), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT25), .B1(new_n263), .B2(G107), .ZN(new_n520));
  OR3_X1    g0320(.A1(new_n263), .A2(KEYINPUT25), .A3(G107), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n520), .B(new_n521), .C1(new_n452), .C2(new_n507), .ZN(new_n522));
  XOR2_X1   g0322(.A(new_n522), .B(KEYINPUT83), .Z(new_n523));
  NAND2_X1  g0323(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT84), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT84), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n519), .A2(new_n526), .A3(new_n523), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n500), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n498), .A2(G190), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n493), .A2(new_n431), .A3(new_n495), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G200), .ZN(new_n531));
  AND4_X1   g0331(.A1(new_n523), .A2(new_n529), .A3(new_n519), .A4(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n368), .A2(new_n372), .A3(G244), .A4(new_n275), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n391), .A2(new_n392), .A3(G250), .A4(G1698), .ZN(new_n536));
  AND2_X1   g0336(.A1(KEYINPUT4), .A2(G244), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n391), .A2(new_n392), .A3(new_n537), .A4(new_n275), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n538), .A3(new_n458), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n279), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n285), .A2(new_n430), .A3(G257), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n540), .A2(G190), .A3(new_n431), .A4(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n539), .B1(new_n533), .B2(new_n534), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n431), .B(new_n541), .C1(new_n543), .C2(new_n285), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G200), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n263), .A2(G97), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n507), .A2(KEYINPUT6), .A3(G97), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n244), .B2(KEYINPUT6), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G20), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n254), .A2(G77), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n549), .B(new_n550), .C1(new_n397), .C2(new_n507), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n546), .B1(new_n551), .B2(new_n262), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n453), .A2(G97), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n542), .A2(new_n545), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n551), .A2(new_n262), .ZN(new_n555));
  INV_X1    g0355(.A(new_n546), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(new_n553), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n540), .A2(new_n296), .A3(new_n431), .A4(new_n541), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n544), .A2(new_n342), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT19), .B1(new_n257), .B2(G97), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n245), .A2(KEYINPUT76), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n245), .A2(KEYINPUT76), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n227), .B(new_n507), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n210), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n561), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n368), .A2(new_n372), .A3(new_n210), .A4(G68), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n266), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n452), .A2(new_n351), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n350), .A2(new_n263), .ZN(new_n571));
  OR3_X1    g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n368), .A2(new_n372), .A3(G244), .A4(G1698), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n368), .A2(new_n372), .A3(G238), .A4(new_n275), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n573), .B(new_n574), .C1(new_n256), .C2(new_n222), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n279), .ZN(new_n576));
  INV_X1    g0376(.A(new_n427), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n282), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n285), .A2(G250), .A3(new_n577), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n576), .A2(new_n296), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n580), .ZN(new_n582));
  AOI211_X1 g0382(.A(new_n578), .B(new_n582), .C1(new_n575), .C2(new_n279), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n572), .B(new_n581), .C1(new_n583), .C2(G169), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n576), .A2(G190), .A3(new_n579), .A4(new_n580), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT77), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n452), .B2(new_n245), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n404), .A2(KEYINPUT77), .A3(G87), .A4(new_n451), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n589), .A2(new_n569), .A3(new_n571), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n585), .B(new_n590), .C1(new_n583), .C2(new_n331), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n554), .A2(new_n560), .A3(new_n584), .A4(new_n591), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n528), .A2(new_n532), .A3(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n423), .A2(new_n488), .A3(new_n593), .ZN(G372));
  INV_X1    g0394(.A(new_n298), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT86), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n409), .A2(new_n412), .A3(KEYINPUT18), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT18), .B1(new_n409), .B2(new_n412), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n415), .A2(KEYINPUT86), .A3(new_n416), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n345), .A2(new_n346), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n336), .B2(new_n422), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT17), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n407), .B(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n599), .B(new_n600), .C1(new_n602), .C2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n595), .B1(new_n605), .B2(new_n295), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n524), .A2(new_n499), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n468), .A2(new_n469), .A3(new_n477), .A4(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n532), .A2(new_n592), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT85), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n608), .A2(KEYINPUT85), .A3(new_n609), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT26), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n584), .A2(new_n591), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(new_n560), .ZN(new_n616));
  INV_X1    g0416(.A(new_n560), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(KEYINPUT26), .A3(new_n584), .A4(new_n591), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n612), .A2(new_n584), .A3(new_n613), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n423), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n606), .A2(new_n622), .ZN(G369));
  NOR2_X1   g0423(.A1(new_n216), .A2(G20), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n214), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n625), .A2(KEYINPUT27), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(KEYINPUT27), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(G213), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(G343), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n484), .A2(new_n487), .B1(new_n466), .B2(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n485), .A2(new_n466), .A3(new_n630), .ZN(new_n632));
  OAI21_X1  g0432(.A(G330), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n525), .A2(new_n527), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n499), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n630), .ZN(new_n637));
  INV_X1    g0437(.A(new_n532), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT87), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT87), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n636), .A2(new_n637), .A3(new_n641), .A4(new_n638), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n640), .B(new_n642), .C1(new_n500), .C2(new_n637), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n607), .A2(new_n630), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n640), .A2(new_n642), .ZN(new_n646));
  INV_X1    g0446(.A(new_n630), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n485), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n645), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n644), .A2(new_n650), .ZN(G399));
  NOR2_X1   g0451(.A1(new_n217), .A2(G41), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n208), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n652), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G1), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n564), .A2(G116), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n657), .B(KEYINPUT28), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n621), .A2(new_n647), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(KEYINPUT29), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT88), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n619), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n609), .B1(new_n485), .B2(new_n528), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n618), .A2(new_n661), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n662), .A2(new_n663), .A3(new_n584), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n647), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(KEYINPUT29), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n593), .B(new_n647), .C1(new_n483), .C2(new_n486), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n475), .A2(new_n296), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n498), .A2(new_n541), .A3(new_n540), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n583), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT30), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n498), .A2(new_n583), .A3(G179), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n675), .A2(new_n475), .A3(new_n544), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n670), .A2(KEYINPUT30), .A3(new_n583), .A4(new_n671), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n630), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n669), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n679), .A2(KEYINPUT31), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G330), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n668), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n658), .B1(new_n684), .B2(G1), .ZN(G364));
  AOI21_X1  g0485(.A(new_n655), .B1(G45), .B2(new_n624), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n251), .A2(G45), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n387), .A2(new_n217), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n208), .A2(new_n426), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n218), .A2(G355), .A3(new_n273), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n691), .B(new_n692), .C1(G116), .C2(new_n218), .ZN(new_n693));
  NOR2_X1   g0493(.A1(G13), .A2(G33), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G20), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n209), .B1(G20), .B2(new_n342), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT89), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n687), .B1(new_n693), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n210), .A2(new_n361), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n296), .A2(G200), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT90), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n705), .A2(new_n706), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n210), .A2(G190), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT92), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n713), .A2(G179), .A3(G200), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n711), .A2(G322), .B1(G329), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n361), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G326), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n296), .A2(new_n331), .A3(G190), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G20), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G294), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n716), .A2(G190), .ZN(new_n724));
  XNOR2_X1  g0524(.A(KEYINPUT33), .B(G317), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n331), .A2(G179), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n703), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G303), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n704), .A2(new_n712), .ZN(new_n731));
  INV_X1    g0531(.A(G311), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n393), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n713), .A2(G179), .A3(new_n331), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n733), .B1(new_n734), .B2(G283), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n715), .A2(new_n726), .A3(new_n730), .A4(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n734), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n507), .ZN(new_n738));
  INV_X1    g0538(.A(new_n717), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n721), .A2(new_n227), .B1(new_n739), .B2(new_n249), .ZN(new_n740));
  INV_X1    g0540(.A(new_n724), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n273), .B1(new_n741), .B2(new_n203), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n738), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n710), .A2(new_n202), .B1(new_n277), .B2(new_n731), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT91), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OR3_X1    g0546(.A1(new_n728), .A2(new_n562), .A3(new_n563), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n744), .A2(new_n745), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n743), .A2(new_n746), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n714), .A2(G159), .ZN(new_n750));
  XNOR2_X1  g0550(.A(KEYINPUT93), .B(KEYINPUT32), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n750), .B(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n736), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT94), .Z(new_n754));
  OR2_X1    g0554(.A1(new_n631), .A2(new_n632), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n696), .B(KEYINPUT95), .Z(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n702), .B1(new_n699), .B2(new_n754), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n755), .A2(G330), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n633), .A2(new_n687), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(G396));
  INV_X1    g0561(.A(new_n354), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n362), .B1(new_n762), .B2(new_n647), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n421), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n421), .A2(new_n630), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n659), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n767), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n621), .A2(new_n647), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  OR3_X1    g0571(.A1(new_n771), .A2(new_n682), .A3(KEYINPUT99), .ZN(new_n772));
  OAI21_X1  g0572(.A(KEYINPUT99), .B1(new_n771), .B2(new_n682), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n771), .A2(new_n682), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n772), .A2(new_n687), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n734), .A2(G68), .ZN(new_n776));
  INV_X1    g0576(.A(new_n387), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(G58), .B2(new_n720), .ZN(new_n778));
  INV_X1    g0578(.A(new_n714), .ZN(new_n779));
  INV_X1    g0579(.A(G132), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n776), .B(new_n778), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G50), .B2(new_n729), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT98), .Z(new_n783));
  AOI22_X1  g0583(.A1(G137), .A2(new_n717), .B1(new_n724), .B2(G150), .ZN(new_n784));
  INV_X1    g0584(.A(G159), .ZN(new_n785));
  INV_X1    g0585(.A(G143), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n784), .B1(new_n785), .B2(new_n731), .C1(new_n710), .C2(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT34), .Z(new_n788));
  NOR2_X1   g0588(.A1(new_n737), .A2(new_n245), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n711), .A2(G294), .B1(G311), .B2(new_n714), .ZN(new_n790));
  INV_X1    g0590(.A(new_n731), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n791), .A2(G116), .B1(G283), .B2(new_n724), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT97), .ZN(new_n793));
  INV_X1    g0593(.A(G303), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n393), .B1(new_n739), .B2(new_n794), .C1(new_n721), .C2(new_n227), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(G107), .B2(new_n729), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n790), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n783), .A2(new_n788), .B1(new_n789), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n698), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n698), .A2(new_n694), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n686), .B1(G77), .B2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT96), .Z(new_n803));
  OAI211_X1 g0603(.A(new_n799), .B(new_n803), .C1(new_n769), .C2(new_n695), .ZN(new_n804));
  AND3_X1   g0604(.A1(new_n775), .A2(KEYINPUT100), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(KEYINPUT100), .B1(new_n775), .B2(new_n804), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G384));
  OAI21_X1  g0608(.A(new_n423), .B1(new_n660), .B2(new_n667), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n606), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT106), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT102), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n613), .A2(new_n584), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n619), .B1(new_n610), .B2(new_n611), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n630), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n765), .B1(new_n815), .B2(new_n769), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n330), .A2(new_n647), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n346), .B(new_n334), .C1(new_n319), .C2(new_n321), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(new_n601), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n336), .B(new_n347), .C1(new_n330), .C2(new_n647), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n812), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT103), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n383), .B1(new_n386), .B2(new_n388), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n399), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n825), .A2(new_n262), .A3(new_n389), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n405), .ZN(new_n827));
  INV_X1    g0627(.A(new_n628), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n412), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n829), .A2(KEYINPUT37), .A3(new_n407), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n827), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n408), .B2(new_n417), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(new_n833), .B2(new_n828), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n409), .A2(new_n828), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n413), .A2(new_n835), .A3(new_n407), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT37), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT38), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n597), .A2(new_n598), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n828), .B(new_n827), .C1(new_n604), .C2(new_n840), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n841), .A2(KEYINPUT38), .A3(new_n838), .A4(new_n830), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n823), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n841), .A2(new_n838), .A3(new_n830), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT38), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(KEYINPUT103), .A3(new_n842), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n770), .A2(new_n766), .ZN(new_n851));
  INV_X1    g0651(.A(new_n821), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(KEYINPUT102), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n822), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n828), .B1(new_n599), .B2(new_n600), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT39), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n847), .B2(new_n842), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n628), .B1(new_n401), .B2(new_n405), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT104), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n836), .B(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n408), .A2(new_n599), .A3(new_n600), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n862), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n842), .B(new_n856), .C1(new_n864), .C2(KEYINPUT38), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n858), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n347), .A2(new_n630), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n855), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n854), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n811), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n767), .B1(new_n819), .B2(new_n820), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n680), .A2(new_n873), .A3(new_n681), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n872), .B1(new_n849), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n680), .A2(new_n681), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n864), .A2(KEYINPUT38), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n877), .B1(new_n878), .B2(new_n842), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n876), .A2(new_n873), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n876), .A2(new_n423), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n881), .B(new_n882), .Z(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(G330), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n870), .B(new_n884), .Z(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n214), .B2(new_n624), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n222), .B1(new_n548), .B2(KEYINPUT35), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n887), .B(new_n211), .C1(KEYINPUT35), .C2(new_n548), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT36), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n208), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT101), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n201), .B2(new_n203), .ZN(new_n892));
  INV_X1    g0692(.A(new_n201), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(KEYINPUT101), .A3(G68), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n890), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(G1), .A3(new_n216), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n886), .A2(new_n889), .A3(new_n896), .ZN(G367));
  INV_X1    g0697(.A(KEYINPUT45), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n646), .A2(new_n649), .ZN(new_n899));
  INV_X1    g0699(.A(new_n645), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n617), .A2(new_n630), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n557), .A2(new_n630), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n554), .A2(new_n560), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n898), .B1(new_n901), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n650), .A2(KEYINPUT45), .A3(new_n905), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n901), .A2(KEYINPUT44), .A3(new_n906), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT44), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n650), .B2(new_n905), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n644), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n644), .A3(new_n913), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n899), .B1(new_n643), .B2(new_n649), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(new_n633), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n919), .A2(new_n683), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n684), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n652), .B(KEYINPUT41), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT108), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n214), .B1(new_n624), .B2(G45), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT108), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n922), .A2(new_n927), .A3(new_n923), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  OR3_X1    g0729(.A1(new_n899), .A2(KEYINPUT42), .A3(new_n904), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n560), .B1(new_n636), .B2(new_n904), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n647), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT42), .B1(new_n899), .B2(new_n904), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n584), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n590), .A2(new_n647), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n615), .B2(new_n936), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT43), .Z(new_n939));
  NAND2_X1  g0739(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT107), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n934), .A2(KEYINPUT43), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n644), .A2(new_n906), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n929), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n729), .A2(G116), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT46), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n720), .A2(G107), .B1(new_n724), .B2(G294), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n948), .A2(new_n777), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n737), .A2(new_n227), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(G283), .ZN(new_n953));
  INV_X1    g0753(.A(G317), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n952), .B1(new_n953), .B2(new_n731), .C1(new_n954), .C2(new_n779), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n710), .A2(new_n794), .B1(new_n732), .B2(new_n739), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n956), .A2(KEYINPUT110), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(KEYINPUT110), .ZN(new_n958));
  OR4_X1    g0758(.A1(new_n950), .A2(new_n955), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n893), .A2(new_n731), .ZN(new_n960));
  INV_X1    g0760(.A(G137), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n779), .A2(new_n961), .B1(new_n202), .B2(new_n728), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT111), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n711), .A2(G150), .B1(G77), .B2(new_n734), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n273), .B1(new_n741), .B2(new_n785), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n721), .A2(new_n203), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(G143), .C2(new_n717), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n964), .A2(new_n965), .A3(new_n966), .A4(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n959), .B1(new_n960), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n687), .B1(new_n973), .B2(new_n698), .ZN(new_n974));
  INV_X1    g0774(.A(new_n689), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n701), .B1(new_n218), .B2(new_n351), .C1(new_n242), .C2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT109), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n974), .B(new_n977), .C1(new_n757), .C2(new_n938), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT113), .Z(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n946), .A2(new_n980), .ZN(G387));
  INV_X1    g0781(.A(new_n920), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n654), .B1(new_n919), .B2(new_n683), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n714), .A2(G326), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G311), .A2(new_n724), .B1(new_n717), .B2(G322), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n794), .B2(new_n731), .C1(new_n710), .C2(new_n954), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT48), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n953), .B2(new_n721), .C1(new_n722), .C2(new_n728), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT49), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n387), .B(new_n985), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n990), .B2(new_n989), .C1(new_n222), .C2(new_n737), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n729), .A2(G77), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n952), .B(new_n993), .C1(new_n203), .C2(new_n731), .ZN(new_n994));
  INV_X1    g0794(.A(G150), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n779), .A2(new_n995), .B1(new_n249), .B2(new_n710), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n994), .A2(new_n777), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n350), .A2(new_n720), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n348), .A2(new_n724), .B1(G159), .B2(new_n717), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT114), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n992), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n687), .B1(new_n1002), .B2(new_n698), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n348), .A2(new_n249), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT50), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n203), .A2(new_n277), .ZN(new_n1006));
  NOR4_X1   g0806(.A1(new_n1005), .A2(G45), .A3(new_n1006), .A4(new_n656), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n689), .B1(new_n239), .B2(new_n426), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n656), .A2(new_n218), .A3(new_n273), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n218), .A2(G107), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n701), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1003), .B(new_n1012), .C1(new_n643), .C2(new_n757), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n984), .B(new_n1013), .C1(new_n926), .C2(new_n919), .ZN(G393));
  NAND2_X1  g0814(.A1(new_n916), .A2(new_n917), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n654), .B1(new_n1015), .B2(new_n982), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1016), .A2(new_n921), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n701), .B1(new_n227), .B2(new_n218), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n247), .B2(new_n689), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n777), .B1(G68), .B2(new_n729), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n720), .A2(G77), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(new_n893), .C2(new_n741), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n245), .A2(new_n737), .B1(new_n779), .B2(new_n786), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT51), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n710), .A2(new_n785), .B1(new_n995), .B2(new_n739), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1022), .B(new_n1023), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n1024), .B2(new_n1025), .C1(new_n259), .C2(new_n731), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n720), .A2(G116), .B1(new_n724), .B2(G303), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1028), .B(new_n393), .C1(new_n722), .C2(new_n731), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1029), .B(new_n738), .C1(G322), .C2(new_n714), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n710), .A2(new_n732), .B1(new_n954), .B2(new_n739), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT52), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1030), .B(new_n1032), .C1(new_n953), .C2(new_n728), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1027), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1019), .B1(new_n1034), .B2(new_n698), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n686), .C1(new_n697), .C2(new_n905), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n1015), .B2(new_n926), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1017), .A2(new_n1037), .ZN(G390));
  INV_X1    g0838(.A(new_n865), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1039), .A2(new_n857), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n821), .B1(new_n770), .B2(new_n766), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1040), .B1(new_n1041), .B2(new_n867), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n764), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n766), .B1(new_n666), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n852), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n867), .B1(new_n878), .B2(new_n842), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n680), .A2(new_n873), .A3(new_n681), .A4(G330), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1042), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n423), .A2(new_n680), .A3(G330), .A4(new_n681), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n809), .A2(new_n606), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n680), .A2(new_n681), .A3(G330), .A4(new_n769), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n821), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1044), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(new_n1059), .A3(new_n1049), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n816), .B1(new_n1058), .B2(new_n1049), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1056), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1053), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n682), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1065), .A2(new_n873), .B1(new_n1057), .B2(new_n821), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1060), .B1(new_n1066), .B2(new_n816), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1067), .A2(new_n1051), .A3(new_n1052), .A4(new_n1056), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1064), .A2(new_n652), .A3(new_n1068), .ZN(new_n1069));
  AND3_X1   g0869(.A1(new_n1042), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1049), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n926), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n686), .B1(new_n348), .B2(new_n801), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT115), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n717), .A2(G128), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n741), .B2(new_n961), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n273), .B1(new_n721), .B2(new_n785), .ZN(new_n1079));
  XOR2_X1   g0879(.A(KEYINPUT54), .B(G143), .Z(new_n1080));
  AOI211_X1 g0880(.A(new_n1078), .B(new_n1079), .C1(new_n791), .C2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n714), .A2(G125), .B1(new_n734), .B2(new_n201), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n711), .A2(G132), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n728), .A2(new_n995), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT53), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n714), .A2(G294), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n273), .B1(new_n729), .B2(G87), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n776), .B(new_n1088), .C1(new_n227), .C2(new_n731), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1021), .B1(new_n739), .B2(new_n953), .C1(new_n507), .C2(new_n741), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n710), .A2(new_n222), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1084), .A2(new_n1086), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT116), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1076), .B1(new_n699), .B2(new_n1094), .C1(new_n866), .C2(new_n695), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1069), .A2(new_n1074), .A3(new_n1095), .ZN(G378));
  AND3_X1   g0896(.A1(new_n875), .A2(G330), .A3(new_n880), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n869), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n269), .A2(new_n828), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n299), .B(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT55), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT56), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT56), .B1(new_n1107), .B2(new_n1102), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n875), .A2(new_n880), .A3(G330), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1110), .A2(new_n868), .A3(new_n854), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1098), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1109), .B1(new_n1098), .B2(new_n1111), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1073), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n351), .A2(new_n731), .B1(new_n721), .B2(new_n203), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n779), .A2(new_n953), .B1(new_n507), .B2(new_n710), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1115), .B(new_n1116), .C1(G116), .C2(new_n717), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n734), .A2(G58), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT117), .Z(new_n1119));
  INV_X1    g0919(.A(G41), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n777), .A2(new_n993), .A3(new_n1120), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT118), .Z(new_n1122));
  NAND3_X1  g0922(.A1(new_n1117), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(G97), .B2(new_n724), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1124), .B(KEYINPUT58), .Z(new_n1125));
  NAND2_X1  g0925(.A1(new_n711), .A2(G128), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n791), .A2(G137), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n720), .A2(G150), .B1(new_n724), .B2(G132), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n729), .A2(new_n1080), .B1(G125), .B2(new_n717), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT59), .Z(new_n1131));
  AOI21_X1  g0931(.A(G41), .B1(new_n714), .B2(G124), .ZN(new_n1132));
  AOI21_X1  g0932(.A(G33), .B1(new_n734), .B2(G159), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(G41), .B1(new_n387), .B2(G33), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1125), .B(new_n1134), .C1(G50), .C2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n687), .B1(new_n1136), .B2(new_n698), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1109), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1137), .B1(new_n201), .B2(new_n801), .C1(new_n1138), .C2(new_n695), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1114), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1055), .B1(new_n1072), .B2(new_n1067), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1098), .A2(new_n1111), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1138), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1098), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1142), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n652), .B1(new_n1146), .B2(KEYINPUT57), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1068), .A2(new_n1056), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1148), .B(KEYINPUT57), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1141), .B1(new_n1147), .B2(new_n1150), .ZN(G375));
  OAI211_X1 g0951(.A(new_n1055), .B(new_n1060), .C1(new_n1066), .C2(new_n816), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT119), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1062), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1155), .A2(KEYINPUT119), .A3(new_n1055), .A4(new_n1060), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1157), .A2(new_n923), .A3(new_n1063), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n387), .B1(new_n785), .B2(new_n728), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n710), .A2(new_n961), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(G128), .C2(new_n714), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n791), .A2(G150), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1080), .A2(new_n724), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n721), .B2(new_n249), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G132), .B2(new_n717), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1119), .A2(new_n1161), .A3(new_n1162), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n273), .B1(new_n717), .B2(G294), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1167), .B1(new_n222), .B2(new_n741), .C1(new_n737), .C2(new_n277), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT121), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n998), .B1(new_n710), .B2(new_n953), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n714), .A2(G303), .B1(G97), .B2(new_n729), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT120), .Z(new_n1173));
  OAI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n731), .A2(new_n507), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1166), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1176), .A2(new_n698), .B1(new_n203), .B2(new_n800), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n686), .B(new_n1177), .C1(new_n852), .C2(new_n695), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1158), .A2(new_n1180), .ZN(G381));
  NOR3_X1   g0981(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT122), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1183), .A2(G381), .A3(G387), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1148), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT57), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1187), .A2(new_n652), .A3(new_n1149), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1140), .A2(G378), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(G390), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1184), .A2(new_n1192), .ZN(G407));
  NAND2_X1  g0993(.A1(new_n1190), .A2(new_n629), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(G407), .A2(G213), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT123), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(G407), .A2(KEYINPUT123), .A3(G213), .A4(new_n1194), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(G409));
  INV_X1    g0999(.A(KEYINPUT60), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1152), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1063), .A2(KEYINPUT60), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n654), .B(new_n1201), .C1(new_n1157), .C2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1180), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n807), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1201), .B1(new_n1157), .B2(new_n1202), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n652), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1207), .A2(G384), .A3(new_n1180), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n629), .A2(G213), .A3(G2897), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1205), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n629), .A2(G213), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1069), .A2(new_n1074), .A3(new_n1095), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1148), .B(new_n923), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1214), .A2(new_n1114), .A3(new_n1139), .A4(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n654), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1140), .B1(new_n1217), .B2(new_n1149), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1213), .B(new_n1216), .C1(new_n1218), .C2(new_n1214), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT61), .B1(new_n1212), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT126), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT62), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1221), .B(new_n1222), .C1(new_n1219), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(G375), .A2(G378), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1189), .A2(new_n1215), .B1(G213), .B2(new_n629), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1225), .A2(KEYINPUT62), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT126), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1214), .B1(new_n1188), .B2(new_n1141), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1216), .A2(new_n1213), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT62), .B1(new_n1232), .B2(new_n1227), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1220), .B(new_n1224), .C1(new_n1229), .C2(new_n1233), .ZN(new_n1234));
  XOR2_X1   g1034(.A(G393), .B(G396), .Z(new_n1235));
  NAND2_X1  g1035(.A1(G387), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1235), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n979), .B1(new_n929), .B2(new_n945), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT124), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1237), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1236), .A2(new_n1240), .A3(G390), .ZN(new_n1241));
  AOI21_X1  g1041(.A(G390), .B1(new_n1236), .B2(new_n1240), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1234), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1209), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1223), .A2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1205), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT63), .B1(new_n1248), .B2(new_n1232), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1232), .A2(new_n1227), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1236), .A2(new_n1240), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1191), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1236), .A2(new_n1240), .A3(G390), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1225), .A2(KEYINPUT63), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT61), .B1(new_n1256), .B2(KEYINPUT125), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1256), .A2(KEYINPUT125), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1251), .A2(new_n1255), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1244), .A2(new_n1259), .ZN(G405));
  INV_X1    g1060(.A(KEYINPUT127), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1253), .A2(KEYINPUT127), .A3(new_n1254), .ZN(new_n1263));
  OR3_X1    g1063(.A1(new_n1190), .A2(new_n1230), .A3(new_n1227), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1227), .B1(new_n1190), .B2(new_n1230), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1262), .A2(new_n1263), .A3(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1243), .A2(KEYINPUT127), .A3(new_n1265), .A4(new_n1264), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(G402));
endmodule


