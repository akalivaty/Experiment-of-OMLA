

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U322 ( .A(n410), .B(n409), .ZN(n417) );
  XNOR2_X1 U323 ( .A(n506), .B(KEYINPUT48), .ZN(n507) );
  XNOR2_X1 U324 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U325 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U326 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n342) );
  XNOR2_X1 U327 ( .A(n343), .B(n342), .ZN(n345) );
  XNOR2_X1 U328 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U329 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n547) );
  XNOR2_X1 U330 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U331 ( .A(n508), .B(n507), .ZN(n541) );
  XNOR2_X1 U332 ( .A(G127GAT), .B(KEYINPUT83), .ZN(n290) );
  XNOR2_X1 U333 ( .A(n290), .B(KEYINPUT82), .ZN(n291) );
  XOR2_X1 U334 ( .A(n291), .B(KEYINPUT0), .Z(n293) );
  XNOR2_X1 U335 ( .A(G113GAT), .B(G134GAT), .ZN(n292) );
  XOR2_X1 U336 ( .A(n293), .B(n292), .Z(n363) );
  INV_X1 U337 ( .A(n363), .ZN(n313) );
  XOR2_X1 U338 ( .A(KEYINPUT5), .B(G57GAT), .Z(n295) );
  XNOR2_X1 U339 ( .A(G1GAT), .B(G148GAT), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U341 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n297) );
  XNOR2_X1 U342 ( .A(KEYINPUT1), .B(KEYINPUT90), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U344 ( .A(n299), .B(n298), .Z(n311) );
  XNOR2_X1 U345 ( .A(KEYINPUT2), .B(KEYINPUT87), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n300), .B(KEYINPUT88), .ZN(n301) );
  XOR2_X1 U347 ( .A(n301), .B(KEYINPUT3), .Z(n303) );
  XNOR2_X1 U348 ( .A(G155GAT), .B(G162GAT), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n385) );
  XOR2_X1 U350 ( .A(G85GAT), .B(G120GAT), .Z(n305) );
  XNOR2_X1 U351 ( .A(G29GAT), .B(G141GAT), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U353 ( .A(KEYINPUT91), .B(n306), .Z(n308) );
  NAND2_X1 U354 ( .A1(G225GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n385), .B(n309), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U358 ( .A(n313), .B(n312), .Z(n543) );
  INV_X1 U359 ( .A(n543), .ZN(n481) );
  XOR2_X1 U360 ( .A(G57GAT), .B(KEYINPUT13), .Z(n427) );
  XOR2_X1 U361 ( .A(G71GAT), .B(G183GAT), .Z(n315) );
  XNOR2_X1 U362 ( .A(G22GAT), .B(G127GAT), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U364 ( .A(n427), .B(n316), .Z(n318) );
  NAND2_X1 U365 ( .A1(G231GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U367 ( .A(n319), .B(KEYINPUT80), .Z(n322) );
  XNOR2_X1 U368 ( .A(G15GAT), .B(G1GAT), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n320), .B(KEYINPUT71), .ZN(n422) );
  XNOR2_X1 U370 ( .A(n422), .B(KEYINPUT79), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n330) );
  XOR2_X1 U372 ( .A(G78GAT), .B(G211GAT), .Z(n324) );
  XNOR2_X1 U373 ( .A(G8GAT), .B(G155GAT), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U375 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n326) );
  XNOR2_X1 U376 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U378 ( .A(n328), .B(n327), .Z(n329) );
  XOR2_X1 U379 ( .A(n330), .B(n329), .Z(n575) );
  INV_X1 U380 ( .A(n575), .ZN(n559) );
  XOR2_X1 U381 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n332) );
  XNOR2_X1 U382 ( .A(G134GAT), .B(G162GAT), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n349) );
  XOR2_X1 U384 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n334) );
  XNOR2_X1 U385 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U387 ( .A(G99GAT), .B(G85GAT), .Z(n434) );
  XOR2_X1 U388 ( .A(n335), .B(n434), .Z(n337) );
  XNOR2_X1 U389 ( .A(G36GAT), .B(G106GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U391 ( .A(G190GAT), .B(KEYINPUT78), .Z(n375) );
  XOR2_X1 U392 ( .A(n375), .B(G92GAT), .Z(n339) );
  NAND2_X1 U393 ( .A1(G232GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U395 ( .A(n341), .B(n340), .Z(n347) );
  XNOR2_X1 U396 ( .A(G43GAT), .B(KEYINPUT70), .ZN(n343) );
  XOR2_X1 U397 ( .A(KEYINPUT7), .B(KEYINPUT69), .Z(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n410) );
  XNOR2_X1 U399 ( .A(n410), .B(G50GAT), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n349), .B(n348), .ZN(n561) );
  INV_X1 U402 ( .A(n561), .ZN(n537) );
  NAND2_X1 U403 ( .A1(n559), .A2(n537), .ZN(n350) );
  XNOR2_X1 U404 ( .A(n350), .B(KEYINPUT16), .ZN(n351) );
  XNOR2_X1 U405 ( .A(KEYINPUT81), .B(n351), .ZN(n405) );
  XOR2_X1 U406 ( .A(G183GAT), .B(KEYINPUT17), .Z(n353) );
  XNOR2_X1 U407 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n371) );
  XOR2_X1 U409 ( .A(G120GAT), .B(G71GAT), .Z(n428) );
  XOR2_X1 U410 ( .A(n371), .B(n428), .Z(n355) );
  NAND2_X1 U411 ( .A1(G227GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U413 ( .A(G176GAT), .B(KEYINPUT20), .Z(n357) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(KEYINPUT84), .ZN(n356) );
  XNOR2_X1 U415 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U416 ( .A(n359), .B(n358), .Z(n365) );
  XOR2_X1 U417 ( .A(G99GAT), .B(G190GAT), .Z(n361) );
  XNOR2_X1 U418 ( .A(G43GAT), .B(G15GAT), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U420 ( .A(n363), .B(n362), .Z(n364) );
  XOR2_X1 U421 ( .A(n365), .B(n364), .Z(n509) );
  INV_X1 U422 ( .A(n509), .ZN(n550) );
  XOR2_X1 U423 ( .A(G64GAT), .B(G92GAT), .Z(n367) );
  XNOR2_X1 U424 ( .A(G176GAT), .B(G204GAT), .ZN(n366) );
  XNOR2_X1 U425 ( .A(n367), .B(n366), .ZN(n429) );
  XOR2_X1 U426 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n373) );
  XOR2_X1 U427 ( .A(KEYINPUT86), .B(G218GAT), .Z(n369) );
  XNOR2_X1 U428 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U430 ( .A(G197GAT), .B(n370), .Z(n383) );
  XNOR2_X1 U431 ( .A(n371), .B(n383), .ZN(n372) );
  XNOR2_X1 U432 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U433 ( .A(n375), .B(n374), .Z(n377) );
  NAND2_X1 U434 ( .A1(G226GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n429), .B(n378), .ZN(n380) );
  XOR2_X1 U437 ( .A(G169GAT), .B(G36GAT), .Z(n379) );
  XNOR2_X1 U438 ( .A(G8GAT), .B(n379), .ZN(n425) );
  XOR2_X1 U439 ( .A(n380), .B(n425), .Z(n484) );
  XNOR2_X1 U440 ( .A(KEYINPUT27), .B(n484), .ZN(n397) );
  NAND2_X1 U441 ( .A1(n481), .A2(n397), .ZN(n523) );
  XOR2_X1 U442 ( .A(G78GAT), .B(G148GAT), .Z(n382) );
  XNOR2_X1 U443 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n382), .B(n381), .ZN(n430) );
  XOR2_X1 U445 ( .A(n430), .B(n383), .Z(n387) );
  XNOR2_X1 U446 ( .A(G50GAT), .B(G22GAT), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n384), .B(G141GAT), .ZN(n408) );
  XNOR2_X1 U448 ( .A(n408), .B(n385), .ZN(n386) );
  XNOR2_X1 U449 ( .A(n387), .B(n386), .ZN(n395) );
  NAND2_X1 U450 ( .A1(G228GAT), .A2(G233GAT), .ZN(n393) );
  XOR2_X1 U451 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n389) );
  XNOR2_X1 U452 ( .A(KEYINPUT85), .B(KEYINPUT23), .ZN(n388) );
  XNOR2_X1 U453 ( .A(n389), .B(n388), .ZN(n391) );
  XOR2_X1 U454 ( .A(KEYINPUT24), .B(G204GAT), .Z(n390) );
  XNOR2_X1 U455 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U457 ( .A(n395), .B(n394), .Z(n546) );
  XNOR2_X1 U458 ( .A(KEYINPUT28), .B(n546), .ZN(n463) );
  INV_X1 U459 ( .A(n463), .ZN(n489) );
  NOR2_X1 U460 ( .A1(n523), .A2(n489), .ZN(n510) );
  NAND2_X1 U461 ( .A1(n550), .A2(n510), .ZN(n404) );
  NOR2_X1 U462 ( .A1(n546), .A2(n509), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n396), .B(KEYINPUT26), .ZN(n567) );
  NAND2_X1 U464 ( .A1(n397), .A2(n567), .ZN(n401) );
  NAND2_X1 U465 ( .A1(n484), .A2(n509), .ZN(n398) );
  NAND2_X1 U466 ( .A1(n546), .A2(n398), .ZN(n399) );
  XOR2_X1 U467 ( .A(KEYINPUT25), .B(n399), .Z(n400) );
  NAND2_X1 U468 ( .A1(n401), .A2(n400), .ZN(n402) );
  NAND2_X1 U469 ( .A1(n402), .A2(n543), .ZN(n403) );
  NAND2_X1 U470 ( .A1(n404), .A2(n403), .ZN(n449) );
  NAND2_X1 U471 ( .A1(n405), .A2(n449), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n406), .B(KEYINPUT94), .ZN(n467) );
  XOR2_X1 U473 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n407) );
  INV_X1 U474 ( .A(n417), .ZN(n416) );
  XOR2_X1 U475 ( .A(KEYINPUT66), .B(KEYINPUT72), .Z(n412) );
  XNOR2_X1 U476 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n414) );
  XOR2_X1 U478 ( .A(G113GAT), .B(G197GAT), .Z(n413) );
  XNOR2_X1 U479 ( .A(n414), .B(n413), .ZN(n418) );
  INV_X1 U480 ( .A(n418), .ZN(n415) );
  NAND2_X1 U481 ( .A1(n416), .A2(n415), .ZN(n420) );
  NAND2_X1 U482 ( .A1(n418), .A2(n417), .ZN(n419) );
  NAND2_X1 U483 ( .A1(n420), .A2(n419), .ZN(n424) );
  NAND2_X1 U484 ( .A1(G229GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n426), .B(n425), .ZN(n492) );
  XNOR2_X1 U486 ( .A(KEYINPUT73), .B(n492), .ZN(n551) );
  XNOR2_X1 U487 ( .A(n428), .B(n427), .ZN(n440) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n438) );
  XOR2_X1 U489 ( .A(KEYINPUT31), .B(KEYINPUT75), .Z(n432) );
  XNOR2_X1 U490 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U492 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U493 ( .A1(G230GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U496 ( .A(n440), .B(n439), .Z(n571) );
  NAND2_X1 U497 ( .A1(n551), .A2(n571), .ZN(n453) );
  NOR2_X1 U498 ( .A1(n467), .A2(n453), .ZN(n447) );
  NAND2_X1 U499 ( .A1(n481), .A2(n447), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n441), .B(KEYINPUT34), .ZN(n442) );
  XNOR2_X1 U501 ( .A(G1GAT), .B(n442), .ZN(G1324GAT) );
  NAND2_X1 U502 ( .A1(n447), .A2(n484), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n443), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U504 ( .A(KEYINPUT95), .B(KEYINPUT35), .Z(n445) );
  NAND2_X1 U505 ( .A1(n447), .A2(n509), .ZN(n444) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U507 ( .A(G15GAT), .B(n446), .Z(G1326GAT) );
  NAND2_X1 U508 ( .A1(n489), .A2(n447), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n448), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U510 ( .A(KEYINPUT36), .B(n561), .Z(n580) );
  NAND2_X1 U511 ( .A1(n575), .A2(n449), .ZN(n450) );
  NOR2_X1 U512 ( .A1(n580), .A2(n450), .ZN(n452) );
  XNOR2_X1 U513 ( .A(KEYINPUT37), .B(KEYINPUT96), .ZN(n451) );
  XNOR2_X1 U514 ( .A(n452), .B(n451), .ZN(n480) );
  NOR2_X1 U515 ( .A1(n480), .A2(n453), .ZN(n454) );
  XOR2_X1 U516 ( .A(KEYINPUT38), .B(n454), .Z(n462) );
  NOR2_X1 U517 ( .A1(n462), .A2(n543), .ZN(n455) );
  XNOR2_X1 U518 ( .A(n455), .B(KEYINPUT39), .ZN(n456) );
  XNOR2_X1 U519 ( .A(G29GAT), .B(n456), .ZN(G1328GAT) );
  INV_X1 U520 ( .A(n484), .ZN(n540) );
  NOR2_X1 U521 ( .A1(n462), .A2(n540), .ZN(n458) );
  XNOR2_X1 U522 ( .A(G36GAT), .B(KEYINPUT97), .ZN(n457) );
  XNOR2_X1 U523 ( .A(n458), .B(n457), .ZN(G1329GAT) );
  XNOR2_X1 U524 ( .A(KEYINPUT40), .B(KEYINPUT98), .ZN(n460) );
  NOR2_X1 U525 ( .A1(n550), .A2(n462), .ZN(n459) );
  XNOR2_X1 U526 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U527 ( .A(G43GAT), .B(n461), .Z(G1330GAT) );
  XNOR2_X1 U528 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n465) );
  NOR2_X1 U529 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U530 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U531 ( .A(G50GAT), .B(n466), .ZN(G1331GAT) );
  XNOR2_X1 U532 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n469) );
  XOR2_X1 U533 ( .A(n571), .B(KEYINPUT41), .Z(n529) );
  XNOR2_X1 U534 ( .A(KEYINPUT101), .B(n529), .ZN(n553) );
  NAND2_X1 U535 ( .A1(n553), .A2(n492), .ZN(n479) );
  NOR2_X1 U536 ( .A1(n467), .A2(n479), .ZN(n474) );
  NAND2_X1 U537 ( .A1(n474), .A2(n481), .ZN(n468) );
  XNOR2_X1 U538 ( .A(n469), .B(n468), .ZN(G1332GAT) );
  NAND2_X1 U539 ( .A1(n474), .A2(n484), .ZN(n470) );
  XNOR2_X1 U540 ( .A(n470), .B(KEYINPUT102), .ZN(n471) );
  XNOR2_X1 U541 ( .A(G64GAT), .B(n471), .ZN(G1333GAT) );
  XOR2_X1 U542 ( .A(G71GAT), .B(KEYINPUT103), .Z(n473) );
  NAND2_X1 U543 ( .A1(n474), .A2(n509), .ZN(n472) );
  XNOR2_X1 U544 ( .A(n473), .B(n472), .ZN(G1334GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n476) );
  NAND2_X1 U546 ( .A1(n474), .A2(n489), .ZN(n475) );
  XNOR2_X1 U547 ( .A(n476), .B(n475), .ZN(n478) );
  XOR2_X1 U548 ( .A(G78GAT), .B(KEYINPUT104), .Z(n477) );
  XNOR2_X1 U549 ( .A(n478), .B(n477), .ZN(G1335GAT) );
  XNOR2_X1 U550 ( .A(G85GAT), .B(KEYINPUT106), .ZN(n483) );
  NOR2_X1 U551 ( .A1(n480), .A2(n479), .ZN(n488) );
  NAND2_X1 U552 ( .A1(n488), .A2(n481), .ZN(n482) );
  XNOR2_X1 U553 ( .A(n483), .B(n482), .ZN(G1336GAT) );
  XOR2_X1 U554 ( .A(G92GAT), .B(KEYINPUT107), .Z(n486) );
  NAND2_X1 U555 ( .A1(n488), .A2(n484), .ZN(n485) );
  XNOR2_X1 U556 ( .A(n486), .B(n485), .ZN(G1337GAT) );
  NAND2_X1 U557 ( .A1(n509), .A2(n488), .ZN(n487) );
  XNOR2_X1 U558 ( .A(n487), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U559 ( .A1(n489), .A2(n488), .ZN(n490) );
  XNOR2_X1 U560 ( .A(n490), .B(KEYINPUT44), .ZN(n491) );
  XNOR2_X1 U561 ( .A(G106GAT), .B(n491), .ZN(G1339GAT) );
  NOR2_X1 U562 ( .A1(n492), .A2(n529), .ZN(n494) );
  XNOR2_X1 U563 ( .A(KEYINPUT46), .B(KEYINPUT109), .ZN(n493) );
  XNOR2_X1 U564 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U565 ( .A(KEYINPUT108), .B(n495), .ZN(n497) );
  AND2_X1 U566 ( .A1(n575), .A2(n537), .ZN(n496) );
  NAND2_X1 U567 ( .A1(n497), .A2(n496), .ZN(n499) );
  XOR2_X1 U568 ( .A(KEYINPUT47), .B(KEYINPUT110), .Z(n498) );
  XNOR2_X1 U569 ( .A(n499), .B(n498), .ZN(n505) );
  NOR2_X1 U570 ( .A1(n575), .A2(n580), .ZN(n501) );
  XNOR2_X1 U571 ( .A(KEYINPUT45), .B(KEYINPUT111), .ZN(n500) );
  XNOR2_X1 U572 ( .A(n501), .B(n500), .ZN(n502) );
  NOR2_X1 U573 ( .A1(n502), .A2(n551), .ZN(n503) );
  NAND2_X1 U574 ( .A1(n571), .A2(n503), .ZN(n504) );
  NAND2_X1 U575 ( .A1(n505), .A2(n504), .ZN(n508) );
  INV_X1 U576 ( .A(KEYINPUT64), .ZN(n506) );
  NAND2_X1 U577 ( .A1(n510), .A2(n509), .ZN(n511) );
  NOR2_X1 U578 ( .A1(n541), .A2(n511), .ZN(n519) );
  NAND2_X1 U579 ( .A1(n519), .A2(n551), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n512), .B(KEYINPUT112), .ZN(n513) );
  XNOR2_X1 U581 ( .A(G113GAT), .B(n513), .ZN(G1340GAT) );
  XOR2_X1 U582 ( .A(G120GAT), .B(KEYINPUT49), .Z(n515) );
  NAND2_X1 U583 ( .A1(n519), .A2(n553), .ZN(n514) );
  XNOR2_X1 U584 ( .A(n515), .B(n514), .ZN(G1341GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n517) );
  NAND2_X1 U586 ( .A1(n519), .A2(n559), .ZN(n516) );
  XNOR2_X1 U587 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U588 ( .A(G127GAT), .B(n518), .ZN(G1342GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n521) );
  NAND2_X1 U590 ( .A1(n519), .A2(n561), .ZN(n520) );
  XNOR2_X1 U591 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U592 ( .A(G134GAT), .B(n522), .ZN(G1343GAT) );
  NOR2_X1 U593 ( .A1(n541), .A2(n523), .ZN(n524) );
  NAND2_X1 U594 ( .A1(n524), .A2(n567), .ZN(n536) );
  NOR2_X1 U595 ( .A1(n492), .A2(n536), .ZN(n526) );
  XNOR2_X1 U596 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n525) );
  XNOR2_X1 U597 ( .A(n526), .B(n525), .ZN(G1344GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n528) );
  XNOR2_X1 U599 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n527) );
  XNOR2_X1 U600 ( .A(n528), .B(n527), .ZN(n533) );
  NOR2_X1 U601 ( .A1(n529), .A2(n536), .ZN(n531) );
  XNOR2_X1 U602 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n530) );
  XNOR2_X1 U603 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U604 ( .A(n533), .B(n532), .ZN(G1345GAT) );
  NOR2_X1 U605 ( .A1(n575), .A2(n536), .ZN(n535) );
  XNOR2_X1 U606 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n534) );
  XNOR2_X1 U607 ( .A(n535), .B(n534), .ZN(G1346GAT) );
  NOR2_X1 U608 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U609 ( .A(KEYINPUT120), .B(n538), .Z(n539) );
  XNOR2_X1 U610 ( .A(G162GAT), .B(n539), .ZN(G1347GAT) );
  NOR2_X1 U611 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U612 ( .A(n542), .B(KEYINPUT54), .ZN(n544) );
  NAND2_X1 U613 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n545), .B(KEYINPUT65), .ZN(n568) );
  NAND2_X1 U615 ( .A1(n546), .A2(n568), .ZN(n548) );
  NOR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n562), .A2(n551), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U619 ( .A1(n553), .A2(n562), .ZN(n558) );
  XOR2_X1 U620 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n555) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U623 ( .A(KEYINPUT122), .B(n556), .Z(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1349GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n562), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1351GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n566) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n579) );
  NOR2_X1 U634 ( .A1(n492), .A2(n579), .ZN(n569) );
  XOR2_X1 U635 ( .A(n570), .B(n569), .Z(G1352GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n579), .ZN(n573) );
  XNOR2_X1 U637 ( .A(KEYINPUT61), .B(KEYINPUT125), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(G204GAT), .B(n574), .Z(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n579), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(n581), .Z(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

