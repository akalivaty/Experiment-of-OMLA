//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n791, new_n792, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896;
  XNOR2_X1  g000(.A(G155gat), .B(G162gat), .ZN(new_n202));
  XOR2_X1   g001(.A(G141gat), .B(G148gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G141gat), .B(G148gat), .ZN(new_n206));
  OR2_X1    g005(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT77), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT77), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G162gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n207), .A2(new_n209), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n206), .B1(new_n213), .B2(KEYINPUT2), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n208), .A2(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G162gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT75), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n218), .B1(new_n215), .B2(new_n217), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n205), .B1(new_n214), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n224));
  OAI21_X1  g023(.A(G113gat), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G113gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G120gat), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT1), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G127gat), .B(G134gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(G127gat), .A2(G134gat), .ZN(new_n230));
  INV_X1    g029(.A(G120gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G113gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n230), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(G134gat), .A3(new_n237), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n228), .A2(new_n229), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n222), .A2(new_n239), .A3(KEYINPUT79), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT79), .B1(new_n222), .B2(new_n239), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT4), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n213), .A2(KEYINPUT2), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n202), .A2(new_n218), .ZN(new_n244));
  INV_X1    g043(.A(new_n220), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n243), .A2(new_n203), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n205), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n229), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n235), .A2(new_n238), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n246), .A2(new_n247), .A3(new_n248), .A4(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n242), .B1(KEYINPUT4), .B2(new_n250), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n251), .A2(KEYINPUT84), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT5), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n254));
  OR3_X1    g053(.A1(new_n222), .A2(KEYINPUT78), .A3(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT78), .B1(new_n222), .B2(new_n254), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n222), .A2(new_n254), .ZN(new_n257));
  INV_X1    g056(.A(new_n239), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n255), .A2(new_n256), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G225gat), .A2(G233gat), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n251), .A2(KEYINPUT84), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n252), .A2(new_n253), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT79), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n250), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n222), .A2(new_n239), .A3(KEYINPUT79), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT80), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n250), .A2(KEYINPUT4), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT80), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n265), .A2(new_n271), .A3(new_n266), .A4(new_n267), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n261), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n222), .A2(new_n239), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n275), .B1(new_n265), .B2(new_n267), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT81), .B1(new_n276), .B2(new_n260), .ZN(new_n277));
  OAI22_X1  g076(.A1(new_n240), .A2(new_n241), .B1(new_n222), .B2(new_n239), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT81), .ZN(new_n279));
  INV_X1    g078(.A(new_n260), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n253), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n274), .A2(new_n282), .A3(KEYINPUT82), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT82), .B1(new_n274), .B2(new_n282), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n263), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G57gat), .B(G85gat), .Z(new_n286));
  XNOR2_X1  g085(.A(G1gat), .B(G29gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n285), .A2(KEYINPUT6), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT85), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n285), .A2(new_n291), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n263), .B(new_n290), .C1(new_n283), .C2(new_n284), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n285), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n291), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n294), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G197gat), .B(G204gat), .Z(new_n301));
  AOI21_X1  g100(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT72), .ZN(new_n304));
  XOR2_X1   g103(.A(G211gat), .B(G218gat), .Z(new_n305));
  OR2_X1    g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT25), .ZN(new_n310));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT24), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G183gat), .ZN(new_n314));
  INV_X1    g113(.A(G190gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT65), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT65), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(G183gat), .B2(G190gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n313), .A2(new_n316), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT23), .ZN(new_n323));
  AND4_X1   g122(.A1(new_n310), .A2(new_n320), .A3(new_n321), .A4(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n322), .A2(KEYINPUT23), .ZN(new_n325));
  INV_X1    g124(.A(G169gat), .ZN(new_n326));
  INV_X1    g125(.A(G176gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT67), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT67), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n329), .B1(G169gat), .B2(G176gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT23), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n313), .B(new_n319), .C1(G183gat), .C2(G190gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT66), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n321), .B(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n332), .A2(new_n325), .A3(new_n333), .A4(new_n335), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n324), .A2(new_n325), .B1(new_n336), .B2(KEYINPUT25), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT27), .B(G183gat), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(new_n315), .ZN(new_n340));
  AND2_X1   g139(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n338), .B(new_n315), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT26), .B1(new_n328), .B2(new_n330), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n321), .B(new_n346), .C1(new_n347), .C2(KEYINPUT68), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n347), .A2(KEYINPUT68), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n311), .B(new_n345), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT29), .B1(new_n337), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G226gat), .A2(G233gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n309), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n352), .B1(new_n337), .B2(new_n350), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n337), .A2(new_n350), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n355), .B1(new_n358), .B2(new_n352), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n308), .B(new_n354), .C1(new_n359), .C2(new_n309), .ZN(new_n360));
  INV_X1    g159(.A(new_n355), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n361), .B1(new_n351), .B2(new_n353), .ZN(new_n362));
  INV_X1    g161(.A(new_n308), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G8gat), .B(G36gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(G64gat), .B(G92gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n365), .A2(new_n369), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT30), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n368), .B1(new_n360), .B2(new_n364), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(KEYINPUT74), .A3(KEYINPUT30), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n370), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n372), .A2(new_n373), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n300), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT31), .B(G22gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(G228gat), .A2(G233gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT3), .B1(new_n363), .B2(new_n357), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(new_n222), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n363), .B1(new_n357), .B2(new_n257), .ZN(new_n388));
  OAI21_X1  g187(.A(G50gat), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n388), .ZN(new_n390));
  INV_X1    g189(.A(G50gat), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n390), .B(new_n391), .C1(new_n222), .C2(new_n386), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n385), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G78gat), .B(G106gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n389), .A2(new_n392), .A3(new_n385), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n395), .ZN(new_n398));
  INV_X1    g197(.A(new_n396), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n398), .B1(new_n399), .B2(new_n393), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n381), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT37), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n365), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n359), .A2(new_n308), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT73), .B1(new_n358), .B2(new_n352), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n406), .B1(new_n362), .B2(KEYINPUT73), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n405), .B(KEYINPUT37), .C1(new_n407), .C2(new_n308), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(new_n368), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT38), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n360), .A2(KEYINPUT37), .A3(new_n364), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n404), .A2(KEYINPUT38), .A3(new_n368), .A4(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n375), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n294), .A2(new_n414), .A3(new_n298), .A4(new_n299), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n252), .A2(new_n259), .A3(new_n262), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n280), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n276), .A2(new_n260), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(KEYINPUT39), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT39), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n416), .A2(new_n420), .A3(new_n280), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n290), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT40), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n419), .A2(KEYINPUT40), .A3(new_n290), .A4(new_n421), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n379), .A2(new_n424), .A3(new_n295), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n397), .A2(new_n400), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n415), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G227gat), .A2(G233gat), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n429), .B(KEYINPUT64), .Z(new_n430));
  NAND2_X1  g229(.A1(new_n356), .A2(new_n258), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n337), .A2(new_n239), .A3(new_n350), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT32), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(G15gat), .B(G43gat), .Z(new_n436));
  XNOR2_X1  g235(.A(G71gat), .B(G99gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n438), .A2(KEYINPUT33), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n438), .B1(new_n433), .B2(KEYINPUT33), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n435), .B(new_n439), .C1(new_n440), .C2(KEYINPUT71), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT71), .ZN(new_n442));
  OAI22_X1  g241(.A1(new_n440), .A2(new_n442), .B1(new_n434), .B2(new_n433), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n431), .A2(new_n430), .A3(new_n432), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n445), .B(KEYINPUT34), .Z(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n444), .A2(new_n447), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n451), .B(KEYINPUT36), .Z(new_n452));
  NAND3_X1  g251(.A1(new_n402), .A2(new_n428), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT35), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT86), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n455), .B1(new_n300), .B2(new_n380), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n451), .A2(KEYINPUT87), .ZN(new_n457));
  INV_X1    g256(.A(new_n450), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n458), .A2(KEYINPUT87), .A3(new_n448), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n427), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n454), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT35), .B1(new_n401), .B2(new_n451), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n454), .A2(KEYINPUT86), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n462), .A2(new_n300), .A3(new_n380), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n453), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G29gat), .A2(G36gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT88), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT15), .ZN(new_n468));
  XOR2_X1   g267(.A(G43gat), .B(G50gat), .Z(new_n469));
  AOI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n468), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NOR3_X1   g271(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n473), .A2(KEYINPUT89), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(KEYINPUT89), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n470), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n476), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(new_n473), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n471), .B1(new_n480), .B2(new_n467), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(KEYINPUT90), .B2(KEYINPUT17), .ZN(new_n483));
  NAND2_X1  g282(.A1(KEYINPUT90), .A2(KEYINPUT17), .ZN(new_n484));
  XOR2_X1   g283(.A(new_n483), .B(new_n484), .Z(new_n485));
  XNOR2_X1  g284(.A(G99gat), .B(G106gat), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT100), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G99gat), .A2(G106gat), .ZN(new_n489));
  INV_X1    g288(.A(G85gat), .ZN(new_n490));
  INV_X1    g289(.A(G92gat), .ZN(new_n491));
  AOI22_X1  g290(.A1(KEYINPUT8), .A2(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT7), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(new_n490), .B2(new_n491), .ZN(new_n494));
  NAND3_X1  g293(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n488), .B(new_n496), .Z(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n485), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT101), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n482), .ZN(new_n502));
  AND2_X1   g301(.A1(G232gat), .A2(G233gat), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n502), .A2(new_n497), .B1(KEYINPUT41), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n485), .A2(KEYINPUT101), .A3(new_n498), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n501), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G190gat), .B(G218gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n506), .A2(new_n507), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n503), .A2(KEYINPUT41), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT99), .ZN(new_n512));
  XOR2_X1   g311(.A(G134gat), .B(G162gat), .Z(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n509), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n506), .A2(new_n507), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n514), .B1(new_n517), .B2(new_n508), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  OR2_X1    g320(.A1(G71gat), .A2(G78gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(G71gat), .A2(G78gat), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n523), .B(KEYINPUT93), .Z(new_n524));
  XNOR2_X1  g323(.A(G57gat), .B(G64gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT94), .ZN(new_n526));
  NOR2_X1   g325(.A1(KEYINPUT93), .A2(KEYINPUT9), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n522), .B(new_n524), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT9), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n523), .B1(new_n522), .B2(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(G57gat), .B(G64gat), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT95), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT21), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT98), .ZN(new_n536));
  INV_X1    g335(.A(G211gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(G127gat), .B(G155gat), .Z(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n536), .B(G211gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n539), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n521), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n541), .A3(new_n521), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n534), .A2(KEYINPUT21), .ZN(new_n547));
  XNOR2_X1  g346(.A(G15gat), .B(G22gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT16), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(G1gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(G1gat), .B2(new_n548), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n551), .B(G8gat), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(G183gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT96), .B(KEYINPUT20), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n559), .B1(new_n557), .B2(new_n556), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n546), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n546), .ZN(new_n564));
  OAI22_X1  g363(.A1(new_n564), .A2(new_n544), .B1(new_n560), .B2(new_n561), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n519), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n465), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n552), .A2(new_n482), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n568), .B1(new_n485), .B2(new_n552), .ZN(new_n569));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT18), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n502), .B(new_n552), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(new_n570), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n571), .A2(new_n572), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT91), .B1(new_n571), .B2(new_n572), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT91), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n569), .A2(new_n580), .A3(KEYINPUT18), .A4(new_n570), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G113gat), .B(G141gat), .ZN(new_n583));
  INV_X1    g382(.A(G197gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT11), .B(G169gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(KEYINPUT12), .Z(new_n588));
  NAND2_X1  g387(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n578), .A2(new_n579), .A3(new_n581), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n534), .A2(new_n497), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n496), .A2(KEYINPUT102), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n496), .A2(KEYINPUT102), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n488), .A3(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n597), .B(KEYINPUT103), .C1(new_n488), .C2(new_n496), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(KEYINPUT103), .B2(new_n597), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n594), .B1(new_n599), .B2(new_n534), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n534), .A2(new_n497), .A3(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G230gat), .A2(G233gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n600), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(G176gat), .B(G204gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT104), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n611), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n593), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n567), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n300), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n379), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT16), .B(G8gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n623), .B(KEYINPUT42), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(G8gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(G1325gat));
  NOR2_X1   g425(.A1(new_n457), .A2(new_n459), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(G15gat), .B1(new_n617), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n452), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n617), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n629), .B1(G15gat), .B2(new_n631), .ZN(G1326gat));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n401), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT43), .B(G22gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(G1327gat));
  INV_X1    g434(.A(new_n519), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n465), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n565), .A2(new_n563), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n616), .A3(new_n639), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n640), .A2(G29gat), .A3(new_n300), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT45), .Z(new_n642));
  XOR2_X1   g441(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n465), .A2(new_n636), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n646), .B1(new_n465), .B2(new_n636), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n639), .A2(new_n616), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(G29gat), .B1(new_n651), .B2(new_n300), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n642), .A2(new_n652), .ZN(G1328gat));
  NOR3_X1   g452(.A1(new_n640), .A2(G36gat), .A3(new_n380), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT46), .ZN(new_n655));
  OAI21_X1  g454(.A(G36gat), .B1(new_n651), .B2(new_n380), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(G1329gat));
  OAI21_X1  g456(.A(G43gat), .B1(new_n651), .B2(new_n452), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT106), .ZN(new_n659));
  AOI21_X1  g458(.A(KEYINPUT47), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n640), .A2(G43gat), .A3(new_n627), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n658), .B(new_n661), .C1(new_n659), .C2(KEYINPUT47), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(G1330gat));
  AOI21_X1  g464(.A(new_n391), .B1(new_n650), .B2(new_n401), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n640), .A2(G50gat), .A3(new_n427), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT107), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g468(.A1(new_n567), .A2(new_n593), .A3(new_n615), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT108), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n300), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g475(.A1(new_n674), .A2(new_n380), .ZN(new_n677));
  NOR2_X1   g476(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n678));
  AND2_X1   g477(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n677), .B2(new_n678), .ZN(G1333gat));
  OAI21_X1  g480(.A(G71gat), .B1(new_n674), .B2(new_n452), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT50), .ZN(new_n683));
  INV_X1    g482(.A(G71gat), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n672), .A2(new_n684), .A3(new_n628), .A4(new_n673), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n683), .B1(new_n682), .B2(new_n685), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(G1334gat));
  NOR2_X1   g487(.A1(new_n674), .A2(new_n427), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT109), .B(G78gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1335gat));
  NAND3_X1  g490(.A1(new_n465), .A2(new_n636), .A3(new_n644), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n637), .B2(new_n646), .ZN(new_n693));
  INV_X1    g492(.A(new_n615), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n638), .A2(new_n694), .A3(new_n592), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n696), .A2(new_n490), .A3(new_n300), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n638), .A2(new_n592), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n465), .A2(new_n636), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT51), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT110), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n465), .A2(KEYINPUT51), .A3(new_n636), .A4(new_n698), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n703), .A2(new_n702), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n704), .A2(new_n705), .A3(new_n618), .A4(new_n615), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n697), .B1(new_n490), .B2(new_n706), .ZN(G1336gat));
  NAND3_X1  g506(.A1(new_n693), .A2(new_n379), .A3(new_n695), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G92gat), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT52), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n380), .A2(G92gat), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n704), .A2(new_n705), .A3(new_n615), .A4(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT112), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n694), .B1(new_n701), .B2(new_n703), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n708), .A2(G92gat), .B1(new_n711), .B2(new_n715), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n716), .A2(KEYINPUT111), .A3(new_n710), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT111), .B1(new_n716), .B2(new_n710), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n714), .A2(new_n719), .ZN(G1337gat));
  OAI21_X1  g519(.A(G99gat), .B1(new_n696), .B2(new_n452), .ZN(new_n721));
  INV_X1    g520(.A(G99gat), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n704), .A2(new_n705), .A3(new_n722), .A4(new_n615), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n627), .B2(new_n723), .ZN(G1338gat));
  OAI211_X1 g523(.A(new_n401), .B(new_n695), .C1(new_n645), .C2(new_n647), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(G106gat), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n427), .A2(G106gat), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n715), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT53), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n729), .A2(new_n615), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n704), .A2(new_n705), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT113), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n704), .A2(new_n705), .A3(new_n735), .A4(new_n732), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n727), .B1(new_n726), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n725), .A2(KEYINPUT114), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT53), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT115), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n693), .A2(new_n738), .A3(new_n401), .A4(new_n695), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n740), .A2(new_n743), .A3(G106gat), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT53), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n744), .A2(new_n734), .A3(new_n745), .A4(new_n736), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n731), .B1(new_n742), .B2(new_n748), .ZN(G1339gat));
  NOR2_X1   g548(.A1(new_n569), .A2(new_n570), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n574), .A2(new_n577), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n587), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n591), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n611), .ZN(new_n754));
  INV_X1    g553(.A(new_n606), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT54), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n604), .A2(new_n605), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(KEYINPUT54), .A3(new_n606), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(KEYINPUT55), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n759), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n753), .A2(new_n760), .A3(new_n613), .A4(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n638), .B1(new_n636), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n592), .A2(new_n613), .A3(new_n763), .A4(new_n760), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n615), .A2(new_n753), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(new_n767), .A3(new_n519), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT116), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n566), .A2(new_n770), .A3(new_n593), .A4(new_n694), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n593), .A2(new_n519), .A3(new_n563), .A4(new_n565), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT116), .B1(new_n772), .B2(new_n615), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n769), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n300), .A2(new_n379), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n460), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n778), .A2(new_n226), .A3(new_n593), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n401), .A2(new_n300), .A3(new_n451), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n774), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n774), .B2(new_n781), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n782), .A2(new_n783), .A3(new_n379), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT118), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n592), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n779), .B1(new_n786), .B2(new_n226), .ZN(G1340gat));
  OAI21_X1  g586(.A(G120gat), .B1(new_n778), .B2(new_n694), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n785), .B1(new_n224), .B2(new_n223), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(new_n694), .ZN(G1341gat));
  NAND2_X1  g589(.A1(new_n236), .A2(new_n237), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n778), .A2(new_n791), .A3(new_n639), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n784), .A2(new_n638), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n793), .B2(new_n791), .ZN(G1342gat));
  INV_X1    g593(.A(G134gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n784), .A2(new_n795), .A3(new_n636), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT119), .B1(new_n796), .B2(KEYINPUT56), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n776), .A2(new_n777), .A3(new_n636), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(G134gat), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n799), .B2(KEYINPUT56), .ZN(new_n800));
  NOR4_X1   g599(.A1(new_n782), .A2(new_n783), .A3(G134gat), .A4(new_n379), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n801), .A2(new_n802), .A3(new_n803), .A4(new_n636), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n797), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n797), .A2(new_n800), .A3(KEYINPUT120), .A4(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1343gat));
  NAND2_X1  g608(.A1(new_n452), .A2(new_n401), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT123), .Z(new_n811));
  AND2_X1   g610(.A1(new_n776), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(G141gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n592), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n774), .A2(new_n401), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n774), .A2(KEYINPUT57), .A3(new_n401), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n452), .A2(new_n775), .ZN(new_n820));
  XOR2_X1   g619(.A(new_n820), .B(KEYINPUT121), .Z(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n592), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G141gat), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n814), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT122), .B1(new_n822), .B2(G141gat), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT58), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT58), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n814), .B2(KEYINPUT124), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT124), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n823), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n827), .B1(new_n829), .B2(new_n831), .ZN(G1344gat));
  INV_X1    g631(.A(G148gat), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n812), .A2(new_n833), .A3(new_n615), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT59), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT125), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n566), .A2(new_n593), .A3(new_n694), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n769), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n769), .B2(new_n837), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n838), .A2(new_n839), .A3(new_n427), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n818), .B1(new_n840), .B2(KEYINPUT57), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n615), .A3(new_n821), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT126), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n833), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n841), .A2(KEYINPUT126), .A3(new_n615), .A4(new_n821), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n835), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n819), .A2(new_n821), .ZN(new_n847));
  AOI211_X1 g646(.A(KEYINPUT59), .B(new_n833), .C1(new_n847), .C2(new_n615), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n834), .B1(new_n846), .B2(new_n848), .ZN(G1345gat));
  NAND2_X1  g648(.A1(new_n207), .A2(new_n212), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n639), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n812), .A2(new_n638), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n847), .A2(new_n851), .B1(new_n852), .B2(new_n850), .ZN(G1346gat));
  NAND2_X1  g652(.A1(new_n209), .A2(new_n211), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n519), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n812), .A2(new_n636), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n847), .A2(new_n855), .B1(new_n856), .B2(new_n854), .ZN(G1347gat));
  AND2_X1   g656(.A1(new_n774), .A2(new_n300), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n401), .A2(new_n451), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n379), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT127), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n326), .A3(new_n592), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n858), .A2(new_n777), .A3(new_n379), .ZN(new_n863));
  OAI21_X1  g662(.A(G169gat), .B1(new_n863), .B2(new_n593), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(G1348gat));
  NOR3_X1   g664(.A1(new_n863), .A2(new_n327), .A3(new_n694), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n861), .A2(new_n615), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(new_n327), .ZN(G1349gat));
  OAI21_X1  g667(.A(G183gat), .B1(new_n863), .B2(new_n639), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n858), .A2(new_n339), .A3(new_n379), .A4(new_n859), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n639), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g671(.A(G190gat), .B1(new_n863), .B2(new_n519), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT61), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n861), .A2(new_n315), .A3(new_n636), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1351gat));
  NOR2_X1   g675(.A1(new_n630), .A2(new_n380), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n300), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n815), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n584), .A3(new_n592), .ZN(new_n880));
  INV_X1    g679(.A(new_n841), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n881), .A2(new_n593), .A3(new_n878), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n880), .B1(new_n882), .B2(new_n584), .ZN(G1352gat));
  INV_X1    g682(.A(G204gat), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n879), .A2(new_n884), .A3(new_n615), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT62), .Z(new_n886));
  NOR3_X1   g685(.A1(new_n881), .A2(new_n694), .A3(new_n878), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n884), .ZN(G1353gat));
  NAND3_X1  g687(.A1(new_n879), .A2(new_n537), .A3(new_n638), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n841), .A2(new_n300), .A3(new_n638), .A4(new_n877), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n890), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT63), .B1(new_n890), .B2(G211gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(G1354gat));
  INV_X1    g692(.A(G218gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n879), .A2(new_n894), .A3(new_n636), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n881), .A2(new_n519), .A3(new_n878), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n894), .ZN(G1355gat));
endmodule


