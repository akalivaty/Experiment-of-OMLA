

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748;

  NOR2_X1 U380 ( .A1(KEYINPUT2), .A2(n736), .ZN(n665) );
  NOR2_X1 U381 ( .A1(n746), .A2(n745), .ZN(n600) );
  INV_X1 U382 ( .A(KEYINPUT41), .ZN(n360) );
  XNOR2_X1 U383 ( .A(n373), .B(n371), .ZN(n722) );
  BUF_X1 U384 ( .A(n485), .Z(n737) );
  XNOR2_X1 U385 ( .A(n448), .B(KEYINPUT68), .ZN(n506) );
  XNOR2_X1 U386 ( .A(n449), .B(G122), .ZN(n472) );
  XNOR2_X2 U387 ( .A(n361), .B(n360), .ZN(n703) );
  NAND2_X1 U388 ( .A1(n693), .A2(n689), .ZN(n361) );
  OR2_X2 U389 ( .A1(n706), .A2(n625), .ZN(n435) );
  NOR2_X1 U390 ( .A1(G902), .A2(n635), .ZN(n516) );
  XNOR2_X2 U391 ( .A(n484), .B(n439), .ZN(n455) );
  XNOR2_X2 U392 ( .A(n424), .B(G143), .ZN(n484) );
  XNOR2_X2 U393 ( .A(n376), .B(KEYINPUT32), .ZN(n744) );
  XNOR2_X2 U394 ( .A(n406), .B(n405), .ZN(n577) );
  XNOR2_X2 U395 ( .A(n548), .B(KEYINPUT99), .ZN(n691) );
  INV_X1 U396 ( .A(n614), .ZN(n535) );
  NAND2_X1 U397 ( .A1(n387), .A2(n389), .ZN(n502) );
  NAND2_X1 U398 ( .A1(n392), .A2(n386), .ZN(n551) );
  NAND2_X1 U399 ( .A1(n385), .A2(n391), .ZN(n388) );
  XNOR2_X1 U400 ( .A(n618), .B(n591), .ZN(n688) );
  XNOR2_X1 U401 ( .A(n681), .B(KEYINPUT6), .ZN(n604) );
  XNOR2_X1 U402 ( .A(n486), .B(n487), .ZN(n519) );
  XNOR2_X1 U403 ( .A(n399), .B(G953), .ZN(n485) );
  INV_X1 U404 ( .A(KEYINPUT64), .ZN(n399) );
  XOR2_X1 U405 ( .A(G125), .B(G146), .Z(n470) );
  XNOR2_X1 U406 ( .A(n408), .B(n407), .ZN(n704) );
  NOR2_X1 U407 ( .A1(G953), .A2(G237), .ZN(n507) );
  XOR2_X1 U408 ( .A(KEYINPUT67), .B(G131), .Z(n475) );
  INV_X1 U409 ( .A(KEYINPUT33), .ZN(n407) );
  NOR2_X1 U410 ( .A1(n549), .A2(n604), .ZN(n408) );
  XNOR2_X1 U411 ( .A(n526), .B(n527), .ZN(n405) );
  OR2_X1 U412 ( .A1(n713), .A2(G902), .ZN(n406) );
  NOR2_X1 U413 ( .A1(n671), .A2(n535), .ZN(n673) );
  NOR2_X1 U414 ( .A1(n637), .A2(n555), .ZN(n556) );
  NAND2_X1 U415 ( .A1(G237), .A2(G234), .ZN(n464) );
  XNOR2_X1 U416 ( .A(G140), .B(G143), .ZN(n476) );
  INV_X1 U417 ( .A(KEYINPUT0), .ZN(n393) );
  XNOR2_X1 U418 ( .A(n506), .B(n411), .ZN(n410) );
  XNOR2_X1 U419 ( .A(n505), .B(n508), .ZN(n409) );
  XNOR2_X1 U420 ( .A(n425), .B(n455), .ZN(n730) );
  XNOR2_X1 U421 ( .A(n440), .B(G134), .ZN(n425) );
  INV_X1 U422 ( .A(G128), .ZN(n424) );
  XNOR2_X1 U423 ( .A(n382), .B(KEYINPUT51), .ZN(n685) );
  OR2_X1 U424 ( .A1(n683), .A2(n684), .ZN(n382) );
  OR2_X1 U425 ( .A1(G902), .A2(G237), .ZN(n461) );
  XNOR2_X1 U426 ( .A(n423), .B(G469), .ZN(n575) );
  OR2_X1 U427 ( .A1(n503), .A2(G902), .ZN(n423) );
  NOR2_X1 U428 ( .A1(n688), .A2(n592), .ZN(n594) );
  XNOR2_X1 U429 ( .A(n481), .B(G475), .ZN(n482) );
  INV_X1 U430 ( .A(n577), .ZN(n675) );
  XNOR2_X1 U431 ( .A(n575), .B(n422), .ZN(n614) );
  INV_X1 U432 ( .A(KEYINPUT1), .ZN(n422) );
  XNOR2_X1 U433 ( .A(n404), .B(n403), .ZN(n524) );
  XNOR2_X1 U434 ( .A(n521), .B(n520), .ZN(n403) );
  NAND2_X1 U435 ( .A1(n519), .A2(G221), .ZN(n404) );
  INV_X1 U436 ( .A(KEYINPUT123), .ZN(n413) );
  OR2_X1 U437 ( .A1(n701), .A2(n365), .ZN(n402) );
  AND2_X1 U438 ( .A1(n601), .A2(n362), .ZN(n431) );
  INV_X1 U439 ( .A(KEYINPUT48), .ZN(n429) );
  NOR2_X1 U440 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U441 ( .A(G137), .B(G140), .Z(n522) );
  XNOR2_X1 U442 ( .A(n559), .B(n558), .ZN(n719) );
  XNOR2_X1 U443 ( .A(n509), .B(n441), .ZN(n453) );
  XNOR2_X1 U444 ( .A(G110), .B(KEYINPUT69), .ZN(n441) );
  XNOR2_X1 U445 ( .A(n522), .B(n381), .ZN(n442) );
  XNOR2_X1 U446 ( .A(G107), .B(G104), .ZN(n381) );
  INV_X1 U447 ( .A(KEYINPUT4), .ZN(n439) );
  XOR2_X1 U448 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n451) );
  XNOR2_X1 U449 ( .A(n596), .B(n380), .ZN(n693) );
  INV_X1 U450 ( .A(KEYINPUT105), .ZN(n380) );
  NOR2_X1 U451 ( .A1(n688), .A2(n687), .ZN(n596) );
  NOR2_X1 U452 ( .A1(n580), .A2(n606), .ZN(n582) );
  XNOR2_X1 U453 ( .A(n480), .B(n479), .ZN(n628) );
  NAND2_X1 U454 ( .A1(n585), .A2(n393), .ZN(n392) );
  NAND2_X1 U455 ( .A1(n469), .A2(n393), .ZN(n391) );
  INV_X1 U456 ( .A(n392), .ZN(n390) );
  AND2_X1 U457 ( .A1(n689), .A2(n499), .ZN(n500) );
  INV_X1 U458 ( .A(n674), .ZN(n499) );
  NAND2_X1 U459 ( .A1(n388), .A2(n500), .ZN(n387) );
  XNOR2_X1 U460 ( .A(n410), .B(n409), .ZN(n511) );
  XNOR2_X1 U461 ( .A(n490), .B(n372), .ZN(n371) );
  XNOR2_X1 U462 ( .A(n506), .B(n472), .ZN(n373) );
  INV_X1 U463 ( .A(KEYINPUT16), .ZN(n372) );
  BUF_X1 U464 ( .A(n719), .Z(n379) );
  XNOR2_X1 U465 ( .A(G128), .B(G110), .ZN(n517) );
  XOR2_X1 U466 ( .A(KEYINPUT24), .B(KEYINPUT93), .Z(n518) );
  XOR2_X1 U467 ( .A(KEYINPUT23), .B(G119), .Z(n520) );
  XOR2_X1 U468 ( .A(G134), .B(G122), .Z(n437) );
  XNOR2_X1 U469 ( .A(n699), .B(n384), .ZN(n383) );
  INV_X1 U470 ( .A(KEYINPUT52), .ZN(n384) );
  NOR2_X1 U471 ( .A1(n606), .A2(n605), .ZN(n613) );
  OR2_X1 U472 ( .A1(n638), .A2(n604), .ZN(n605) );
  XNOR2_X1 U473 ( .A(n460), .B(n434), .ZN(n433) );
  INV_X1 U474 ( .A(KEYINPUT88), .ZN(n434) );
  XNOR2_X1 U475 ( .A(n599), .B(KEYINPUT42), .ZN(n745) );
  NOR2_X1 U476 ( .A1(n703), .A2(n598), .ZN(n599) );
  NAND2_X1 U477 ( .A1(n421), .A2(n571), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n537), .B(n536), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n545), .B(KEYINPUT98), .ZN(n647) );
  AND2_X1 U480 ( .A1(n531), .A2(n364), .ZN(n528) );
  XNOR2_X1 U481 ( .A(n414), .B(n412), .ZN(n714) );
  XNOR2_X1 U482 ( .A(n713), .B(n413), .ZN(n412) );
  INV_X1 U483 ( .A(KEYINPUT56), .ZN(n394) );
  INV_X1 U484 ( .A(KEYINPUT53), .ZN(n426) );
  AND2_X1 U485 ( .A1(n610), .A2(n663), .ZN(n362) );
  OR2_X1 U486 ( .A1(n469), .A2(n393), .ZN(n363) );
  XNOR2_X1 U487 ( .A(n483), .B(n482), .ZN(n543) );
  AND2_X1 U488 ( .A1(n614), .A2(n580), .ZN(n364) );
  AND2_X1 U489 ( .A1(n705), .A2(n704), .ZN(n365) );
  XNOR2_X1 U490 ( .A(n635), .B(n634), .ZN(n366) );
  XNOR2_X1 U491 ( .A(KEYINPUT35), .B(KEYINPUT79), .ZN(n367) );
  XOR2_X1 U492 ( .A(n708), .B(n707), .Z(n368) );
  XOR2_X1 U493 ( .A(n633), .B(KEYINPUT65), .Z(n369) );
  XOR2_X1 U494 ( .A(KEYINPUT63), .B(KEYINPUT107), .Z(n370) );
  INV_X1 U495 ( .A(n715), .ZN(n396) );
  NAND2_X1 U496 ( .A1(n712), .A2(G469), .ZN(n417) );
  NOR2_X4 U497 ( .A1(n669), .A2(n626), .ZN(n712) );
  NAND2_X1 U498 ( .A1(n390), .A2(n500), .ZN(n389) );
  NOR2_X2 U499 ( .A1(n702), .A2(n402), .ZN(n401) );
  XNOR2_X1 U500 ( .A(n600), .B(KEYINPUT46), .ZN(n432) );
  XNOR2_X1 U501 ( .A(n374), .B(n369), .ZN(G60) );
  NAND2_X1 U502 ( .A1(n378), .A2(n396), .ZN(n374) );
  XNOR2_X1 U503 ( .A(n375), .B(n370), .ZN(G57) );
  NAND2_X1 U504 ( .A1(n377), .A2(n396), .ZN(n375) );
  INV_X1 U505 ( .A(n742), .ZN(n620) );
  XNOR2_X1 U506 ( .A(n619), .B(KEYINPUT101), .ZN(n742) );
  XNOR2_X1 U507 ( .A(n504), .B(KEYINPUT75), .ZN(n411) );
  NAND2_X1 U508 ( .A1(n531), .A2(n532), .ZN(n376) );
  XNOR2_X1 U509 ( .A(n636), .B(n366), .ZN(n377) );
  XNOR2_X1 U510 ( .A(n632), .B(n631), .ZN(n378) );
  AND2_X2 U511 ( .A1(n618), .A2(n463), .ZN(n607) );
  NAND2_X1 U512 ( .A1(n744), .A2(n646), .ZN(n534) );
  NAND2_X1 U513 ( .A1(n557), .A2(n556), .ZN(n559) );
  XNOR2_X1 U514 ( .A(n513), .B(n445), .ZN(n503) );
  NOR2_X1 U515 ( .A1(n383), .A2(n700), .ZN(n701) );
  NAND2_X1 U516 ( .A1(n531), .A2(n614), .ZN(n542) );
  OR2_X2 U517 ( .A1(n585), .A2(n363), .ZN(n385) );
  XNOR2_X2 U518 ( .A(n607), .B(KEYINPUT19), .ZN(n585) );
  INV_X1 U519 ( .A(n388), .ZN(n386) );
  XNOR2_X1 U520 ( .A(n395), .B(n394), .ZN(G51) );
  NAND2_X1 U521 ( .A1(n397), .A2(n396), .ZN(n395) );
  XNOR2_X1 U522 ( .A(n398), .B(n368), .ZN(n397) );
  NAND2_X1 U523 ( .A1(n712), .A2(G210), .ZN(n398) );
  NAND2_X1 U524 ( .A1(n400), .A2(n428), .ZN(n427) );
  XNOR2_X1 U525 ( .A(n401), .B(KEYINPUT118), .ZN(n400) );
  NAND2_X1 U526 ( .A1(n704), .A2(n551), .ZN(n537) );
  NAND2_X1 U527 ( .A1(n712), .A2(G217), .ZN(n414) );
  XNOR2_X2 U528 ( .A(n502), .B(n501), .ZN(n531) );
  NOR2_X2 U529 ( .A1(n719), .A2(n664), .ZN(n624) );
  NAND2_X1 U530 ( .A1(n432), .A2(n431), .ZN(n430) );
  NOR2_X2 U531 ( .A1(n674), .A2(n675), .ZN(n671) );
  AND2_X2 U532 ( .A1(n624), .A2(KEYINPUT2), .ZN(n623) );
  XNOR2_X1 U533 ( .A(n430), .B(n429), .ZN(n622) );
  XNOR2_X2 U534 ( .A(n623), .B(KEYINPUT76), .ZN(n669) );
  XNOR2_X1 U535 ( .A(n415), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U536 ( .A1(n416), .A2(n396), .ZN(n415) );
  XNOR2_X1 U537 ( .A(n417), .B(n627), .ZN(n416) );
  NAND2_X1 U538 ( .A1(n419), .A2(n418), .ZN(n539) );
  INV_X1 U539 ( .A(KEYINPUT44), .ZN(n418) );
  INV_X1 U540 ( .A(n743), .ZN(n419) );
  XNOR2_X2 U541 ( .A(n420), .B(n367), .ZN(n743) );
  XNOR2_X1 U542 ( .A(n427), .B(n426), .ZN(G75) );
  INV_X1 U543 ( .A(G953), .ZN(n428) );
  XNOR2_X2 U544 ( .A(n435), .B(n433), .ZN(n618) );
  XNOR2_X2 U545 ( .A(G119), .B(KEYINPUT3), .ZN(n448) );
  XNOR2_X2 U546 ( .A(G104), .B(G113), .ZN(n449) );
  XNOR2_X1 U547 ( .A(n490), .B(n437), .ZN(n491) );
  XOR2_X1 U548 ( .A(n477), .B(n476), .Z(n436) );
  OR2_X1 U549 ( .A1(n624), .A2(KEYINPUT2), .ZN(n438) );
  INV_X1 U550 ( .A(n691), .ZN(n692) );
  XNOR2_X1 U551 ( .A(n478), .B(n436), .ZN(n479) );
  INV_X1 U552 ( .A(KEYINPUT13), .ZN(n481) );
  INV_X1 U553 ( .A(n687), .ZN(n463) );
  XNOR2_X1 U554 ( .A(n514), .B(G472), .ZN(n515) );
  INV_X1 U555 ( .A(KEYINPUT45), .ZN(n558) );
  NAND2_X1 U556 ( .A1(n438), .A2(n625), .ZN(n626) );
  XNOR2_X1 U557 ( .A(KEYINPUT84), .B(KEYINPUT39), .ZN(n593) );
  NAND2_X1 U558 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U559 ( .A1(n737), .A2(G952), .ZN(n715) );
  XNOR2_X1 U560 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n447) );
  INV_X1 U561 ( .A(n475), .ZN(n440) );
  XNOR2_X1 U562 ( .A(G146), .B(n730), .ZN(n513) );
  XOR2_X1 U563 ( .A(G101), .B(KEYINPUT66), .Z(n509) );
  XOR2_X1 U564 ( .A(n453), .B(n442), .Z(n444) );
  NAND2_X1 U565 ( .A1(G227), .A2(n737), .ZN(n443) );
  XNOR2_X1 U566 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U567 ( .A(n503), .B(KEYINPUT57), .ZN(n446) );
  XNOR2_X1 U568 ( .A(n447), .B(n446), .ZN(n627) );
  XOR2_X1 U569 ( .A(G107), .B(G116), .Z(n490) );
  NAND2_X1 U570 ( .A1(G224), .A2(n737), .ZN(n450) );
  XOR2_X1 U571 ( .A(n451), .B(n450), .Z(n452) );
  XNOR2_X1 U572 ( .A(n722), .B(n452), .ZN(n459) );
  INV_X1 U573 ( .A(KEYINPUT78), .ZN(n454) );
  XNOR2_X1 U574 ( .A(n454), .B(n453), .ZN(n457) );
  XNOR2_X1 U575 ( .A(n470), .B(n455), .ZN(n456) );
  XNOR2_X1 U576 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U577 ( .A(n459), .B(n458), .ZN(n706) );
  XOR2_X1 U578 ( .A(KEYINPUT15), .B(G902), .Z(n625) );
  NAND2_X1 U579 ( .A1(G210), .A2(n461), .ZN(n460) );
  NAND2_X1 U580 ( .A1(G214), .A2(n461), .ZN(n462) );
  XNOR2_X1 U581 ( .A(KEYINPUT89), .B(n462), .ZN(n687) );
  XNOR2_X1 U582 ( .A(n464), .B(KEYINPUT90), .ZN(n465) );
  XNOR2_X1 U583 ( .A(KEYINPUT14), .B(n465), .ZN(n467) );
  NAND2_X1 U584 ( .A1(G952), .A2(n467), .ZN(n700) );
  NOR2_X1 U585 ( .A1(G953), .A2(n700), .ZN(n466) );
  XOR2_X1 U586 ( .A(KEYINPUT91), .B(n466), .Z(n564) );
  NAND2_X1 U587 ( .A1(G902), .A2(n467), .ZN(n565) );
  XOR2_X1 U588 ( .A(G898), .B(KEYINPUT92), .Z(n718) );
  NAND2_X1 U589 ( .A1(G953), .A2(n718), .ZN(n725) );
  NOR2_X1 U590 ( .A1(n565), .A2(n725), .ZN(n468) );
  NOR2_X1 U591 ( .A1(n564), .A2(n468), .ZN(n469) );
  INV_X1 U592 ( .A(n470), .ZN(n471) );
  XNOR2_X1 U593 ( .A(KEYINPUT10), .B(n471), .ZN(n523) );
  XOR2_X1 U594 ( .A(n472), .B(n523), .Z(n474) );
  NAND2_X1 U595 ( .A1(n507), .A2(G214), .ZN(n473) );
  XNOR2_X1 U596 ( .A(n474), .B(n473), .ZN(n480) );
  XNOR2_X1 U597 ( .A(n475), .B(KEYINPUT12), .ZN(n478) );
  XOR2_X1 U598 ( .A(KEYINPUT11), .B(KEYINPUT96), .Z(n477) );
  NOR2_X1 U599 ( .A1(G902), .A2(n628), .ZN(n483) );
  XOR2_X1 U600 ( .A(n484), .B(KEYINPUT97), .Z(n489) );
  XOR2_X1 U601 ( .A(KEYINPUT82), .B(KEYINPUT8), .Z(n487) );
  NAND2_X1 U602 ( .A1(n485), .A2(G234), .ZN(n486) );
  NAND2_X1 U603 ( .A1(G217), .A2(n519), .ZN(n488) );
  XNOR2_X1 U604 ( .A(n489), .B(n488), .ZN(n492) );
  XNOR2_X1 U605 ( .A(n492), .B(n491), .ZN(n494) );
  XOR2_X1 U606 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n493) );
  XNOR2_X1 U607 ( .A(n494), .B(n493), .ZN(n710) );
  NOR2_X1 U608 ( .A1(G902), .A2(n710), .ZN(n495) );
  XNOR2_X1 U609 ( .A(G478), .B(n495), .ZN(n546) );
  AND2_X1 U610 ( .A1(n543), .A2(n546), .ZN(n689) );
  INV_X1 U611 ( .A(n625), .ZN(n496) );
  NAND2_X1 U612 ( .A1(G234), .A2(n496), .ZN(n497) );
  XNOR2_X1 U613 ( .A(KEYINPUT20), .B(n497), .ZN(n525) );
  NAND2_X1 U614 ( .A1(n525), .A2(G221), .ZN(n498) );
  XNOR2_X1 U615 ( .A(n498), .B(KEYINPUT21), .ZN(n674) );
  XNOR2_X1 U616 ( .A(KEYINPUT22), .B(KEYINPUT72), .ZN(n501) );
  XOR2_X1 U617 ( .A(G113), .B(G116), .Z(n505) );
  XNOR2_X1 U618 ( .A(KEYINPUT5), .B(KEYINPUT94), .ZN(n504) );
  AND2_X1 U619 ( .A1(n507), .A2(G210), .ZN(n508) );
  XOR2_X1 U620 ( .A(G137), .B(n509), .Z(n510) );
  XNOR2_X1 U621 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U622 ( .A(n512), .B(n513), .ZN(n635) );
  XNOR2_X1 U623 ( .A(KEYINPUT71), .B(KEYINPUT95), .ZN(n514) );
  XNOR2_X2 U624 ( .A(n516), .B(n515), .ZN(n580) );
  INV_X1 U625 ( .A(n580), .ZN(n681) );
  XNOR2_X1 U626 ( .A(KEYINPUT25), .B(KEYINPUT77), .ZN(n527) );
  XNOR2_X1 U627 ( .A(n518), .B(n517), .ZN(n521) );
  XNOR2_X1 U628 ( .A(n523), .B(n522), .ZN(n731) );
  XNOR2_X1 U629 ( .A(n524), .B(n731), .ZN(n713) );
  NAND2_X1 U630 ( .A1(G217), .A2(n525), .ZN(n526) );
  NAND2_X1 U631 ( .A1(n528), .A2(n675), .ZN(n646) );
  NAND2_X1 U632 ( .A1(n535), .A2(n604), .ZN(n529) );
  NOR2_X1 U633 ( .A1(n577), .A2(n529), .ZN(n530) );
  XNOR2_X1 U634 ( .A(KEYINPUT80), .B(n530), .ZN(n532) );
  NOR2_X1 U635 ( .A1(KEYINPUT44), .A2(KEYINPUT85), .ZN(n533) );
  XNOR2_X1 U636 ( .A(n534), .B(n533), .ZN(n538) );
  NAND2_X1 U637 ( .A1(n671), .A2(n535), .ZN(n549) );
  XOR2_X1 U638 ( .A(KEYINPUT70), .B(KEYINPUT34), .Z(n536) );
  NOR2_X1 U639 ( .A1(n543), .A2(n546), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n538), .A2(n743), .ZN(n540) );
  NAND2_X1 U641 ( .A1(n540), .A2(n539), .ZN(n557) );
  NAND2_X1 U642 ( .A1(n577), .A2(n604), .ZN(n541) );
  NOR2_X1 U643 ( .A1(n542), .A2(n541), .ZN(n637) );
  INV_X1 U644 ( .A(n546), .ZN(n544) );
  INV_X1 U645 ( .A(n543), .ZN(n547) );
  NAND2_X1 U646 ( .A1(n547), .A2(n546), .ZN(n638) );
  NAND2_X1 U647 ( .A1(n647), .A2(n638), .ZN(n548) );
  NOR2_X1 U648 ( .A1(n580), .A2(n549), .ZN(n684) );
  NAND2_X1 U649 ( .A1(n551), .A2(n684), .ZN(n550) );
  XNOR2_X1 U650 ( .A(n550), .B(KEYINPUT31), .ZN(n659) );
  NAND2_X1 U651 ( .A1(n671), .A2(n575), .ZN(n563) );
  NAND2_X1 U652 ( .A1(n580), .A2(n551), .ZN(n552) );
  NOR2_X1 U653 ( .A1(n563), .A2(n552), .ZN(n641) );
  NOR2_X1 U654 ( .A1(n659), .A2(n641), .ZN(n553) );
  NOR2_X1 U655 ( .A1(n691), .A2(n553), .ZN(n554) );
  XNOR2_X1 U656 ( .A(n554), .B(KEYINPUT100), .ZN(n555) );
  INV_X1 U657 ( .A(KEYINPUT30), .ZN(n561) );
  NOR2_X1 U658 ( .A1(n687), .A2(n580), .ZN(n560) );
  XNOR2_X1 U659 ( .A(n561), .B(n560), .ZN(n562) );
  NOR2_X1 U660 ( .A1(n563), .A2(n562), .ZN(n570) );
  INV_X1 U661 ( .A(n564), .ZN(n569) );
  NOR2_X1 U662 ( .A1(G900), .A2(n565), .ZN(n567) );
  INV_X1 U663 ( .A(n737), .ZN(n566) );
  NAND2_X1 U664 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U665 ( .A1(n569), .A2(n568), .ZN(n578) );
  NAND2_X1 U666 ( .A1(n570), .A2(n578), .ZN(n592) );
  INV_X1 U667 ( .A(n592), .ZN(n573) );
  AND2_X1 U668 ( .A1(n618), .A2(n571), .ZN(n572) );
  NAND2_X1 U669 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U670 ( .A(KEYINPUT102), .B(n574), .ZN(n748) );
  XNOR2_X1 U671 ( .A(KEYINPUT81), .B(n748), .ZN(n590) );
  INV_X1 U672 ( .A(n575), .ZN(n576) );
  XNOR2_X1 U673 ( .A(KEYINPUT103), .B(n576), .ZN(n584) );
  NOR2_X1 U674 ( .A1(n674), .A2(n577), .ZN(n579) );
  NAND2_X1 U675 ( .A1(n579), .A2(n578), .ZN(n606) );
  XNOR2_X1 U676 ( .A(KEYINPUT28), .B(KEYINPUT104), .ZN(n581) );
  XNOR2_X1 U677 ( .A(n582), .B(n581), .ZN(n583) );
  NAND2_X1 U678 ( .A1(n584), .A2(n583), .ZN(n598) );
  NOR2_X1 U679 ( .A1(n598), .A2(n585), .ZN(n653) );
  INV_X1 U680 ( .A(n653), .ZN(n648) );
  XNOR2_X1 U681 ( .A(n691), .B(KEYINPUT73), .ZN(n587) );
  INV_X1 U682 ( .A(KEYINPUT47), .ZN(n586) );
  NAND2_X1 U683 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U684 ( .A1(n648), .A2(n588), .ZN(n589) );
  NOR2_X1 U685 ( .A1(n590), .A2(n589), .ZN(n601) );
  XNOR2_X1 U686 ( .A(KEYINPUT74), .B(KEYINPUT38), .ZN(n591) );
  XNOR2_X1 U687 ( .A(n594), .B(n593), .ZN(n611) );
  NOR2_X1 U688 ( .A1(n638), .A2(n611), .ZN(n595) );
  XNOR2_X1 U689 ( .A(n595), .B(KEYINPUT40), .ZN(n746) );
  NOR2_X1 U690 ( .A1(n691), .A2(KEYINPUT73), .ZN(n602) );
  NAND2_X1 U691 ( .A1(n602), .A2(n653), .ZN(n603) );
  NAND2_X1 U692 ( .A1(n603), .A2(KEYINPUT47), .ZN(n610) );
  AND2_X1 U693 ( .A1(n607), .A2(n613), .ZN(n608) );
  XNOR2_X1 U694 ( .A(n608), .B(KEYINPUT36), .ZN(n609) );
  NAND2_X1 U695 ( .A1(n609), .A2(n535), .ZN(n663) );
  NOR2_X1 U696 ( .A1(n647), .A2(n611), .ZN(n612) );
  XNOR2_X1 U697 ( .A(n612), .B(KEYINPUT106), .ZN(n747) );
  NAND2_X1 U698 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U699 ( .A1(n687), .A2(n615), .ZN(n616) );
  XNOR2_X1 U700 ( .A(n616), .B(KEYINPUT43), .ZN(n617) );
  NOR2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U702 ( .A1(n747), .A2(n620), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n622), .A2(n621), .ZN(n664) );
  NAND2_X1 U704 ( .A1(n712), .A2(G475), .ZN(n632) );
  XOR2_X1 U705 ( .A(KEYINPUT87), .B(KEYINPUT59), .Z(n630) );
  XNOR2_X1 U706 ( .A(n628), .B(KEYINPUT122), .ZN(n629) );
  XNOR2_X1 U707 ( .A(n630), .B(n629), .ZN(n631) );
  INV_X1 U708 ( .A(KEYINPUT60), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n712), .A2(G472), .ZN(n636) );
  XOR2_X1 U710 ( .A(KEYINPUT62), .B(KEYINPUT86), .Z(n634) );
  XOR2_X1 U711 ( .A(G101), .B(n637), .Z(G3) );
  INV_X1 U712 ( .A(n638), .ZN(n656) );
  NAND2_X1 U713 ( .A1(n641), .A2(n656), .ZN(n639) );
  XNOR2_X1 U714 ( .A(n639), .B(KEYINPUT108), .ZN(n640) );
  XNOR2_X1 U715 ( .A(G104), .B(n640), .ZN(G6) );
  XOR2_X1 U716 ( .A(KEYINPUT109), .B(KEYINPUT26), .Z(n643) );
  INV_X1 U717 ( .A(n647), .ZN(n658) );
  NAND2_X1 U718 ( .A1(n641), .A2(n658), .ZN(n642) );
  XNOR2_X1 U719 ( .A(n643), .B(n642), .ZN(n645) );
  XOR2_X1 U720 ( .A(G107), .B(KEYINPUT27), .Z(n644) );
  XNOR2_X1 U721 ( .A(n645), .B(n644), .ZN(G9) );
  XNOR2_X1 U722 ( .A(n646), .B(G110), .ZN(G12) );
  NOR2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n652) );
  XOR2_X1 U724 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n650) );
  XNOR2_X1 U725 ( .A(G128), .B(KEYINPUT29), .ZN(n649) );
  XNOR2_X1 U726 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n652), .B(n651), .ZN(G30) );
  NAND2_X1 U728 ( .A1(n653), .A2(n656), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n654), .B(KEYINPUT112), .ZN(n655) );
  XNOR2_X1 U730 ( .A(G146), .B(n655), .ZN(G48) );
  NAND2_X1 U731 ( .A1(n656), .A2(n659), .ZN(n657) );
  XNOR2_X1 U732 ( .A(G113), .B(n657), .ZN(G15) );
  XOR2_X1 U733 ( .A(G116), .B(KEYINPUT113), .Z(n661) );
  NAND2_X1 U734 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U735 ( .A(n661), .B(n660), .ZN(G18) );
  XOR2_X1 U736 ( .A(G125), .B(KEYINPUT37), .Z(n662) );
  XNOR2_X1 U737 ( .A(n663), .B(n662), .ZN(G27) );
  INV_X1 U738 ( .A(n664), .ZN(n736) );
  XNOR2_X1 U739 ( .A(n665), .B(KEYINPUT83), .ZN(n668) );
  INV_X1 U740 ( .A(KEYINPUT2), .ZN(n666) );
  NAND2_X1 U741 ( .A1(n666), .A2(n379), .ZN(n667) );
  NAND2_X1 U742 ( .A1(n668), .A2(n667), .ZN(n670) );
  NOR2_X1 U743 ( .A1(n670), .A2(n669), .ZN(n702) );
  XNOR2_X1 U744 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n672) );
  XNOR2_X1 U745 ( .A(n673), .B(n672), .ZN(n679) );
  XOR2_X1 U746 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n677) );
  NAND2_X1 U747 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U748 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U750 ( .A(n682), .B(KEYINPUT116), .ZN(n683) );
  NOR2_X1 U751 ( .A1(n703), .A2(n685), .ZN(n686) );
  XNOR2_X1 U752 ( .A(n686), .B(KEYINPUT117), .ZN(n698) );
  NAND2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n690) );
  NAND2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n695) );
  NAND2_X1 U755 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U756 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U757 ( .A1(n704), .A2(n696), .ZN(n697) );
  NAND2_X1 U758 ( .A1(n698), .A2(n697), .ZN(n699) );
  INV_X1 U759 ( .A(n703), .ZN(n705) );
  XNOR2_X1 U760 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n708) );
  XNOR2_X1 U761 ( .A(n706), .B(KEYINPUT55), .ZN(n707) );
  NAND2_X1 U762 ( .A1(G478), .A2(n712), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n715), .A2(n711), .ZN(G63) );
  NOR2_X1 U765 ( .A1(n715), .A2(n714), .ZN(G66) );
  NAND2_X1 U766 ( .A1(G953), .A2(G224), .ZN(n716) );
  XOR2_X1 U767 ( .A(KEYINPUT61), .B(n716), .Z(n717) );
  NOR2_X1 U768 ( .A1(n718), .A2(n717), .ZN(n721) );
  NOR2_X1 U769 ( .A1(G953), .A2(n379), .ZN(n720) );
  NOR2_X1 U770 ( .A1(n721), .A2(n720), .ZN(n729) );
  XNOR2_X1 U771 ( .A(n722), .B(G101), .ZN(n723) );
  XNOR2_X1 U772 ( .A(n723), .B(KEYINPUT125), .ZN(n724) );
  XNOR2_X1 U773 ( .A(G110), .B(n724), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U775 ( .A(n727), .B(KEYINPUT124), .ZN(n728) );
  XNOR2_X1 U776 ( .A(n729), .B(n728), .ZN(G69) );
  XNOR2_X1 U777 ( .A(n731), .B(n730), .ZN(n735) );
  XOR2_X1 U778 ( .A(G227), .B(n735), .Z(n732) );
  NAND2_X1 U779 ( .A1(n732), .A2(G900), .ZN(n733) );
  XNOR2_X1 U780 ( .A(n733), .B(KEYINPUT126), .ZN(n734) );
  NAND2_X1 U781 ( .A1(n734), .A2(G953), .ZN(n740) );
  XNOR2_X1 U782 ( .A(n736), .B(n735), .ZN(n738) );
  NAND2_X1 U783 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U784 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U785 ( .A(KEYINPUT127), .B(n741), .Z(G72) );
  XNOR2_X1 U786 ( .A(G140), .B(n742), .ZN(G42) );
  XNOR2_X1 U787 ( .A(G122), .B(n743), .ZN(G24) );
  XNOR2_X1 U788 ( .A(n744), .B(G119), .ZN(G21) );
  XOR2_X1 U789 ( .A(n745), .B(G137), .Z(G39) );
  XOR2_X1 U790 ( .A(G131), .B(n746), .Z(G33) );
  XOR2_X1 U791 ( .A(G134), .B(n747), .Z(G36) );
  XNOR2_X1 U792 ( .A(G143), .B(n748), .ZN(G45) );
endmodule

