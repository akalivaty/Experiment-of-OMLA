

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745;

  XNOR2_X1 U378 ( .A(n400), .B(G110), .ZN(n402) );
  INV_X2 U379 ( .A(G953), .ZN(n738) );
  AND2_X2 U380 ( .A1(n363), .A2(n362), .ZN(n366) );
  AND2_X4 U381 ( .A1(n608), .A2(n607), .ZN(n637) );
  NAND2_X2 U382 ( .A1(n488), .A2(n533), .ZN(n517) );
  XNOR2_X2 U383 ( .A(n592), .B(KEYINPUT103), .ZN(n618) );
  XNOR2_X2 U384 ( .A(n408), .B(n407), .ZN(n504) );
  NOR2_X1 U385 ( .A1(n616), .A2(KEYINPUT44), .ZN(n582) );
  AND2_X1 U386 ( .A1(n573), .A2(n572), .ZN(n581) );
  NOR2_X1 U387 ( .A1(n588), .A2(n587), .ZN(n589) );
  AND2_X2 U388 ( .A1(n622), .A2(n644), .ZN(n624) );
  AND2_X2 U389 ( .A1(n634), .A2(n644), .ZN(n636) );
  AND2_X2 U390 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U391 ( .A1(n736), .A2(n718), .ZN(n669) );
  XNOR2_X1 U392 ( .A(KEYINPUT4), .B(G101), .ZN(n464) );
  XOR2_X1 U393 ( .A(KEYINPUT89), .B(KEYINPUT75), .Z(n462) );
  XNOR2_X1 U394 ( .A(KEYINPUT88), .B(KEYINPUT17), .ZN(n463) );
  XNOR2_X1 U395 ( .A(n474), .B(KEYINPUT90), .ZN(n475) );
  OR2_X2 U396 ( .A1(n588), .A2(n569), .ZN(n368) );
  XNOR2_X1 U397 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U398 ( .A(G128), .B(G110), .ZN(n409) );
  XNOR2_X1 U399 ( .A(n500), .B(n499), .ZN(n711) );
  XNOR2_X1 U400 ( .A(n494), .B(KEYINPUT39), .ZN(n531) );
  AND2_X1 U401 ( .A1(n529), .A2(n355), .ZN(n530) );
  INV_X1 U402 ( .A(KEYINPUT104), .ZN(n603) );
  XNOR2_X1 U403 ( .A(n498), .B(KEYINPUT109), .ZN(n682) );
  XNOR2_X1 U404 ( .A(G122), .B(G107), .ZN(n445) );
  NAND2_X1 U405 ( .A1(n669), .A2(n374), .ZN(n370) );
  NAND2_X1 U406 ( .A1(n605), .A2(n374), .ZN(n373) );
  NAND2_X1 U407 ( .A1(n375), .A2(KEYINPUT2), .ZN(n372) );
  INV_X1 U408 ( .A(G146), .ZN(n387) );
  XNOR2_X1 U409 ( .A(n724), .B(n472), .ZN(n638) );
  NOR2_X1 U410 ( .A1(n669), .A2(n606), .ZN(n673) );
  NOR2_X1 U411 ( .A1(n481), .A2(n425), .ZN(n493) );
  XNOR2_X1 U412 ( .A(n397), .B(n396), .ZN(n424) );
  XNOR2_X1 U413 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n396) );
  XNOR2_X1 U414 ( .A(n368), .B(n570), .ZN(n573) );
  XNOR2_X1 U415 ( .A(n731), .B(n411), .ZN(n418) );
  NOR2_X1 U416 ( .A1(n711), .A2(n506), .ZN(n507) );
  AND2_X1 U417 ( .A1(n370), .A2(n357), .ZN(n354) );
  AND2_X1 U418 ( .A1(n528), .A2(n376), .ZN(n355) );
  XOR2_X1 U419 ( .A(KEYINPUT72), .B(KEYINPUT22), .Z(n356) );
  AND2_X1 U420 ( .A1(n373), .A2(n372), .ZN(n357) );
  XOR2_X1 U421 ( .A(n610), .B(n609), .Z(n358) );
  XOR2_X1 U422 ( .A(n632), .B(n631), .Z(n359) );
  XNOR2_X1 U423 ( .A(n620), .B(KEYINPUT62), .ZN(n360) );
  XOR2_X1 U424 ( .A(n639), .B(n641), .Z(n361) );
  XNOR2_X1 U425 ( .A(G902), .B(KEYINPUT15), .ZN(n605) );
  NOR2_X1 U426 ( .A1(n738), .A2(G952), .ZN(n643) );
  INV_X1 U427 ( .A(KEYINPUT84), .ZN(n374) );
  NAND2_X1 U428 ( .A1(n579), .A2(n578), .ZN(n362) );
  NAND2_X1 U429 ( .A1(n585), .A2(n584), .ZN(n363) );
  XNOR2_X2 U430 ( .A(n364), .B(KEYINPUT45), .ZN(n718) );
  NAND2_X2 U431 ( .A1(n366), .A2(n365), .ZN(n364) );
  XNOR2_X2 U432 ( .A(n367), .B(n603), .ZN(n365) );
  NAND2_X1 U433 ( .A1(n618), .A2(n602), .ZN(n367) );
  XNOR2_X2 U434 ( .A(n369), .B(n356), .ZN(n588) );
  NOR2_X2 U435 ( .A1(n594), .A2(n565), .ZN(n369) );
  NAND2_X1 U436 ( .A1(n371), .A2(n354), .ZN(n608) );
  NAND2_X1 U437 ( .A1(n604), .A2(n375), .ZN(n371) );
  INV_X1 U438 ( .A(n605), .ZN(n375) );
  NOR2_X2 U439 ( .A1(n591), .A2(n590), .ZN(n592) );
  OR2_X1 U440 ( .A1(n527), .A2(n526), .ZN(n376) );
  AND2_X1 U441 ( .A1(G217), .A2(n422), .ZN(n377) );
  INV_X1 U442 ( .A(n742), .ZN(n509) );
  INV_X1 U443 ( .A(G902), .ZN(n452) );
  AND2_X1 U444 ( .A1(n543), .A2(n542), .ZN(n736) );
  INV_X1 U445 ( .A(n581), .ZN(n617) );
  NOR2_X1 U446 ( .A1(G900), .A2(n738), .ZN(n378) );
  NAND2_X1 U447 ( .A1(n378), .A2(G902), .ZN(n379) );
  NAND2_X1 U448 ( .A1(n738), .A2(G952), .ZN(n548) );
  NAND2_X1 U449 ( .A1(n379), .A2(n548), .ZN(n381) );
  NAND2_X1 U450 ( .A1(G234), .A2(G237), .ZN(n380) );
  XNOR2_X1 U451 ( .A(n380), .B(KEYINPUT14), .ZN(n676) );
  NAND2_X1 U452 ( .A1(n381), .A2(n676), .ZN(n481) );
  NOR2_X1 U453 ( .A1(G902), .A2(G237), .ZN(n382) );
  XNOR2_X1 U454 ( .A(KEYINPUT73), .B(n382), .ZN(n473) );
  NAND2_X1 U455 ( .A1(n473), .A2(G214), .ZN(n384) );
  INV_X1 U456 ( .A(KEYINPUT91), .ZN(n383) );
  XNOR2_X1 U457 ( .A(n384), .B(n383), .ZN(n533) );
  XOR2_X1 U458 ( .A(G137), .B(KEYINPUT5), .Z(n386) );
  NOR2_X1 U459 ( .A1(G953), .A2(G237), .ZN(n432) );
  NAND2_X1 U460 ( .A1(n432), .A2(G210), .ZN(n385) );
  XNOR2_X1 U461 ( .A(n386), .B(n385), .ZN(n388) );
  XNOR2_X1 U462 ( .A(n464), .B(n387), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n388), .B(n404), .ZN(n392) );
  XNOR2_X1 U464 ( .A(G119), .B(G116), .ZN(n389) );
  XNOR2_X1 U465 ( .A(n389), .B(KEYINPUT3), .ZN(n391) );
  XNOR2_X1 U466 ( .A(G113), .B(KEYINPUT71), .ZN(n390) );
  XNOR2_X1 U467 ( .A(n391), .B(n390), .ZN(n458) );
  XNOR2_X1 U468 ( .A(n392), .B(n458), .ZN(n394) );
  XNOR2_X1 U469 ( .A(G131), .B(KEYINPUT68), .ZN(n393) );
  XNOR2_X1 U470 ( .A(n393), .B(KEYINPUT67), .ZN(n429) );
  XNOR2_X2 U471 ( .A(G143), .B(G128), .ZN(n460) );
  XNOR2_X1 U472 ( .A(n460), .B(G134), .ZN(n448) );
  XOR2_X1 U473 ( .A(n429), .B(n448), .Z(n399) );
  XNOR2_X1 U474 ( .A(n394), .B(n399), .ZN(n620) );
  NAND2_X1 U475 ( .A1(n620), .A2(n452), .ZN(n395) );
  XNOR2_X1 U476 ( .A(n395), .B(G472), .ZN(n501) );
  NAND2_X1 U477 ( .A1(n533), .A2(n501), .ZN(n397) );
  XOR2_X1 U478 ( .A(G137), .B(G140), .Z(n410) );
  INV_X1 U479 ( .A(n410), .ZN(n398) );
  XNOR2_X1 U480 ( .A(n399), .B(n398), .ZN(n730) );
  INV_X2 U481 ( .A(KEYINPUT74), .ZN(n400) );
  XNOR2_X1 U482 ( .A(G107), .B(G104), .ZN(n401) );
  XNOR2_X1 U483 ( .A(n402), .B(n401), .ZN(n455) );
  NAND2_X1 U484 ( .A1(G227), .A2(n738), .ZN(n403) );
  XNOR2_X1 U485 ( .A(n455), .B(n403), .ZN(n405) );
  XNOR2_X1 U486 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U487 ( .A(n730), .B(n406), .ZN(n610) );
  NAND2_X1 U488 ( .A1(n610), .A2(n452), .ZN(n408) );
  XOR2_X1 U489 ( .A(KEYINPUT70), .B(G469), .Z(n407) );
  XNOR2_X2 U490 ( .A(G146), .B(G125), .ZN(n469) );
  XOR2_X1 U491 ( .A(KEYINPUT10), .B(n469), .Z(n731) );
  NAND2_X1 U492 ( .A1(G234), .A2(n738), .ZN(n412) );
  XOR2_X1 U493 ( .A(KEYINPUT8), .B(n412), .Z(n447) );
  NAND2_X1 U494 ( .A1(n447), .A2(G221), .ZN(n416) );
  XOR2_X1 U495 ( .A(KEYINPUT24), .B(KEYINPUT94), .Z(n414) );
  XNOR2_X1 U496 ( .A(G119), .B(KEYINPUT23), .ZN(n413) );
  XNOR2_X1 U497 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U498 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U499 ( .A(n418), .B(n417), .ZN(n626) );
  NAND2_X1 U500 ( .A1(n626), .A2(n452), .ZN(n421) );
  NAND2_X1 U501 ( .A1(n605), .A2(G234), .ZN(n419) );
  XNOR2_X1 U502 ( .A(n419), .B(KEYINPUT20), .ZN(n422) );
  XNOR2_X1 U503 ( .A(KEYINPUT25), .B(n377), .ZN(n420) );
  XNOR2_X2 U504 ( .A(n421), .B(n420), .ZN(n571) );
  AND2_X1 U505 ( .A1(n422), .A2(G221), .ZN(n423) );
  XNOR2_X1 U506 ( .A(n423), .B(KEYINPUT21), .ZN(n688) );
  NAND2_X1 U507 ( .A1(n571), .A2(n688), .ZN(n692) );
  NOR2_X1 U508 ( .A1(n504), .A2(n692), .ZN(n596) );
  NAND2_X1 U509 ( .A1(n424), .A2(n596), .ZN(n425) );
  XOR2_X1 U510 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n427) );
  XNOR2_X1 U511 ( .A(G113), .B(KEYINPUT96), .ZN(n426) );
  XNOR2_X1 U512 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U513 ( .A(n429), .B(n428), .Z(n436) );
  XOR2_X1 U514 ( .A(G140), .B(G104), .Z(n431) );
  XNOR2_X1 U515 ( .A(G143), .B(G122), .ZN(n430) );
  XNOR2_X1 U516 ( .A(n431), .B(n430), .ZN(n434) );
  AND2_X1 U517 ( .A1(G214), .A2(n432), .ZN(n433) );
  XNOR2_X1 U518 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U519 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U520 ( .A(n437), .B(n731), .ZN(n632) );
  NAND2_X1 U521 ( .A1(n632), .A2(n452), .ZN(n441) );
  XOR2_X1 U522 ( .A(KEYINPUT98), .B(KEYINPUT13), .Z(n439) );
  XNOR2_X1 U523 ( .A(KEYINPUT97), .B(G475), .ZN(n438) );
  XNOR2_X1 U524 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U525 ( .A(n441), .B(n440), .ZN(n515) );
  XOR2_X1 U526 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n443) );
  XNOR2_X1 U527 ( .A(G116), .B(KEYINPUT7), .ZN(n442) );
  XNOR2_X1 U528 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U529 ( .A(n444), .B(KEYINPUT99), .Z(n446) );
  XNOR2_X1 U530 ( .A(n446), .B(n445), .ZN(n451) );
  NAND2_X1 U531 ( .A1(n447), .A2(G217), .ZN(n449) );
  XNOR2_X1 U532 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U533 ( .A(n451), .B(n450), .ZN(n629) );
  NAND2_X1 U534 ( .A1(n629), .A2(n452), .ZN(n454) );
  INV_X1 U535 ( .A(G478), .ZN(n453) );
  XNOR2_X1 U536 ( .A(n454), .B(n453), .ZN(n513) );
  OR2_X1 U537 ( .A1(n515), .A2(n513), .ZN(n557) );
  INV_X1 U538 ( .A(n455), .ZN(n457) );
  XNOR2_X1 U539 ( .A(KEYINPUT16), .B(G122), .ZN(n456) );
  XNOR2_X2 U540 ( .A(n457), .B(n456), .ZN(n459) );
  XNOR2_X2 U541 ( .A(n459), .B(n458), .ZN(n724) );
  INV_X1 U542 ( .A(n460), .ZN(n461) );
  XNOR2_X1 U543 ( .A(n462), .B(n461), .ZN(n466) );
  XNOR2_X1 U544 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U545 ( .A(n466), .B(n465), .ZN(n471) );
  NAND2_X1 U546 ( .A1(G224), .A2(n738), .ZN(n467) );
  XNOR2_X1 U547 ( .A(n467), .B(KEYINPUT18), .ZN(n468) );
  XNOR2_X1 U548 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U549 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U550 ( .A1(n638), .A2(n605), .ZN(n476) );
  NAND2_X1 U551 ( .A1(n473), .A2(G210), .ZN(n474) );
  XNOR2_X2 U552 ( .A(n476), .B(n475), .ZN(n487) );
  BUF_X2 U553 ( .A(n487), .Z(n538) );
  NOR2_X1 U554 ( .A1(n557), .A2(n538), .ZN(n477) );
  NAND2_X1 U555 ( .A1(n493), .A2(n477), .ZN(n614) );
  INV_X1 U556 ( .A(n614), .ZN(n480) );
  INV_X1 U557 ( .A(KEYINPUT83), .ZN(n478) );
  NOR2_X1 U558 ( .A1(KEYINPUT47), .A2(n478), .ZN(n479) );
  NOR2_X1 U559 ( .A1(n480), .A2(n479), .ZN(n492) );
  INV_X1 U560 ( .A(n688), .ZN(n482) );
  NOR2_X1 U561 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U562 ( .A(n483), .B(KEYINPUT69), .ZN(n484) );
  NOR2_X1 U563 ( .A1(n571), .A2(n484), .ZN(n502) );
  INV_X1 U564 ( .A(n515), .ZN(n485) );
  NAND2_X1 U565 ( .A1(n485), .A2(n513), .ZN(n661) );
  INV_X1 U566 ( .A(n661), .ZN(n658) );
  NAND2_X1 U567 ( .A1(n502), .A2(n658), .ZN(n486) );
  XNOR2_X1 U568 ( .A(n501), .B(KEYINPUT6), .ZN(n586) );
  OR2_X1 U569 ( .A1(n486), .A2(n586), .ZN(n532) );
  INV_X1 U570 ( .A(n487), .ZN(n488) );
  INV_X1 U571 ( .A(n533), .ZN(n677) );
  NOR2_X1 U572 ( .A1(n532), .A2(n517), .ZN(n489) );
  XOR2_X1 U573 ( .A(KEYINPUT36), .B(n489), .Z(n490) );
  XNOR2_X1 U574 ( .A(KEYINPUT111), .B(n490), .ZN(n491) );
  XNOR2_X2 U575 ( .A(n504), .B(KEYINPUT1), .ZN(n691) );
  INV_X1 U576 ( .A(n691), .ZN(n536) );
  NAND2_X1 U577 ( .A1(n491), .A2(n536), .ZN(n667) );
  NAND2_X1 U578 ( .A1(n492), .A2(n667), .ZN(n512) );
  XOR2_X1 U579 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n496) );
  XNOR2_X2 U580 ( .A(n538), .B(KEYINPUT38), .ZN(n497) );
  NAND2_X1 U581 ( .A1(n493), .A2(n497), .ZN(n494) );
  NAND2_X1 U582 ( .A1(n531), .A2(n658), .ZN(n495) );
  XNOR2_X1 U583 ( .A(n496), .B(n495), .ZN(n742) );
  NAND2_X1 U584 ( .A1(n497), .A2(n533), .ZN(n498) );
  AND2_X1 U585 ( .A1(n515), .A2(n513), .ZN(n679) );
  NAND2_X1 U586 ( .A1(n682), .A2(n679), .ZN(n500) );
  XOR2_X1 U587 ( .A(KEYINPUT110), .B(KEYINPUT41), .Z(n499) );
  INV_X1 U588 ( .A(n501), .ZN(n599) );
  INV_X1 U589 ( .A(n599), .ZN(n695) );
  AND2_X1 U590 ( .A1(n695), .A2(n502), .ZN(n503) );
  XOR2_X1 U591 ( .A(n503), .B(KEYINPUT28), .Z(n505) );
  NOR2_X1 U592 ( .A1(n505), .A2(n504), .ZN(n518) );
  INV_X1 U593 ( .A(n518), .ZN(n506) );
  XNOR2_X1 U594 ( .A(n507), .B(KEYINPUT42), .ZN(n745) );
  INV_X1 U595 ( .A(n745), .ZN(n508) );
  NAND2_X1 U596 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U597 ( .A(n510), .B(KEYINPUT46), .ZN(n511) );
  NOR2_X1 U598 ( .A1(n512), .A2(n511), .ZN(n529) );
  INV_X1 U599 ( .A(n513), .ZN(n514) );
  NAND2_X1 U600 ( .A1(n515), .A2(n514), .ZN(n664) );
  INV_X1 U601 ( .A(n664), .ZN(n654) );
  NOR2_X1 U602 ( .A1(n654), .A2(n658), .ZN(n516) );
  XNOR2_X1 U603 ( .A(KEYINPUT101), .B(n516), .ZN(n681) );
  XNOR2_X2 U604 ( .A(n517), .B(KEYINPUT19), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n518), .A2(n552), .ZN(n519) );
  XNOR2_X1 U606 ( .A(n519), .B(KEYINPUT80), .ZN(n527) );
  NOR2_X1 U607 ( .A1(n527), .A2(KEYINPUT66), .ZN(n521) );
  INV_X1 U608 ( .A(n527), .ZN(n657) );
  NOR2_X1 U609 ( .A1(KEYINPUT83), .A2(n657), .ZN(n520) );
  NOR2_X1 U610 ( .A1(n521), .A2(n520), .ZN(n522) );
  NAND2_X1 U611 ( .A1(n681), .A2(n522), .ZN(n523) );
  NAND2_X1 U612 ( .A1(n523), .A2(KEYINPUT47), .ZN(n528) );
  NAND2_X1 U613 ( .A1(n681), .A2(KEYINPUT66), .ZN(n524) );
  NOR2_X1 U614 ( .A1(KEYINPUT47), .A2(n524), .ZN(n525) );
  NOR2_X1 U615 ( .A1(KEYINPUT83), .A2(n525), .ZN(n526) );
  XNOR2_X1 U616 ( .A(n530), .B(KEYINPUT48), .ZN(n543) );
  NAND2_X1 U617 ( .A1(n531), .A2(n654), .ZN(n668) );
  INV_X1 U618 ( .A(n668), .ZN(n541) );
  INV_X1 U619 ( .A(n532), .ZN(n534) );
  NAND2_X1 U620 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U621 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U622 ( .A(n537), .B(KEYINPUT43), .ZN(n540) );
  INV_X1 U623 ( .A(n538), .ZN(n539) );
  NOR2_X1 U624 ( .A1(n540), .A2(n539), .ZN(n615) );
  NOR2_X1 U625 ( .A1(n541), .A2(n615), .ZN(n542) );
  OR2_X1 U626 ( .A1(n586), .A2(n692), .ZN(n544) );
  NOR2_X1 U627 ( .A1(n544), .A2(n691), .ZN(n546) );
  XNOR2_X1 U628 ( .A(KEYINPUT106), .B(KEYINPUT33), .ZN(n545) );
  XNOR2_X1 U629 ( .A(n546), .B(n545), .ZN(n710) );
  INV_X1 U630 ( .A(n710), .ZN(n554) );
  NOR2_X1 U631 ( .A1(G898), .A2(n738), .ZN(n547) );
  XNOR2_X1 U632 ( .A(KEYINPUT92), .B(n547), .ZN(n725) );
  NAND2_X1 U633 ( .A1(n725), .A2(G902), .ZN(n549) );
  NAND2_X1 U634 ( .A1(n549), .A2(n548), .ZN(n550) );
  AND2_X1 U635 ( .A1(n550), .A2(n676), .ZN(n551) );
  NAND2_X1 U636 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X2 U637 ( .A(n553), .B(KEYINPUT0), .ZN(n594) );
  XNOR2_X1 U638 ( .A(n594), .B(KEYINPUT93), .ZN(n597) );
  NAND2_X1 U639 ( .A1(n554), .A2(n597), .ZN(n556) );
  XNOR2_X1 U640 ( .A(KEYINPUT77), .B(KEYINPUT34), .ZN(n555) );
  XNOR2_X1 U641 ( .A(n556), .B(n555), .ZN(n559) );
  INV_X1 U642 ( .A(n557), .ZN(n558) );
  NAND2_X1 U643 ( .A1(n559), .A2(n558), .ZN(n561) );
  XNOR2_X1 U644 ( .A(KEYINPUT76), .B(KEYINPUT35), .ZN(n560) );
  XNOR2_X2 U645 ( .A(n561), .B(n560), .ZN(n619) );
  NAND2_X1 U646 ( .A1(n619), .A2(KEYINPUT86), .ZN(n576) );
  XNOR2_X1 U647 ( .A(n571), .B(KEYINPUT102), .ZN(n689) );
  NOR2_X1 U648 ( .A1(n691), .A2(n689), .ZN(n562) );
  XOR2_X1 U649 ( .A(KEYINPUT105), .B(n562), .Z(n564) );
  XOR2_X1 U650 ( .A(KEYINPUT79), .B(n586), .Z(n563) );
  NAND2_X1 U651 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U652 ( .A1(n679), .A2(n688), .ZN(n565) );
  NOR2_X1 U653 ( .A1(n566), .A2(n588), .ZN(n568) );
  XOR2_X1 U654 ( .A(KEYINPUT78), .B(KEYINPUT32), .Z(n567) );
  XNOR2_X1 U655 ( .A(n568), .B(n567), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n580), .A2(KEYINPUT44), .ZN(n574) );
  NAND2_X1 U657 ( .A1(n691), .A2(n599), .ZN(n569) );
  INV_X1 U658 ( .A(KEYINPUT64), .ZN(n570) );
  INV_X1 U659 ( .A(n571), .ZN(n572) );
  NOR2_X1 U660 ( .A1(n574), .A2(n581), .ZN(n575) );
  NAND2_X1 U661 ( .A1(n576), .A2(n575), .ZN(n579) );
  INV_X1 U662 ( .A(KEYINPUT44), .ZN(n577) );
  NAND2_X1 U663 ( .A1(n577), .A2(KEYINPUT86), .ZN(n578) );
  INV_X1 U664 ( .A(n580), .ZN(n616) );
  NAND2_X1 U665 ( .A1(n582), .A2(n617), .ZN(n583) );
  NAND2_X1 U666 ( .A1(n583), .A2(KEYINPUT86), .ZN(n585) );
  INV_X1 U667 ( .A(n619), .ZN(n584) );
  INV_X1 U668 ( .A(n586), .ZN(n587) );
  XNOR2_X1 U669 ( .A(n589), .B(KEYINPUT85), .ZN(n591) );
  NAND2_X1 U670 ( .A1(n691), .A2(n689), .ZN(n590) );
  NOR2_X1 U671 ( .A1(n691), .A2(n692), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n593), .A2(n695), .ZN(n700) );
  NOR2_X1 U673 ( .A1(n700), .A2(n594), .ZN(n595) );
  XNOR2_X1 U674 ( .A(n595), .B(KEYINPUT31), .ZN(n663) );
  NAND2_X1 U675 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U676 ( .A(n598), .B(KEYINPUT95), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n650) );
  NAND2_X1 U678 ( .A1(n663), .A2(n650), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n601), .A2(n681), .ZN(n602) );
  NOR2_X1 U680 ( .A1(n669), .A2(n374), .ZN(n604) );
  INV_X1 U681 ( .A(KEYINPUT2), .ZN(n606) );
  INV_X1 U682 ( .A(n673), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n637), .A2(G469), .ZN(n611) );
  XNOR2_X1 U684 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n611), .B(n358), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n612), .A2(n644), .ZN(n613) );
  XNOR2_X1 U687 ( .A(n613), .B(KEYINPUT121), .ZN(G54) );
  XNOR2_X1 U688 ( .A(n614), .B(G143), .ZN(G45) );
  XOR2_X1 U689 ( .A(G140), .B(n615), .Z(G42) );
  XNOR2_X1 U690 ( .A(n580), .B(G119), .ZN(G21) );
  XNOR2_X1 U691 ( .A(n617), .B(G110), .ZN(G12) );
  XNOR2_X1 U692 ( .A(n618), .B(G101), .ZN(G3) );
  XOR2_X1 U693 ( .A(n619), .B(G122), .Z(G24) );
  NAND2_X1 U694 ( .A1(n637), .A2(G472), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n621), .B(n360), .ZN(n622) );
  XOR2_X1 U696 ( .A(KEYINPUT112), .B(KEYINPUT63), .Z(n623) );
  XNOR2_X1 U697 ( .A(n624), .B(n623), .ZN(G57) );
  NAND2_X1 U698 ( .A1(n637), .A2(G217), .ZN(n625) );
  XOR2_X1 U699 ( .A(n626), .B(n625), .Z(n627) );
  NOR2_X1 U700 ( .A1(n627), .A2(n643), .ZN(G66) );
  NAND2_X1 U701 ( .A1(n637), .A2(G478), .ZN(n628) );
  XOR2_X1 U702 ( .A(n629), .B(n628), .Z(n630) );
  NOR2_X1 U703 ( .A1(n630), .A2(n643), .ZN(G63) );
  NAND2_X1 U704 ( .A1(n637), .A2(G475), .ZN(n633) );
  XOR2_X1 U705 ( .A(KEYINPUT65), .B(KEYINPUT59), .Z(n631) );
  XNOR2_X1 U706 ( .A(n633), .B(n359), .ZN(n634) );
  XNOR2_X1 U707 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(G60) );
  NAND2_X1 U709 ( .A1(n637), .A2(G210), .ZN(n642) );
  BUF_X1 U710 ( .A(n638), .Z(n639) );
  XNOR2_X1 U711 ( .A(KEYINPUT87), .B(KEYINPUT54), .ZN(n640) );
  XOR2_X1 U712 ( .A(n640), .B(KEYINPUT55), .Z(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n361), .ZN(n645) );
  INV_X1 U714 ( .A(n643), .ZN(n644) );
  XNOR2_X1 U715 ( .A(n646), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X1 U716 ( .A1(n661), .A2(n650), .ZN(n648) );
  XNOR2_X1 U717 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U719 ( .A(G104), .B(n649), .ZN(G6) );
  NOR2_X1 U720 ( .A1(n664), .A2(n650), .ZN(n652) );
  XNOR2_X1 U721 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U723 ( .A(G107), .B(n653), .ZN(G9) );
  XOR2_X1 U724 ( .A(G128), .B(KEYINPUT29), .Z(n656) );
  NAND2_X1 U725 ( .A1(n654), .A2(n657), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n656), .B(n655), .ZN(G30) );
  XOR2_X1 U727 ( .A(G146), .B(KEYINPUT115), .Z(n660) );
  NAND2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n660), .B(n659), .ZN(G48) );
  NOR2_X1 U730 ( .A1(n661), .A2(n663), .ZN(n662) );
  XOR2_X1 U731 ( .A(G113), .B(n662), .Z(G15) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U733 ( .A(G116), .B(n665), .Z(G18) );
  XOR2_X1 U734 ( .A(G125), .B(KEYINPUT37), .Z(n666) );
  XNOR2_X1 U735 ( .A(n667), .B(n666), .ZN(G27) );
  XNOR2_X1 U736 ( .A(G134), .B(n668), .ZN(G36) );
  XOR2_X1 U737 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n717) );
  BUF_X1 U738 ( .A(n669), .Z(n671) );
  XOR2_X1 U739 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n670) );
  NAND2_X1 U740 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U741 ( .A(n672), .B(KEYINPUT81), .ZN(n674) );
  NOR2_X1 U742 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U743 ( .A1(n675), .A2(G953), .ZN(n715) );
  INV_X1 U744 ( .A(n676), .ZN(n707) );
  INV_X1 U745 ( .A(n497), .ZN(n678) );
  NAND2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n680) );
  NAND2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n684) );
  NAND2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U750 ( .A(KEYINPUT117), .B(n685), .ZN(n686) );
  NOR2_X1 U751 ( .A1(n710), .A2(n686), .ZN(n687) );
  XNOR2_X1 U752 ( .A(n687), .B(KEYINPUT118), .ZN(n704) );
  NOR2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U754 ( .A(KEYINPUT49), .B(n690), .ZN(n698) );
  XOR2_X1 U755 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n694) );
  NAND2_X1 U756 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U757 ( .A(n694), .B(n693), .ZN(n696) );
  NOR2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U759 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U760 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U761 ( .A(KEYINPUT51), .B(n701), .ZN(n702) );
  NOR2_X1 U762 ( .A1(n702), .A2(n711), .ZN(n703) );
  NOR2_X1 U763 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U764 ( .A(n705), .B(KEYINPUT52), .ZN(n706) );
  NOR2_X1 U765 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U766 ( .A1(n708), .A2(G952), .ZN(n709) );
  XNOR2_X1 U767 ( .A(n709), .B(KEYINPUT119), .ZN(n713) );
  NOR2_X1 U768 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U769 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U770 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U771 ( .A(n717), .B(n716), .ZN(G75) );
  NAND2_X1 U772 ( .A1(n718), .A2(n738), .ZN(n723) );
  NAND2_X1 U773 ( .A1(G953), .A2(G224), .ZN(n719) );
  XNOR2_X1 U774 ( .A(KEYINPUT61), .B(n719), .ZN(n720) );
  NAND2_X1 U775 ( .A1(n720), .A2(G898), .ZN(n721) );
  XOR2_X1 U776 ( .A(KEYINPUT123), .B(n721), .Z(n722) );
  NAND2_X1 U777 ( .A1(n723), .A2(n722), .ZN(n728) );
  XOR2_X1 U778 ( .A(n724), .B(G101), .Z(n726) );
  NOR2_X1 U779 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U780 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U781 ( .A(KEYINPUT124), .B(n729), .ZN(G69) );
  XNOR2_X1 U782 ( .A(KEYINPUT4), .B(n730), .ZN(n732) );
  XOR2_X1 U783 ( .A(n732), .B(n731), .Z(n737) );
  XNOR2_X1 U784 ( .A(n737), .B(KEYINPUT125), .ZN(n733) );
  XNOR2_X1 U785 ( .A(G227), .B(n733), .ZN(n734) );
  NAND2_X1 U786 ( .A1(G900), .A2(n734), .ZN(n735) );
  NAND2_X1 U787 ( .A1(n735), .A2(G953), .ZN(n741) );
  XNOR2_X1 U788 ( .A(n737), .B(n736), .ZN(n739) );
  NAND2_X1 U789 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U790 ( .A1(n741), .A2(n740), .ZN(G72) );
  XNOR2_X1 U791 ( .A(n742), .B(G131), .ZN(n743) );
  XNOR2_X1 U792 ( .A(n743), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U793 ( .A(G137), .B(KEYINPUT126), .Z(n744) );
  XNOR2_X1 U794 ( .A(n745), .B(n744), .ZN(G39) );
endmodule

