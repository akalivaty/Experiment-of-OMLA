//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT75), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT22), .ZN(new_n205));
  INV_X1    g004(.A(G211gat), .ZN(new_n206));
  INV_X1    g005(.A(G218gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT71), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n204), .A3(new_n208), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n209), .A2(KEYINPUT71), .A3(new_n211), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT73), .ZN(new_n219));
  XOR2_X1   g018(.A(KEYINPUT27), .B(G183gat), .Z(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G190gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT67), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n222), .A2(new_n223), .B1(G183gat), .B2(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226));
  INV_X1    g025(.A(G169gat), .ZN(new_n227));
  INV_X1    g026(.A(G176gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n226), .B1(new_n229), .B2(KEYINPUT26), .ZN(new_n230));
  NOR2_X1   g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n231), .A2(KEYINPUT68), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n231), .B(KEYINPUT64), .ZN(new_n234));
  OAI221_X1 g033(.A(new_n225), .B1(new_n230), .B2(new_n233), .C1(new_n234), .C2(KEYINPUT26), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n224), .B(new_n235), .C1(new_n223), .C2(new_n222), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(new_n221), .B2(G183gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n225), .A2(KEYINPUT23), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(new_n229), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT23), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT25), .B(new_n245), .C1(new_n234), .C2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n229), .ZN(new_n248));
  OR2_X1    g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n238), .A2(new_n240), .A3(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  OAI22_X1  g050(.A1(new_n243), .A2(new_n247), .B1(new_n251), .B2(KEYINPUT25), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT29), .B1(new_n236), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G226gat), .ZN(new_n254));
  INV_X1    g053(.A(G233gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n219), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n256), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(new_n236), .B2(new_n252), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n236), .A2(new_n252), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT29), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n259), .B1(new_n262), .B2(new_n258), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n218), .B(new_n257), .C1(new_n263), .C2(new_n219), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n217), .A2(KEYINPUT72), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n217), .A2(KEYINPUT72), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n253), .A2(new_n256), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n267), .B1(new_n268), .B2(new_n259), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G8gat), .B(G36gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(G64gat), .B(G92gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n264), .A2(new_n269), .A3(new_n273), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(KEYINPUT30), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT30), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n264), .A2(new_n278), .A3(new_n269), .A4(new_n273), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT2), .ZN(new_n281));
  INV_X1    g080(.A(G148gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(G141gat), .ZN(new_n283));
  INV_X1    g082(.A(G141gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(G148gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n281), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287));
  INV_X1    g086(.A(G155gat), .ZN(new_n288));
  INV_X1    g087(.A(G162gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n286), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT74), .B1(new_n282), .B2(G141gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT74), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(new_n284), .A3(G148gat), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n292), .B(new_n294), .C1(new_n284), .C2(G148gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n287), .B1(new_n290), .B2(KEYINPUT2), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT3), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G113gat), .B(G120gat), .Z(new_n301));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G127gat), .B(G134gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(new_n302), .A3(new_n304), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n297), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT3), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n300), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n306), .A2(new_n307), .A3(new_n291), .A4(new_n297), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT4), .ZN(new_n314));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT4), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n311), .A2(new_n314), .A3(new_n315), .A4(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n315), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n307), .A2(new_n306), .B1(new_n291), .B2(new_n297), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n319), .B1(new_n313), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT5), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G1gat), .B(G29gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT0), .ZN(new_n325));
  XNOR2_X1  g124(.A(G57gat), .B(G85gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT4), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n328), .A2(KEYINPUT5), .A3(new_n315), .A4(new_n311), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n323), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT6), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n323), .A2(new_n329), .ZN(new_n333));
  INV_X1    g132(.A(new_n327), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT6), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n332), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n203), .B1(new_n280), .B2(new_n337), .ZN(new_n338));
  AOI211_X1 g137(.A(KEYINPUT75), .B(new_n336), .C1(new_n277), .C2(new_n279), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n300), .A2(new_n261), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n265), .A2(new_n341), .A3(new_n266), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n299), .B1(new_n217), .B2(KEYINPUT29), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n309), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n342), .A2(G228gat), .A3(G233gat), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G228gat), .A2(G233gat), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n218), .B1(new_n261), .B2(new_n300), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n212), .A2(new_n214), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(new_n261), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n298), .B1(new_n349), .B2(new_n299), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n346), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G22gat), .ZN(new_n353));
  INV_X1    g152(.A(G22gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n345), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G78gat), .B(G106gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT31), .B(G50gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n354), .B1(new_n345), .B2(new_n351), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n359), .B1(new_n360), .B2(KEYINPUT76), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n353), .A2(KEYINPUT76), .A3(new_n355), .A4(new_n359), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(KEYINPUT69), .B(G71gat), .Z(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(G99gat), .ZN(new_n366));
  XOR2_X1   g165(.A(G15gat), .B(G43gat), .Z(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G227gat), .A2(G233gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n260), .A2(new_n308), .ZN(new_n371));
  INV_X1    g170(.A(new_n308), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n236), .A2(new_n252), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n370), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n369), .B1(new_n374), .B2(KEYINPUT33), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n371), .A2(new_n370), .A3(new_n373), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT34), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n236), .A2(new_n252), .A3(new_n372), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n372), .B1(new_n236), .B2(new_n252), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT34), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(new_n370), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n375), .A2(new_n377), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n370), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(new_n378), .B2(new_n379), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT33), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n368), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n381), .B1(new_n380), .B2(new_n370), .ZN(new_n388));
  NOR4_X1   g187(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT34), .A4(new_n384), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n383), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n385), .A2(KEYINPUT32), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n392), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n383), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n364), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n383), .A2(new_n390), .A3(new_n394), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n394), .B1(new_n383), .B2(new_n390), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(KEYINPUT81), .A3(new_n364), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n202), .B1(new_n340), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n327), .B(KEYINPUT78), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT79), .B1(new_n333), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n405), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n323), .A2(new_n407), .A3(new_n408), .A4(new_n329), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n335), .ZN(new_n411));
  INV_X1    g210(.A(new_n332), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT35), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n280), .A2(new_n401), .A3(new_n413), .A4(new_n364), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT80), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n364), .A2(new_n393), .A3(new_n395), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT80), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n416), .A2(new_n417), .A3(new_n280), .A4(new_n413), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n364), .B(KEYINPUT77), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n280), .A2(new_n337), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT75), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n280), .A2(new_n203), .A3(new_n337), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n425));
  AND2_X1   g224(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n393), .B(new_n395), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n401), .B2(new_n426), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n328), .A2(new_n311), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n319), .ZN(new_n430));
  OR2_X1    g229(.A1(new_n313), .A2(new_n320), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n430), .B(KEYINPUT39), .C1(new_n319), .C2(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n432), .B(new_n405), .C1(KEYINPUT39), .C2(new_n430), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT40), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n410), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n364), .B1(new_n435), .B2(new_n280), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n411), .A2(new_n412), .A3(new_n276), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT38), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n270), .B2(KEYINPUT37), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n439), .B(new_n274), .C1(KEYINPUT37), .C2(new_n270), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n274), .B1(new_n270), .B2(KEYINPUT37), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT37), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n257), .B1(new_n263), .B2(new_n219), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n217), .ZN(new_n444));
  OR3_X1    g243(.A1(new_n268), .A2(new_n267), .A3(new_n259), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n438), .B1(new_n441), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n437), .B1(new_n440), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n428), .B1(new_n436), .B2(new_n448), .ZN(new_n449));
  OAI22_X1  g248(.A1(new_n404), .A2(new_n419), .B1(new_n424), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT88), .ZN(new_n451));
  NAND2_X1  g250(.A1(G229gat), .A2(G233gat), .ZN(new_n452));
  INV_X1    g251(.A(G50gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G43gat), .ZN(new_n454));
  INV_X1    g253(.A(G43gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G50gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n456), .A3(KEYINPUT15), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT82), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT82), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n460), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT14), .ZN(new_n462));
  INV_X1    g261(.A(G29gat), .ZN(new_n463));
  INV_X1    g262(.A(G36gat), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n459), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  AND3_X1   g265(.A1(KEYINPUT83), .A2(G29gat), .A3(G36gat), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT83), .B1(G29gat), .B2(G36gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n457), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n465), .A2(new_n458), .ZN(new_n472));
  XNOR2_X1  g271(.A(G43gat), .B(G50gat), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n472), .B1(KEYINPUT15), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n469), .A2(new_n457), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n454), .A2(new_n456), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT15), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n477), .A2(new_n478), .B1(new_n458), .B2(new_n465), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n479), .A2(KEYINPUT84), .A3(new_n457), .A4(new_n469), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n470), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT16), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(G1gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n487));
  INV_X1    g286(.A(G8gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n482), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n482), .B2(new_n487), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n486), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n482), .A2(new_n487), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G8gat), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n494), .A2(new_n485), .A3(new_n484), .A4(new_n489), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n452), .B1(new_n481), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n470), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n474), .A2(new_n475), .A3(new_n471), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n469), .A2(new_n457), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT84), .B1(new_n500), .B2(new_n479), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n498), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT86), .ZN(new_n503));
  XOR2_X1   g302(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT86), .B1(new_n481), .B2(new_n504), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n492), .A2(new_n495), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(KEYINPUT17), .B2(new_n481), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n497), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n451), .B1(new_n511), .B2(KEYINPUT18), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n452), .B(KEYINPUT13), .Z(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n502), .A2(new_n509), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n481), .A2(new_n496), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n511), .B2(KEYINPUT18), .ZN(new_n518));
  XNOR2_X1  g317(.A(G113gat), .B(G141gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(G197gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT11), .B(G169gat), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n520), .B(new_n521), .Z(new_n522));
  XOR2_X1   g321(.A(new_n522), .B(KEYINPUT12), .Z(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT18), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT17), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n496), .B1(new_n502), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n527), .B1(new_n507), .B2(new_n506), .ZN(new_n528));
  OAI211_X1 g327(.A(KEYINPUT88), .B(new_n525), .C1(new_n528), .C2(new_n497), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n512), .A2(new_n518), .A3(new_n524), .A4(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n503), .B1(new_n502), .B2(new_n505), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n481), .A2(KEYINPUT86), .A3(new_n504), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n510), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n497), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(KEYINPUT18), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n517), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n511), .A2(KEYINPUT18), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n523), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n530), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n450), .A2(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G64gat), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT90), .B1(new_n548), .B2(G57gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n550));
  INV_X1    g349(.A(G57gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n551), .A3(G64gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n548), .A2(G57gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n547), .B1(KEYINPUT91), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n549), .A2(new_n552), .A3(new_n556), .A4(new_n553), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n551), .A2(G64gat), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n545), .B1(new_n558), .B2(new_n553), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n559), .B1(KEYINPUT89), .B2(new_n544), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n561), .A3(new_n543), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n555), .A2(new_n557), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G127gat), .B(G155gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n509), .B1(KEYINPUT21), .B2(new_n563), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n568), .B(new_n569), .Z(new_n570));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT93), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(new_n576), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(KEYINPUT41), .ZN(new_n581));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n581), .B(new_n582), .Z(new_n583));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n580), .A2(KEYINPUT41), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  INV_X1    g386(.A(G92gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT7), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n590), .B1(new_n587), .B2(new_n588), .ZN(new_n591));
  NAND3_X1  g390(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n589), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G99gat), .B(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT94), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n589), .A2(new_n594), .A3(new_n591), .A4(new_n592), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n593), .A2(KEYINPUT94), .A3(new_n595), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n585), .B1(new_n602), .B2(new_n481), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n481), .B2(KEYINPUT17), .ZN(new_n604));
  AOI211_X1 g403(.A(new_n584), .B(new_n603), .C1(new_n508), .C2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n584), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n604), .B1(new_n531), .B2(new_n532), .ZN(new_n607));
  INV_X1    g406(.A(new_n603), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n583), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g411(.A(KEYINPUT95), .B(new_n583), .C1(new_n605), .C2(new_n609), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(KEYINPUT96), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT96), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n603), .B1(new_n508), .B2(new_n604), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n615), .B1(new_n616), .B2(new_n606), .ZN(new_n617));
  INV_X1    g416(.A(new_n583), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n607), .A2(new_n606), .A3(new_n608), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n614), .A2(new_n617), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n612), .A2(new_n613), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n602), .A2(new_n564), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n554), .A2(KEYINPUT91), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n625), .A2(new_n557), .A3(new_n544), .A4(new_n546), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n544), .A2(KEYINPUT89), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n558), .A2(new_n553), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n627), .B(new_n562), .C1(new_n545), .C2(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n626), .A2(new_n629), .A3(new_n596), .A4(new_n598), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n623), .B1(new_n624), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n630), .B(new_n633), .C1(new_n601), .C2(new_n563), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n626), .A2(KEYINPUT10), .A3(new_n629), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n601), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n623), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  NAND3_X1  g440(.A1(new_n632), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n634), .A2(new_n636), .B1(G230gat), .B2(G233gat), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n631), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n579), .A2(new_n622), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n541), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n337), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT97), .B(G1gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1324gat));
  INV_X1    g452(.A(new_n280), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n541), .A2(new_n654), .A3(new_n649), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT16), .B(G8gat), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n658), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n655), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(KEYINPUT42), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT98), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n661), .B(new_n663), .C1(new_n655), .C2(new_n657), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n659), .B1(new_n662), .B2(new_n665), .ZN(G1325gat));
  INV_X1    g465(.A(new_n650), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n401), .ZN(new_n668));
  INV_X1    g467(.A(G15gat), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT99), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n668), .A2(new_n672), .A3(new_n669), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n428), .A2(new_n669), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT100), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n671), .A2(new_n673), .B1(new_n667), .B2(new_n675), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n650), .A2(new_n420), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  INV_X1    g478(.A(KEYINPUT45), .ZN(new_n680));
  INV_X1    g479(.A(new_n579), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n647), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n622), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n541), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n337), .A2(G29gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n685), .B1(new_n684), .B2(new_n686), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n680), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n689), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(KEYINPUT45), .A3(new_n687), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n403), .A2(new_n422), .A3(new_n423), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n419), .B1(KEYINPUT35), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n449), .A2(new_n424), .ZN(new_n695));
  OAI211_X1 g494(.A(KEYINPUT103), .B(new_n621), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n450), .A2(KEYINPUT103), .A3(KEYINPUT44), .A4(new_n621), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n540), .A2(KEYINPUT102), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n530), .B2(new_n539), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n682), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n698), .A2(new_n699), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(G29gat), .B1(new_n705), .B2(new_n337), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n692), .A3(new_n706), .ZN(G1328gat));
  OAI21_X1  g506(.A(G36gat), .B1(new_n705), .B2(new_n280), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n280), .A2(G36gat), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n450), .A2(new_n540), .A3(new_n683), .A4(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT46), .Z(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT104), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n708), .A2(new_n714), .A3(new_n711), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(G1329gat));
  NAND2_X1  g515(.A1(new_n541), .A2(new_n683), .ZN(new_n717));
  INV_X1    g516(.A(new_n401), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n455), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n428), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G43gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n705), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g522(.A(G50gat), .B1(new_n705), .B2(new_n364), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n420), .A2(G50gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n684), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n724), .A2(KEYINPUT48), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n420), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n698), .A2(new_n728), .A3(new_n699), .A4(new_n704), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n729), .A2(G50gat), .B1(new_n684), .B2(new_n725), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n727), .B1(new_n730), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g530(.A(new_n703), .ZN(new_n732));
  NOR4_X1   g531(.A1(new_n732), .A2(new_n681), .A3(new_n621), .A4(new_n647), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n450), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n337), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(new_n551), .ZN(G1332gat));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n734), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n654), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n740));
  XOR2_X1   g539(.A(KEYINPUT49), .B(G64gat), .Z(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n739), .B2(new_n741), .ZN(G1333gat));
  NAND3_X1  g541(.A1(new_n738), .A2(G71gat), .A3(new_n720), .ZN(new_n743));
  INV_X1    g542(.A(G71gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n734), .B2(new_n718), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n743), .A2(new_n745), .A3(new_n747), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(G1334gat));
  NAND2_X1  g550(.A1(new_n738), .A2(new_n728), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g552(.A1(new_n703), .A2(new_n681), .A3(new_n646), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT107), .Z(new_n755));
  NAND3_X1  g554(.A1(new_n698), .A2(new_n699), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G85gat), .B1(new_n756), .B2(new_n337), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n732), .A2(new_n579), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n450), .A2(new_n621), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n450), .A2(KEYINPUT51), .A3(new_n621), .A4(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n336), .A2(new_n587), .A3(new_n646), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n757), .B1(new_n764), .B2(new_n765), .ZN(G1336gat));
  OAI21_X1  g565(.A(G92gat), .B1(new_n756), .B2(new_n280), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n761), .A2(KEYINPUT108), .A3(new_n762), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n759), .A2(new_n769), .A3(new_n760), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n280), .A2(G92gat), .A3(new_n647), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n768), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT52), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(new_n763), .B2(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n767), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(G1337gat));
  NAND4_X1  g576(.A1(new_n698), .A2(new_n720), .A3(new_n699), .A4(new_n755), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT109), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G99gat), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n778), .A2(KEYINPUT109), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n718), .A2(G99gat), .A3(new_n647), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT110), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n780), .A2(new_n781), .B1(new_n764), .B2(new_n783), .ZN(G1338gat));
  NOR3_X1   g583(.A1(new_n364), .A2(G106gat), .A3(new_n647), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT53), .B1(new_n763), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n364), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n698), .A2(new_n787), .A3(new_n699), .A4(new_n755), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT111), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G106gat), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n788), .A2(KEYINPUT111), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n786), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G106gat), .B1(new_n756), .B2(new_n420), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n768), .A2(new_n770), .A3(new_n785), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT53), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n796), .ZN(G1339gat));
  AOI21_X1  g596(.A(new_n623), .B1(new_n635), .B2(new_n601), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n634), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT54), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT55), .B1(new_n800), .B2(new_n644), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n643), .B1(new_n638), .B2(KEYINPUT54), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n642), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n641), .B1(new_n644), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n798), .B2(new_n634), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n638), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT55), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n700), .A2(new_n702), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n515), .A2(new_n516), .A3(new_n514), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n812), .B(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n452), .B1(new_n533), .B2(new_n515), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n522), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n530), .A2(new_n646), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n622), .B1(new_n811), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n522), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n812), .B(KEYINPUT112), .ZN(new_n821));
  INV_X1    g620(.A(new_n452), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n481), .A2(new_n496), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n528), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n820), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n512), .A2(new_n529), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n537), .A2(new_n523), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n621), .A2(new_n828), .A3(new_n809), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n819), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n681), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n732), .A2(new_n648), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n337), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n834), .A2(new_n280), .A3(new_n403), .ZN(new_n835));
  INV_X1    g634(.A(G113gat), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n836), .A3(new_n732), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n728), .B1(new_n831), .B2(new_n833), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n654), .A2(new_n718), .A3(new_n337), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n540), .A3(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n840), .A2(new_n841), .A3(G113gat), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n840), .B2(G113gat), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n837), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT114), .ZN(G1340gat));
  NAND2_X1  g644(.A1(new_n838), .A2(new_n839), .ZN(new_n846));
  INV_X1    g645(.A(G120gat), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n846), .A2(new_n847), .A3(new_n647), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n835), .A2(new_n646), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(new_n847), .ZN(G1341gat));
  INV_X1    g649(.A(G127gat), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n835), .A2(new_n851), .A3(new_n579), .ZN(new_n852));
  OAI21_X1  g651(.A(G127gat), .B1(new_n846), .B2(new_n681), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1342gat));
  NOR2_X1   g653(.A1(new_n622), .A2(G134gat), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n835), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT115), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n835), .A2(new_n858), .A3(new_n855), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n857), .A2(KEYINPUT56), .A3(new_n859), .ZN(new_n863));
  OAI21_X1  g662(.A(G134gat), .B1(new_n846), .B2(new_n622), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(G1343gat));
  NOR2_X1   g664(.A1(new_n720), .A2(new_n364), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n834), .A2(new_n866), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(KEYINPUT118), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(KEYINPUT118), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n868), .A2(new_n280), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n540), .A2(new_n284), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n428), .A2(new_n336), .A3(new_n280), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n828), .A2(new_n646), .B1(new_n540), .B2(new_n809), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n829), .B1(new_n876), .B2(new_n621), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n877), .A2(new_n681), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n728), .B1(new_n878), .B2(new_n832), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n875), .B1(new_n879), .B2(KEYINPUT57), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n579), .B1(new_n819), .B2(new_n829), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n881), .B(new_n787), .C1(new_n882), .C2(new_n832), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n539), .B2(new_n530), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n874), .B1(new_n885), .B2(new_n284), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n834), .A2(new_n280), .A3(new_n866), .A4(new_n872), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n887), .B(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n880), .A2(new_n732), .A3(new_n883), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n890), .A2(KEYINPUT116), .A3(G141gat), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT116), .B1(new_n890), .B2(G141gat), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n889), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n873), .A2(new_n886), .B1(new_n893), .B2(new_n874), .ZN(G1344gat));
  NAND3_X1  g693(.A1(new_n870), .A2(new_n282), .A3(new_n646), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n896), .B(G148gat), .C1(new_n884), .C2(new_n647), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n648), .A2(new_n540), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n579), .B1(new_n877), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(KEYINPUT119), .B(new_n829), .C1(new_n876), .C2(new_n621), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n898), .B(new_n881), .C1(new_n903), .C2(new_n420), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n540), .A2(new_n809), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n621), .B1(new_n905), .B2(new_n817), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n805), .A2(new_n807), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT55), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n644), .A2(new_n631), .A3(new_n643), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n908), .B1(new_n638), .B2(new_n806), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n805), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n530), .A2(new_n816), .A3(new_n909), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n607), .A2(new_n608), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT96), .B1(new_n914), .B2(new_n584), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n619), .A2(new_n618), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI22_X1  g716(.A1(new_n917), .A2(new_n614), .B1(new_n610), .B2(new_n611), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n913), .B1(new_n613), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n900), .B1(new_n906), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n902), .A3(new_n681), .ZN(new_n921));
  INV_X1    g720(.A(new_n899), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n420), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT120), .B1(new_n923), .B2(KEYINPUT57), .ZN(new_n924));
  OAI211_X1 g723(.A(KEYINPUT57), .B(new_n787), .C1(new_n882), .C2(new_n832), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n904), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n875), .A2(new_n647), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n282), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n897), .B1(new_n928), .B2(new_n896), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n895), .A2(new_n929), .ZN(G1345gat));
  NAND3_X1  g729(.A1(new_n870), .A2(new_n288), .A3(new_n579), .ZN(new_n931));
  OAI21_X1  g730(.A(G155gat), .B1(new_n884), .B2(new_n681), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1346gat));
  NAND3_X1  g732(.A1(new_n870), .A2(new_n289), .A3(new_n621), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n880), .A2(new_n621), .A3(new_n883), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n289), .B1(new_n935), .B2(KEYINPUT121), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n936), .B1(KEYINPUT121), .B2(new_n935), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(G1347gat));
  AOI21_X1  g737(.A(new_n336), .B1(new_n831), .B2(new_n833), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n280), .B1(new_n398), .B2(new_n402), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n227), .A3(new_n732), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n654), .A2(new_n337), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(new_n718), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n838), .A2(new_n540), .A3(new_n945), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n946), .A2(KEYINPUT122), .A3(G169gat), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT122), .B1(new_n946), .B2(G169gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n943), .B1(new_n947), .B2(new_n948), .ZN(G1348gat));
  NAND2_X1  g748(.A1(new_n838), .A2(new_n945), .ZN(new_n950));
  OAI21_X1  g749(.A(G176gat), .B1(new_n950), .B2(new_n647), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n646), .A2(new_n228), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n941), .B2(new_n952), .ZN(G1349gat));
  OAI21_X1  g752(.A(G183gat), .B1(new_n950), .B2(new_n681), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT123), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n681), .A2(new_n220), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n954), .B(new_n955), .C1(new_n941), .C2(new_n956), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g757(.A(G190gat), .B1(new_n950), .B2(new_n622), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n959), .A2(KEYINPUT124), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n962), .B1(KEYINPUT124), .B2(new_n959), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n941), .A2(new_n221), .A3(new_n622), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n964), .B1(new_n960), .B2(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1351gat));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n720), .A2(new_n944), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(new_n540), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n926), .A2(KEYINPUT125), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT125), .B1(new_n926), .B2(new_n969), .ZN(new_n971));
  INV_X1    g770(.A(G197gat), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n939), .A2(new_n654), .A3(new_n866), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n974), .A2(new_n972), .A3(new_n732), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n967), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n926), .A2(new_n969), .ZN(new_n978));
  OAI21_X1  g777(.A(G197gat), .B1(new_n978), .B2(KEYINPUT125), .ZN(new_n979));
  OAI211_X1 g778(.A(KEYINPUT126), .B(new_n975), .C1(new_n979), .C2(new_n970), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n977), .A2(new_n980), .ZN(G1352gat));
  XNOR2_X1  g780(.A(KEYINPUT127), .B(G204gat), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n647), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n974), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g783(.A(new_n984), .B(KEYINPUT62), .Z(new_n985));
  NAND2_X1  g784(.A1(new_n926), .A2(new_n968), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n982), .B1(new_n986), .B2(new_n647), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n985), .A2(new_n987), .ZN(G1353gat));
  NAND3_X1  g787(.A1(new_n974), .A2(new_n206), .A3(new_n579), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n926), .A2(new_n579), .A3(new_n968), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n990), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n991));
  AOI21_X1  g790(.A(KEYINPUT63), .B1(new_n990), .B2(G211gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(G1354gat));
  OAI21_X1  g792(.A(G218gat), .B1(new_n986), .B2(new_n622), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n974), .A2(new_n207), .A3(new_n621), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(G1355gat));
endmodule


