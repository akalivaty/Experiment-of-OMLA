//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953;
  INV_X1    g000(.A(KEYINPUT5), .ZN(new_n202));
  OR2_X1    g001(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(G134gat), .A3(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G134gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT67), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT67), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G134gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n209), .A3(G127gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G120gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G113gat), .ZN(new_n213));
  INV_X1    g012(.A(G113gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G120gat), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT1), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G141gat), .B(G148gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n223), .B1(G155gat), .B2(G162gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n221), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G141gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G148gat), .ZN(new_n227));
  INV_X1    g026(.A(G148gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G141gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G155gat), .B(G162gat), .ZN(new_n231));
  INV_X1    g030(.A(G155gat), .ZN(new_n232));
  INV_X1    g031(.A(G162gat), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT2), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G127gat), .B(G134gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n218), .A2(new_n225), .A3(new_n235), .A4(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n225), .A2(new_n235), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n216), .B1(new_n210), .B2(new_n205), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n216), .A2(new_n236), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n202), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n238), .A2(KEYINPUT4), .ZN(new_n247));
  XOR2_X1   g046(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n248));
  NOR2_X1   g047(.A1(new_n240), .A2(new_n241), .ZN(new_n249));
  INV_X1    g048(.A(new_n239), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n239), .A2(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n218), .A2(new_n237), .ZN(new_n254));
  XOR2_X1   g053(.A(KEYINPUT75), .B(KEYINPUT3), .Z(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n253), .B(new_n254), .C1(new_n239), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n244), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n246), .B1(new_n252), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n238), .A2(KEYINPUT4), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n249), .A2(new_n250), .A3(new_n248), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT78), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n225), .A2(new_n235), .A3(new_n255), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT3), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n264), .B1(new_n225), .B2(new_n235), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n245), .B1(new_n266), .B2(new_n254), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT78), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n249), .A2(new_n268), .A3(new_n250), .A4(new_n248), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n262), .A2(new_n267), .A3(new_n202), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n259), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G1gat), .B(G29gat), .Z(new_n272));
  XNOR2_X1  g071(.A(G57gat), .B(G85gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT80), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n276), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n280), .B1(new_n259), .B2(new_n270), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT80), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT79), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n244), .B(new_n257), .C1(new_n247), .C2(new_n251), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n276), .B1(new_n284), .B2(new_n246), .ZN(new_n285));
  AOI211_X1 g084(.A(new_n283), .B(KEYINPUT6), .C1(new_n285), .C2(new_n270), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n259), .A2(new_n270), .A3(new_n280), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT79), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n279), .B(new_n282), .C1(new_n286), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT81), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n288), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n283), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n287), .A2(KEYINPUT79), .A3(new_n288), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n281), .B(new_n278), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT81), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n271), .A2(KEYINPUT6), .A3(new_n276), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n291), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT26), .ZN(new_n302));
  INV_X1    g101(.A(G169gat), .ZN(new_n303));
  INV_X1    g102(.A(G176gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n305), .A2(KEYINPUT65), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  NOR3_X1   g108(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT65), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G183gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT27), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT27), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G183gat), .ZN(new_n317));
  INV_X1    g116(.A(G190gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT28), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT27), .B(G183gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(KEYINPUT28), .A3(new_n318), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n313), .A2(new_n324), .A3(KEYINPUT66), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT66), .B1(new_n313), .B2(new_n324), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(G169gat), .B2(G176gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n318), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n330), .A3(new_n306), .ZN(new_n331));
  NAND2_X1  g130(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G190gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT23), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT64), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n336), .B(new_n337), .C1(new_n338), .C2(KEYINPUT25), .ZN(new_n339));
  AND2_X1   g138(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n340), .A2(new_n318), .B1(G169gat), .B2(G176gat), .ZN(new_n341));
  OR2_X1    g140(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(G190gat), .A3(new_n332), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n341), .A2(new_n343), .A3(new_n338), .A4(new_n329), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n341), .A2(new_n343), .A3(new_n329), .A4(new_n337), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT25), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT29), .B1(new_n327), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n301), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n339), .A2(new_n347), .B1(new_n324), .B2(new_n313), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(KEYINPUT72), .A3(new_n351), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n356), .B1(new_n353), .B2(new_n350), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n313), .A2(new_n324), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT66), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n313), .A2(new_n324), .A3(KEYINPUT66), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n348), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n365), .A2(KEYINPUT71), .A3(new_n350), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n352), .A2(new_n358), .A3(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(G211gat), .B(G218gat), .Z(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT70), .B(G197gat), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n370), .A2(G204gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(G204gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n369), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  AOI211_X1 g175(.A(new_n368), .B(new_n374), .C1(new_n371), .C2(new_n372), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n367), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n348), .B2(new_n359), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT73), .B1(new_n380), .B2(new_n351), .ZN(new_n381));
  INV_X1    g180(.A(new_n378), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n363), .A2(new_n351), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT73), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n384), .B(new_n350), .C1(new_n353), .C2(KEYINPUT29), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n381), .A2(new_n382), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(G8gat), .B(G36gat), .Z(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT74), .ZN(new_n388));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT30), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n379), .A2(new_n386), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n386), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n395), .B1(new_n378), .B2(new_n367), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n394), .B1(new_n396), .B2(new_n390), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT30), .B1(new_n396), .B2(new_n390), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n300), .A2(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(KEYINPUT31), .B(G50gat), .Z(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT82), .ZN(new_n402));
  XOR2_X1   g201(.A(G78gat), .B(G106gat), .Z(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G22gat), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n364), .B1(new_n376), .B2(new_n377), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n264), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n239), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n263), .A2(KEYINPUT29), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n409), .A2(new_n376), .A3(new_n377), .ZN(new_n410));
  AND2_X1   g209(.A1(G228gat), .A2(G233gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n250), .B1(new_n406), .B2(new_n255), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n412), .B1(new_n415), .B2(new_n410), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n405), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n404), .B1(new_n417), .B2(KEYINPUT83), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n414), .A2(new_n416), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G22gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n414), .A2(new_n416), .A3(new_n405), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT83), .A4(new_n404), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n363), .A2(new_n249), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n327), .A2(new_n254), .A3(new_n348), .ZN(new_n427));
  AND2_X1   g226(.A1(G227gat), .A2(G233gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(G15gat), .B(G43gat), .Z(new_n432));
  XNOR2_X1  g231(.A(G71gat), .B(G99gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n428), .B1(new_n426), .B2(new_n427), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT34), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI211_X1 g237(.A(KEYINPUT34), .B(new_n428), .C1(new_n426), .C2(new_n427), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n435), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n436), .A2(new_n437), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n431), .B(new_n434), .C1(new_n442), .C2(new_n439), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n429), .A2(KEYINPUT32), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n441), .B2(new_n443), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT36), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT36), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n449), .B1(new_n445), .B2(new_n446), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n400), .A2(new_n425), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n425), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n262), .A2(new_n269), .A3(new_n257), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n245), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT84), .B1(new_n243), .B2(new_n245), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT84), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n238), .A2(new_n242), .A3(new_n457), .A4(new_n244), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n455), .A2(KEYINPUT39), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n460), .A2(KEYINPUT40), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT39), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n454), .A2(new_n463), .A3(new_n245), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n459), .A2(new_n280), .A3(new_n462), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n280), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n456), .A2(KEYINPUT39), .A3(new_n458), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n467), .B1(new_n454), .B2(new_n245), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n461), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n465), .A2(new_n277), .A3(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n453), .B(new_n470), .C1(new_n397), .C2(new_n398), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n379), .A2(new_n386), .A3(new_n390), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n392), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n379), .A2(new_n386), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n391), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n476), .A3(new_n394), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n453), .B1(new_n477), .B2(new_n470), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n452), .B1(new_n472), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT38), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n391), .A2(KEYINPUT37), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n475), .A2(KEYINPUT37), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n367), .A2(new_n382), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n381), .A2(new_n378), .A3(new_n383), .A4(new_n385), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n486), .A2(KEYINPUT37), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT38), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n390), .B1(new_n379), .B2(new_n386), .ZN(new_n489));
  INV_X1    g288(.A(new_n481), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g290(.A(KEYINPUT87), .B(new_n299), .C1(new_n292), .C2(new_n281), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n281), .A2(new_n493), .A3(KEYINPUT6), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n492), .A2(new_n494), .B1(new_n396), .B2(new_n390), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n491), .A2(new_n495), .A3(KEYINPUT88), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n484), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n451), .B1(new_n479), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n452), .A2(new_n447), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT35), .B1(new_n400), .B2(new_n502), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n425), .A2(new_n445), .A3(new_n446), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT35), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n492), .A2(new_n505), .A3(new_n494), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n477), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n501), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT93), .ZN(new_n511));
  XNOR2_X1  g310(.A(G113gat), .B(G141gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(G197gat), .ZN(new_n513));
  XOR2_X1   g312(.A(KEYINPUT11), .B(G169gat), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(new_n515), .B(KEYINPUT12), .Z(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(G29gat), .A2(G36gat), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n518), .B(KEYINPUT14), .Z(new_n519));
  XOR2_X1   g318(.A(KEYINPUT89), .B(G36gat), .Z(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(G29gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(KEYINPUT15), .A3(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G43gat), .B(G50gat), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n519), .A2(new_n521), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n524), .B1(KEYINPUT15), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n522), .A2(new_n523), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530));
  INV_X1    g329(.A(G1gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT16), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(G1gat), .B2(new_n530), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(G8gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n529), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT91), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n529), .B2(new_n537), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n539), .A2(new_n541), .B1(new_n529), .B2(new_n537), .ZN(new_n542));
  NAND2_X1  g341(.A1(G229gat), .A2(G233gat), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n543), .B(KEYINPUT13), .Z(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n539), .A2(new_n541), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n529), .A2(KEYINPUT17), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n535), .B1(new_n528), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(KEYINPUT18), .A3(new_n543), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT18), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n549), .A2(new_n553), .ZN(new_n557));
  INV_X1    g356(.A(new_n543), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n517), .B1(new_n548), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n546), .A2(new_n547), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n542), .A2(KEYINPUT92), .A3(new_n545), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n555), .A2(new_n559), .ZN(new_n565));
  NOR3_X1   g364(.A1(new_n564), .A2(new_n565), .A3(new_n516), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n511), .B1(new_n561), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n516), .B1(new_n564), .B2(new_n565), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n548), .A2(new_n560), .A3(new_n517), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT93), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G85gat), .A2(G92gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT7), .ZN(new_n574));
  NAND2_X1  g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  INV_X1    g374(.A(G85gat), .ZN(new_n576));
  INV_X1    g375(.A(G92gat), .ZN(new_n577));
  AOI22_X1  g376(.A1(KEYINPUT8), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G99gat), .B(G106gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n581), .B1(new_n528), .B2(new_n551), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n550), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n528), .A2(new_n581), .B1(KEYINPUT41), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n584), .A2(KEYINPUT41), .ZN(new_n589));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n588), .B(new_n591), .Z(new_n592));
  AND2_X1   g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n593), .A2(KEYINPUT9), .ZN(new_n594));
  XOR2_X1   g393(.A(G57gat), .B(G64gat), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G71gat), .B(G78gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G127gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n598), .B(KEYINPUT94), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n537), .B1(new_n605), .B2(new_n599), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n603), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G155gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n607), .B(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n592), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n581), .B(new_n598), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT10), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n581), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(G230gat), .ZN(new_n619));
  INV_X1    g418(.A(G233gat), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OR3_X1    g420(.A1(new_n614), .A2(new_n619), .A3(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n623), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT95), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n630), .ZN(new_n631));
  OR3_X1    g430(.A1(new_n510), .A2(new_n572), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(new_n300), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n531), .ZN(G1324gat));
  NOR2_X1   g433(.A1(new_n632), .A2(new_n399), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT16), .B(G8gat), .Z(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(G8gat), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n637), .B1(new_n638), .B2(new_n635), .ZN(new_n639));
  MUX2_X1   g438(.A(new_n637), .B(new_n639), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g439(.A1(new_n448), .A2(new_n450), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT96), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n448), .A2(KEYINPUT96), .A3(new_n450), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(G15gat), .B1(new_n632), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n447), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n647), .A2(G15gat), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n646), .B1(new_n632), .B2(new_n648), .ZN(G1326gat));
  NOR2_X1   g448(.A1(new_n632), .A2(new_n452), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT43), .B(G22gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  INV_X1    g451(.A(new_n592), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n630), .A2(new_n612), .ZN(new_n654));
  NOR4_X1   g453(.A1(new_n510), .A2(new_n572), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(G29gat), .ZN(new_n656));
  INV_X1    g455(.A(new_n300), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT45), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT44), .B1(new_n510), .B2(new_n653), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT97), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n290), .A2(KEYINPUT81), .B1(KEYINPUT6), .B2(new_n281), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n477), .B1(new_n298), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n505), .B1(new_n663), .B2(new_n504), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n504), .A2(new_n507), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n503), .A2(new_n508), .A3(KEYINPUT97), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n501), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n653), .A2(KEYINPUT44), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n668), .A2(KEYINPUT98), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT98), .B1(new_n668), .B2(new_n669), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n660), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n568), .A2(new_n569), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n654), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G29gat), .B1(new_n676), .B2(new_n300), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n659), .A2(new_n677), .ZN(G1328gat));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n520), .B1(new_n679), .B2(KEYINPUT46), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n655), .A2(new_n477), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n679), .A2(KEYINPUT46), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n520), .B1(new_n676), .B2(new_n399), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(G1329gat));
  OAI21_X1  g484(.A(G43gat), .B1(new_n676), .B2(new_n641), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n647), .A2(G43gat), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n655), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n686), .A2(KEYINPUT47), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n645), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n672), .A2(new_n690), .A3(new_n675), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n691), .A2(KEYINPUT100), .A3(G43gat), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n688), .B(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT100), .B1(new_n691), .B2(G43gat), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n692), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n689), .B1(new_n696), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g496(.A1(new_n672), .A2(new_n425), .A3(new_n675), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n452), .A2(G50gat), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n698), .A2(G50gat), .B1(new_n655), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT48), .ZN(G1331gat));
  AND3_X1   g500(.A1(new_n674), .A2(new_n613), .A3(new_n629), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n668), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n657), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g505(.A1(new_n399), .A2(KEYINPUT102), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n399), .A2(KEYINPUT102), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  AND2_X1   g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n711), .B2(new_n712), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n703), .B2(new_n645), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n647), .A2(G71gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n703), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT103), .B(KEYINPUT50), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1334gat));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n425), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G78gat), .ZN(G1335gat));
  INV_X1    g521(.A(KEYINPUT51), .ZN(new_n723));
  INV_X1    g522(.A(new_n612), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n673), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n668), .A2(new_n592), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n668), .A2(KEYINPUT104), .A3(new_n592), .A4(new_n725), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n668), .A2(new_n674), .A3(new_n612), .A4(new_n592), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n723), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n733), .A2(new_n576), .A3(new_n657), .A4(new_n629), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n673), .A2(new_n724), .A3(new_n630), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n672), .A2(new_n735), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n736), .A2(new_n657), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n734), .B1(new_n737), .B2(new_n576), .ZN(G1336gat));
  AOI21_X1  g537(.A(new_n577), .B1(new_n736), .B2(new_n477), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n732), .A2(new_n726), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n710), .A2(G92gat), .A3(new_n630), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT52), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n733), .A2(new_n745), .A3(new_n741), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n728), .A2(new_n729), .B1(new_n723), .B2(new_n731), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT105), .B1(new_n747), .B2(new_n742), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT106), .B(KEYINPUT52), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n672), .A2(new_n709), .A3(new_n735), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(G92gat), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n749), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n750), .B1(new_n749), .B2(new_n753), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n744), .B1(new_n754), .B2(new_n755), .ZN(G1337gat));
  INV_X1    g555(.A(G99gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n736), .A2(new_n690), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n759), .B2(new_n758), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n733), .A2(new_n757), .A3(new_n447), .A4(new_n629), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1338gat));
  INV_X1    g562(.A(G106gat), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n736), .B2(new_n425), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n629), .A2(new_n764), .A3(new_n425), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n740), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT53), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n747), .B2(new_n766), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n765), .B2(new_n770), .ZN(G1339gat));
  NOR2_X1   g570(.A1(new_n554), .A2(new_n543), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n542), .A2(new_n545), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n515), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n569), .A2(new_n629), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n616), .A2(G230gat), .A3(G233gat), .A4(new_n617), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n621), .A2(KEYINPUT54), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n626), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n777), .B(new_n778), .C1(KEYINPUT54), .C2(new_n621), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n621), .A2(new_n622), .A3(new_n626), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n780), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n568), .B2(new_n569), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n653), .B1(new_n775), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n569), .A2(new_n774), .ZN(new_n787));
  INV_X1    g586(.A(new_n784), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n592), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n724), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n631), .A2(new_n673), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(new_n300), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n709), .A2(new_n502), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G113gat), .B1(new_n795), .B2(new_n572), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT109), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n795), .B(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n799), .A2(new_n214), .A3(new_n673), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n797), .A2(new_n800), .ZN(G1340gat));
  OAI21_X1  g600(.A(G120gat), .B1(new_n795), .B2(new_n630), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT111), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n799), .A2(new_n212), .A3(new_n629), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1341gat));
  OAI21_X1  g605(.A(KEYINPUT112), .B1(new_n795), .B2(new_n612), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n793), .A2(new_n808), .A3(new_n724), .A4(new_n794), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n203), .A2(new_n204), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n810), .B(new_n811), .ZN(G1342gat));
  NAND2_X1  g611(.A1(new_n592), .A2(new_n399), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n504), .A2(new_n207), .A3(new_n209), .ZN(new_n814));
  NOR4_X1   g613(.A1(new_n792), .A2(new_n300), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT56), .ZN(new_n816));
  OAI21_X1  g615(.A(G134gat), .B1(new_n795), .B2(new_n653), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1343gat));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n819), .B(new_n425), .C1(new_n790), .C2(new_n791), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n710), .A2(new_n657), .A3(new_n641), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  XOR2_X1   g622(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n824));
  AOI21_X1  g623(.A(new_n824), .B1(new_n779), .B2(KEYINPUT113), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n825), .B1(KEYINPUT113), .B2(new_n779), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n782), .A3(new_n781), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT93), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT93), .B1(new_n568), .B2(new_n569), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n569), .A2(new_n629), .A3(new_n774), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n592), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n787), .A2(new_n592), .A3(new_n788), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n612), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n791), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n452), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n823), .B(new_n571), .C1(new_n837), .C2(new_n819), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G141gat), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n840), .B(new_n657), .C1(new_n790), .C2(new_n791), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n425), .A3(new_n645), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n673), .A2(new_n788), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n592), .B1(new_n843), .B2(new_n832), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n612), .B1(new_n844), .B2(new_n834), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n836), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n840), .B1(new_n846), .B2(new_n657), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n571), .A2(new_n226), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n850), .B(KEYINPUT116), .Z(new_n851));
  NAND4_X1  g650(.A1(new_n848), .A2(new_n849), .A3(new_n710), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n839), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n823), .B1(new_n837), .B2(new_n819), .ZN(new_n855));
  OAI211_X1 g654(.A(KEYINPUT58), .B(G141gat), .C1(new_n855), .C2(new_n674), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n842), .A2(new_n847), .A3(new_n709), .ZN(new_n857));
  AOI22_X1  g656(.A1(new_n857), .A2(new_n851), .B1(new_n849), .B2(new_n854), .ZN(new_n858));
  AOI22_X1  g657(.A1(new_n853), .A2(new_n854), .B1(new_n856), .B2(new_n858), .ZN(G1344gat));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n228), .A3(new_n629), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n820), .A2(new_n822), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n827), .B1(new_n567), .B2(new_n570), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n653), .B1(new_n862), .B2(new_n775), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n724), .B1(new_n863), .B2(new_n789), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n425), .B1(new_n864), .B2(new_n791), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n861), .B1(new_n865), .B2(KEYINPUT57), .ZN(new_n866));
  AOI211_X1 g665(.A(KEYINPUT59), .B(new_n228), .C1(new_n866), .C2(new_n629), .ZN(new_n867));
  XNOR2_X1  g666(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n452), .A2(KEYINPUT57), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n571), .A2(new_n631), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT57), .B1(new_n792), .B2(new_n452), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n821), .A2(KEYINPUT119), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n630), .B1(new_n821), .B2(KEYINPUT119), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n871), .A2(new_n872), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n868), .B1(new_n875), .B2(G148gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n860), .B1(new_n867), .B2(new_n876), .ZN(G1345gat));
  OAI21_X1  g676(.A(G155gat), .B1(new_n855), .B2(new_n612), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n857), .A2(new_n232), .A3(new_n724), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1346gat));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n233), .B1(new_n866), .B2(new_n592), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n813), .A2(G162gat), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n848), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n881), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(G162gat), .B1(new_n855), .B2(new_n653), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n848), .A2(new_n883), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(KEYINPUT120), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(new_n888), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n792), .A2(new_n657), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n710), .A2(new_n502), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(KEYINPUT121), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n846), .A2(new_n300), .A3(new_n891), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n892), .A2(new_n895), .A3(new_n303), .A4(new_n673), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n846), .A2(new_n300), .A3(new_n477), .A4(new_n504), .ZN(new_n897));
  OAI21_X1  g696(.A(G169gat), .B1(new_n897), .B2(new_n572), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT122), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n896), .A2(new_n901), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1348gat));
  NAND4_X1  g702(.A1(new_n892), .A2(new_n895), .A3(new_n304), .A4(new_n629), .ZN(new_n904));
  OAI21_X1  g703(.A(G176gat), .B1(new_n897), .B2(new_n630), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n904), .A2(KEYINPUT123), .A3(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1349gat));
  OAI21_X1  g709(.A(G183gat), .B1(new_n897), .B2(new_n612), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n724), .A2(new_n322), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n911), .B(new_n912), .C1(new_n893), .C2(new_n913), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n897), .B2(new_n653), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n916), .A2(KEYINPUT61), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(KEYINPUT61), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n892), .A2(new_n895), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n592), .A2(new_n318), .ZN(new_n920));
  OAI22_X1  g719(.A1(new_n917), .A2(new_n918), .B1(new_n919), .B2(new_n920), .ZN(G1351gat));
  INV_X1    g720(.A(G197gat), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n690), .A2(new_n657), .A3(new_n399), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n871), .A2(new_n872), .A3(new_n571), .A4(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n925), .B2(new_n924), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n690), .A2(new_n452), .A3(new_n710), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n928), .A2(KEYINPUT125), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(KEYINPUT125), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n890), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n922), .A3(new_n673), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n927), .A2(new_n933), .ZN(G1352gat));
  OR2_X1    g733(.A1(new_n630), .A2(G204gat), .ZN(new_n935));
  OR3_X1    g734(.A1(new_n931), .A2(KEYINPUT62), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n871), .A2(new_n872), .A3(new_n923), .ZN(new_n937));
  OAI21_X1  g736(.A(G204gat), .B1(new_n937), .B2(new_n630), .ZN(new_n938));
  OAI21_X1  g737(.A(KEYINPUT62), .B1(new_n931), .B2(new_n935), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(G1353gat));
  OR3_X1    g739(.A1(new_n931), .A2(G211gat), .A3(new_n612), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n871), .A2(new_n872), .A3(new_n724), .A4(new_n923), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n942), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT63), .B1(new_n942), .B2(G211gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(G1354gat));
  NAND4_X1  g744(.A1(new_n871), .A2(new_n872), .A3(new_n592), .A4(new_n923), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G218gat), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n653), .A2(G218gat), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT127), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n947), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1355gat));
endmodule


