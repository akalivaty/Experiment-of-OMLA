//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1350, new_n1351,
    new_n1352, new_n1353, new_n1354, new_n1355, new_n1356, new_n1357,
    new_n1358, new_n1359, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1423, new_n1424,
    new_n1425, new_n1426, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1432, new_n1433, new_n1434, new_n1435, new_n1436, new_n1437,
    new_n1438, new_n1439, new_n1440;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n211), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT65), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n220), .B1(new_n211), .B2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G13), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n222), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  AND2_X1   g0026(.A1(KEYINPUT66), .A2(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(KEYINPUT66), .A2(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n206), .A2(new_n207), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n219), .B(new_n226), .C1(new_n231), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n207), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n203), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n244), .B(new_n249), .ZN(G351));
  NAND2_X1  g0050(.A1(G33), .A2(G97), .ZN(new_n251));
  INV_X1    g0051(.A(G232), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G1698), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(G226), .B2(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n251), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(KEYINPUT71), .A3(new_n230), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT71), .ZN(new_n263));
  AND2_X1   g0063(.A1(G1), .A2(G13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT13), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n270), .A2(new_n273), .B1(new_n264), .B2(new_n265), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT67), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n271), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT67), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n272), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G1), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n274), .A2(G238), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n268), .A2(new_n269), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT73), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n278), .A2(new_n280), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n274), .A2(G238), .ZN(new_n286));
  INV_X1    g0086(.A(new_n251), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G226), .A2(G1698), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n252), .B2(G1698), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n287), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(KEYINPUT71), .B1(new_n261), .B2(new_n230), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n264), .A2(new_n263), .A3(new_n265), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n285), .B(new_n286), .C1(new_n291), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT13), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n268), .A2(KEYINPUT73), .A3(new_n269), .A4(new_n281), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n284), .A2(G190), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(KEYINPUT74), .A2(KEYINPUT12), .ZN(new_n299));
  NAND2_X1  g0099(.A1(KEYINPUT74), .A2(KEYINPUT12), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n270), .A2(G13), .A3(G20), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n299), .B(new_n300), .C1(new_n301), .C2(G68), .ZN(new_n302));
  INV_X1    g0102(.A(new_n301), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n203), .ZN(new_n304));
  OAI211_X1 g0104(.A(KEYINPUT75), .B(new_n302), .C1(new_n304), .C2(KEYINPUT12), .ZN(new_n305));
  NAND3_X1  g0105(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n230), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G20), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G1), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n308), .A2(G68), .A3(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n305), .B(new_n312), .C1(KEYINPUT75), .C2(new_n302), .ZN(new_n313));
  NOR2_X1   g0113(.A1(G20), .A2(G33), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n314), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n229), .A2(G33), .ZN(new_n316));
  INV_X1    g0116(.A(G77), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n318), .A2(KEYINPUT11), .A3(new_n307), .ZN(new_n319));
  AOI21_X1  g0119(.A(KEYINPUT11), .B1(new_n318), .B2(new_n307), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n313), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n282), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n269), .B1(new_n268), .B2(new_n281), .ZN(new_n323));
  OAI21_X1  g0123(.A(G200), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n298), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G179), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n326), .B1(new_n295), .B2(KEYINPUT13), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n284), .A2(new_n327), .A3(new_n297), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n296), .A2(new_n282), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT14), .B1(new_n329), .B2(G169), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT14), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  AOI211_X1 g0132(.A(new_n331), .B(new_n332), .C1(new_n296), .C2(new_n282), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n328), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n321), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n325), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G1698), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n290), .A2(G232), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G107), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(new_n290), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT70), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n259), .B2(new_n337), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n290), .A2(KEYINPUT70), .A3(G1698), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n340), .B1(new_n344), .B2(G238), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n294), .ZN(new_n346));
  INV_X1    g0146(.A(new_n274), .ZN(new_n347));
  INV_X1    g0147(.A(G244), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n285), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n326), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT66), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n309), .ZN(new_n353));
  NAND2_X1  g0153(.A1(KEYINPUT66), .A2(G20), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(new_n255), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT15), .B(G87), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n356), .A2(new_n358), .B1(G77), .B2(new_n355), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT8), .B(G58), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT72), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n309), .A2(new_n255), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n307), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n310), .A2(new_n317), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n308), .A2(new_n365), .B1(new_n317), .B2(new_n303), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n332), .B1(new_n346), .B2(new_n349), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n351), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G200), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n350), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n350), .A2(G190), .ZN(new_n372));
  INV_X1    g0172(.A(new_n367), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n336), .B(new_n369), .C1(new_n371), .C2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT69), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n290), .A2(new_n376), .A3(G222), .A4(new_n337), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n290), .A2(G222), .A3(new_n337), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT69), .B1(new_n259), .B2(G77), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G223), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n342), .B2(new_n343), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n267), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  XOR2_X1   g0183(.A(KEYINPUT68), .B(G226), .Z(new_n384));
  AOI22_X1  g0184(.A1(new_n274), .A2(new_n384), .B1(new_n278), .B2(new_n280), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(G179), .ZN(new_n387));
  INV_X1    g0187(.A(new_n307), .ZN(new_n388));
  INV_X1    g0188(.A(new_n360), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n356), .A2(new_n389), .B1(G150), .B2(new_n314), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n208), .A2(G20), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n388), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n388), .A2(new_n301), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n311), .A2(G50), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n393), .A2(new_n394), .B1(G50), .B2(new_n301), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(G169), .B1(new_n383), .B2(new_n385), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n387), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT10), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n386), .A2(G200), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT9), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n392), .B2(new_n395), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n390), .A2(new_n391), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n307), .ZN(new_n405));
  INV_X1    g0205(.A(new_n395), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(KEYINPUT9), .A3(new_n406), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n401), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n383), .A2(G190), .A3(new_n385), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n400), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n407), .A2(new_n403), .ZN(new_n411));
  AND4_X1   g0211(.A1(new_n400), .A2(new_n411), .A3(new_n409), .A4(new_n401), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n399), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n389), .A2(new_n311), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n393), .B1(new_n414), .B2(KEYINPUT77), .ZN(new_n415));
  OR3_X1    g0215(.A1(new_n360), .A2(KEYINPUT77), .A3(new_n310), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n415), .A2(new_n416), .B1(new_n303), .B2(new_n360), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT76), .B1(new_n257), .B2(G33), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT76), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(new_n255), .A3(KEYINPUT3), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(new_n420), .A3(new_n258), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT7), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n227), .A2(new_n228), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n422), .B1(new_n290), .B2(G20), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G68), .ZN(new_n427));
  INV_X1    g0227(.A(G159), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n362), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G58), .A2(G68), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n204), .A2(new_n205), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n429), .B1(new_n431), .B2(G20), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT16), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(G20), .B1(new_n256), .B2(new_n258), .ZN(new_n434));
  OAI21_X1  g0234(.A(G68), .B1(new_n434), .B2(new_n422), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n353), .A2(new_n422), .A3(new_n354), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(new_n290), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n432), .B(KEYINPUT16), .C1(new_n435), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n307), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n417), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n256), .A2(new_n258), .A3(G223), .A4(new_n337), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G87), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n256), .A2(new_n258), .A3(G226), .A4(G1698), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n441), .B(new_n442), .C1(new_n443), .C2(KEYINPUT78), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n443), .A2(KEYINPUT78), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n267), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n274), .A2(G232), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n285), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(G179), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n443), .A2(KEYINPUT78), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT78), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n290), .A2(new_n452), .A3(G226), .A4(G1698), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n451), .A2(new_n453), .A3(new_n441), .A4(new_n442), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n448), .B1(new_n454), .B2(new_n267), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n450), .B1(new_n332), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n440), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT18), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT17), .ZN(new_n459));
  INV_X1    g0259(.A(G190), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n446), .A2(new_n460), .A3(new_n449), .ZN(new_n461));
  AOI21_X1  g0261(.A(G200), .B1(new_n446), .B2(new_n449), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n459), .B1(new_n463), .B2(new_n440), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT18), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n440), .A2(new_n465), .A3(new_n456), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n414), .A2(KEYINPUT77), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(new_n416), .A3(new_n308), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n301), .B2(new_n389), .ZN(new_n469));
  INV_X1    g0269(.A(new_n439), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT16), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n203), .B1(new_n424), .B2(new_n425), .ZN(new_n472));
  INV_X1    g0272(.A(new_n432), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n469), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n446), .A2(new_n460), .A3(new_n449), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(G200), .B2(new_n455), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(KEYINPUT17), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n458), .A2(new_n464), .A3(new_n466), .A4(new_n478), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n375), .A2(new_n413), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n256), .A2(new_n258), .A3(G244), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(new_n348), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n484), .A2(new_n337), .A3(new_n256), .A4(new_n258), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n256), .A2(new_n258), .A3(G250), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n337), .B1(new_n488), .B2(KEYINPUT4), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n267), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT81), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n264), .A2(new_n265), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT5), .B1(new_n276), .B2(new_n277), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT5), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n270), .B(G45), .C1(new_n495), .C2(G41), .ZN(new_n496));
  OAI211_X1 g0296(.A(G257), .B(new_n493), .C1(new_n494), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT82), .ZN(new_n498));
  INV_X1    g0298(.A(new_n496), .ZN(new_n499));
  AND2_X1   g0299(.A1(KEYINPUT67), .A2(G41), .ZN(new_n500));
  NOR2_X1   g0300(.A1(KEYINPUT67), .A2(G41), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n495), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT82), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n503), .A2(new_n504), .A3(G257), .A4(new_n493), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n494), .A2(new_n496), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n261), .A2(new_n230), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(new_n279), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n498), .A2(new_n505), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(KEYINPUT81), .B(new_n267), .C1(new_n487), .C2(new_n489), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n492), .A2(new_n509), .A3(new_n326), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n498), .A2(new_n505), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n506), .A2(new_n508), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n490), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n332), .ZN(new_n515));
  AND2_X1   g0315(.A1(G97), .A2(G107), .ZN(new_n516));
  NOR2_X1   g0316(.A1(G97), .A2(G107), .ZN(new_n517));
  OAI22_X1  g0317(.A1(new_n516), .A2(new_n517), .B1(KEYINPUT79), .B2(KEYINPUT6), .ZN(new_n518));
  NOR2_X1   g0318(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g0319(.A(G97), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n519), .B1(KEYINPUT6), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g0321(.A(G97), .B(G107), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI22_X1  g0323(.A1(new_n523), .A2(new_n229), .B1(new_n317), .B2(new_n362), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n339), .B1(new_n424), .B2(new_n425), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n307), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n270), .A2(G33), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n301), .A2(new_n527), .A3(new_n230), .A4(new_n306), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G97), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n301), .A2(new_n520), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT80), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n529), .A2(KEYINPUT80), .A3(new_n530), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n526), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n511), .A2(new_n515), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT83), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n514), .A2(new_n332), .B1(new_n526), .B2(new_n535), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(KEYINPUT83), .A3(new_n511), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n492), .A2(new_n509), .A3(new_n510), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G200), .ZN(new_n543));
  INV_X1    g0343(.A(new_n536), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n512), .A2(new_n490), .A3(new_n513), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G190), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n539), .A2(new_n541), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT25), .B1(new_n303), .B2(new_n339), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n303), .A2(KEYINPUT25), .A3(new_n339), .ZN(new_n551));
  INV_X1    g0351(.A(new_n528), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n550), .A2(new_n551), .B1(G107), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n355), .A2(new_n259), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT22), .B1(new_n555), .B2(G87), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n229), .A2(new_n290), .A3(KEYINPUT22), .A4(G87), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n355), .A2(new_n558), .A3(new_n339), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT24), .ZN(new_n560));
  OAI22_X1  g0360(.A1(new_n558), .A2(new_n339), .B1(new_n560), .B2(KEYINPUT85), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G33), .A2(G116), .ZN(new_n562));
  AOI21_X1  g0362(.A(G20), .B1(new_n562), .B2(new_n558), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n557), .A2(new_n559), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT85), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n556), .A2(new_n565), .B1(new_n566), .B2(KEYINPUT24), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n559), .A2(new_n564), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT22), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n229), .A2(new_n290), .ZN(new_n570));
  INV_X1    g0370(.A(G87), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n566), .A2(KEYINPUT24), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n568), .A2(new_n572), .A3(new_n573), .A4(new_n557), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n554), .B1(new_n575), .B2(new_n307), .ZN(new_n576));
  OAI211_X1 g0376(.A(G264), .B(new_n493), .C1(new_n494), .C2(new_n496), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT86), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n507), .B1(new_n499), .B2(new_n502), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(KEYINPUT86), .A3(G264), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n290), .A2(G257), .A3(G1698), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n256), .A2(new_n258), .A3(G250), .A4(new_n337), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G294), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n586), .A2(new_n267), .B1(new_n506), .B2(new_n508), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G169), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n582), .A2(G179), .A3(new_n587), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT87), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n576), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(KEYINPUT87), .A3(new_n590), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n588), .A2(new_n370), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G190), .B2(new_n588), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n593), .A2(new_n594), .B1(new_n576), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n255), .A2(G97), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n353), .A2(new_n598), .A3(new_n354), .A4(new_n486), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n306), .A2(new_n230), .B1(G20), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT20), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n599), .A2(KEYINPUT20), .A3(new_n601), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n301), .A2(G116), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n552), .B2(G116), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n290), .A2(G264), .A3(G1698), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n259), .A2(G303), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n256), .A2(new_n258), .A3(G257), .A4(new_n337), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n267), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n580), .A2(G270), .B1(new_n506), .B2(new_n508), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n609), .A2(G179), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n614), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(new_n609), .A3(G169), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT21), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT21), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n618), .A2(new_n609), .A3(new_n621), .A4(G169), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n617), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  AND4_X1   g0423(.A1(KEYINPUT84), .A2(new_n571), .A3(new_n520), .A4(new_n339), .ZN(new_n624));
  NOR2_X1   g0424(.A1(G87), .A2(G97), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT84), .B1(new_n625), .B2(new_n339), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT19), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n251), .A2(new_n627), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n624), .A2(new_n626), .B1(new_n355), .B2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n353), .A2(G33), .A3(G97), .A4(new_n354), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n627), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n229), .A2(new_n290), .A3(G68), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n307), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n357), .A2(new_n303), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n552), .A2(new_n358), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n280), .A2(G45), .ZN(new_n638));
  OAI21_X1  g0438(.A(G250), .B1(new_n272), .B2(G1), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n507), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n256), .A2(new_n258), .A3(G244), .A4(G1698), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n256), .A2(new_n258), .A3(G238), .A4(new_n337), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n642), .A3(new_n562), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n640), .B1(new_n643), .B2(new_n267), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n326), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(G169), .B2(new_n644), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n643), .A2(new_n267), .ZN(new_n647));
  INV_X1    g0447(.A(new_n640), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G190), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n370), .B2(new_n644), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n552), .A2(G87), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n634), .A2(new_n635), .A3(new_n651), .ZN(new_n652));
  OAI22_X1  g0452(.A1(new_n637), .A2(new_n646), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n609), .B1(new_n618), .B2(G200), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n460), .B2(new_n618), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n623), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  AND4_X1   g0457(.A1(new_n480), .A2(new_n548), .A3(new_n597), .A4(new_n657), .ZN(G372));
  AND3_X1   g0458(.A1(new_n440), .A2(new_n465), .A3(new_n456), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n465), .B1(new_n440), .B2(new_n456), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n369), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n298), .A2(new_n321), .A3(new_n324), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n662), .A2(new_n663), .B1(new_n335), .B2(new_n334), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n463), .A2(new_n440), .A3(new_n459), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT17), .B1(new_n475), .B2(new_n477), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n661), .B1(new_n664), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n411), .A2(new_n409), .A3(new_n401), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT10), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n408), .A2(new_n400), .A3(new_n409), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n398), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n480), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n676));
  INV_X1    g0476(.A(new_n644), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n332), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n676), .A2(new_n678), .A3(new_n645), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(G200), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n633), .A2(new_n307), .B1(new_n303), .B2(new_n357), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(new_n651), .A4(new_n649), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n540), .A2(new_n511), .A3(new_n679), .A4(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n679), .B1(new_n683), .B2(KEYINPUT26), .ZN(new_n684));
  AND4_X1   g0484(.A1(KEYINPUT83), .A2(new_n511), .A3(new_n515), .A4(new_n536), .ZN(new_n685));
  AOI21_X1  g0485(.A(KEYINPUT83), .B1(new_n540), .B2(new_n511), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n654), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n684), .B1(new_n687), .B2(KEYINPUT26), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n685), .A2(new_n686), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n575), .A2(new_n307), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n553), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n591), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n623), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n653), .B1(new_n576), .B2(new_n596), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n689), .A2(new_n547), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n688), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n674), .B1(new_n675), .B2(new_n697), .ZN(G369));
  NOR2_X1   g0498(.A1(new_n222), .A2(G1), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n229), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT27), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n229), .A2(new_n702), .A3(new_n699), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(G213), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G343), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n609), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n623), .A2(new_n656), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT88), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n708), .B(new_n709), .C1(new_n623), .C2(new_n707), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n620), .A2(new_n622), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n616), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(KEYINPUT88), .A3(new_n609), .A4(new_n706), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(G330), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n590), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n332), .B1(new_n582), .B2(new_n587), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n592), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n691), .A3(new_n594), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n596), .A2(new_n576), .ZN(new_n719));
  INV_X1    g0519(.A(new_n706), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n718), .B(new_n719), .C1(new_n576), .C2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n593), .A2(new_n594), .A3(new_n706), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n714), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT89), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n706), .B(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n692), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n623), .A2(new_n706), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n597), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n726), .A2(new_n731), .ZN(G399));
  NOR3_X1   g0532(.A1(new_n624), .A2(new_n626), .A3(G116), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT90), .ZN(new_n734));
  INV_X1    g0534(.A(new_n224), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n276), .A2(new_n277), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n270), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n734), .A2(new_n738), .B1(new_n232), .B2(new_n737), .ZN(new_n739));
  XNOR2_X1  g0539(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n694), .A2(new_n539), .A3(new_n541), .A4(new_n547), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n718), .A2(new_n623), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n679), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n683), .B2(KEYINPUT26), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(new_n687), .B2(KEYINPUT26), .ZN(new_n747));
  OAI211_X1 g0547(.A(KEYINPUT29), .B(new_n720), .C1(new_n744), .C2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n728), .B1(new_n688), .B2(new_n695), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n748), .B1(KEYINPUT29), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n326), .B1(new_n586), .B2(new_n267), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n577), .A2(new_n578), .ZN(new_n752));
  AOI21_X1  g0552(.A(KEYINPUT86), .B1(new_n580), .B2(G264), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n615), .A2(new_n644), .A3(new_n614), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n545), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT30), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n756), .A2(KEYINPUT30), .A3(new_n545), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n644), .A2(G179), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n542), .A2(new_n588), .A3(new_n618), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n728), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT31), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n763), .A2(KEYINPUT92), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(KEYINPUT92), .B1(new_n763), .B2(new_n766), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n548), .A2(new_n597), .A3(new_n657), .A4(new_n764), .ZN(new_n770));
  AOI21_X1  g0570(.A(KEYINPUT30), .B1(new_n756), .B2(new_n545), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT93), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n760), .B(new_n762), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n514), .A2(new_n754), .A3(new_n755), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n774), .A2(KEYINPUT93), .A3(KEYINPUT30), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n706), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n765), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n769), .A2(new_n770), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G330), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n750), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n741), .B1(new_n781), .B2(G1), .ZN(G364));
  NOR2_X1   g0582(.A1(new_n355), .A2(new_n222), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n270), .B1(new_n783), .B2(G45), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n737), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n224), .A2(G355), .A3(new_n290), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n735), .A2(new_n290), .ZN(new_n789));
  INV_X1    g0589(.A(new_n232), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n789), .B1(new_n790), .B2(G45), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n249), .A2(new_n272), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n788), .B1(G116), .B2(new_n224), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n230), .B1(G20), .B2(new_n332), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n787), .B1(new_n793), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT94), .Z(new_n800));
  NAND2_X1  g0600(.A1(new_n710), .A2(new_n713), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n796), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n229), .A2(new_n326), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n460), .A2(G200), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G190), .A2(G200), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n202), .A2(new_n807), .B1(new_n809), .B2(new_n317), .ZN(new_n810));
  NOR2_X1   g0610(.A1(G179), .A2(G200), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n355), .A2(new_n460), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G159), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT32), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n805), .A2(G200), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n460), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n810), .B(new_n815), .C1(G50), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n806), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n355), .B1(new_n819), .B2(G179), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT97), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n520), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT96), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n816), .B2(G190), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n805), .A2(KEYINPUT96), .A3(new_n460), .A4(G200), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G68), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n370), .A2(G179), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n833), .A2(G20), .A3(G190), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(G87), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n355), .A2(new_n460), .A3(new_n833), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n836), .B(new_n290), .C1(new_n339), .C2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT95), .Z(new_n839));
  NAND4_X1  g0639(.A1(new_n818), .A2(new_n827), .A3(new_n832), .A4(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n824), .A2(G294), .B1(G326), .B2(new_n817), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT98), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(G322), .ZN(new_n844));
  INV_X1    g0644(.A(G283), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n807), .A2(new_n844), .B1(new_n845), .B2(new_n837), .ZN(new_n846));
  INV_X1    g0646(.A(G303), .ZN(new_n847));
  INV_X1    g0647(.A(G311), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n259), .B1(new_n847), .B2(new_n834), .C1(new_n809), .C2(new_n848), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n846), .B(new_n849), .C1(G329), .C2(new_n813), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n841), .A2(new_n842), .ZN(new_n851));
  XNOR2_X1  g0651(.A(KEYINPUT33), .B(G317), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n831), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n843), .A2(new_n850), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n840), .A2(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n800), .B(new_n804), .C1(new_n797), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n802), .A2(G330), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n710), .A2(G330), .A3(new_n713), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n859), .A2(new_n786), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n856), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(G396));
  NOR2_X1   g0662(.A1(new_n369), .A2(new_n706), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n367), .A2(new_n706), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n374), .B2(new_n371), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n863), .B1(new_n369), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n749), .B(new_n866), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n867), .A2(new_n779), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n786), .B1(new_n867), .B2(new_n779), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n797), .A2(new_n794), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT99), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n786), .B1(new_n872), .B2(G77), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n290), .B1(new_n835), .B2(G107), .ZN(new_n874));
  INV_X1    g0674(.A(new_n817), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n874), .B1(new_n600), .B2(new_n809), .C1(new_n875), .C2(new_n847), .ZN(new_n876));
  INV_X1    g0676(.A(new_n807), .ZN(new_n877));
  INV_X1    g0677(.A(new_n837), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n877), .A2(G294), .B1(new_n878), .B2(G87), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n848), .B2(new_n812), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n876), .A2(new_n826), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n831), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n881), .B1(new_n845), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n809), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n884), .A2(G159), .B1(new_n877), .B2(G143), .ZN(new_n885));
  INV_X1    g0685(.A(G137), .ZN(new_n886));
  INV_X1    g0686(.A(G150), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n885), .B1(new_n886), .B2(new_n875), .C1(new_n882), .C2(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT34), .Z(new_n889));
  NAND2_X1  g0689(.A1(new_n878), .A2(G68), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n290), .B1(new_n834), .B2(new_n207), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n813), .B2(G132), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n890), .B(new_n892), .C1(new_n825), .C2(new_n202), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n883), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n873), .B1(new_n894), .B2(new_n797), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n795), .B2(new_n866), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT100), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n870), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(G384));
  NOR2_X1   g0699(.A1(new_n783), .A2(new_n270), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  OAI221_X1 g0701(.A(G68), .B1(new_n436), .B2(new_n290), .C1(new_n422), .C2(new_n434), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT16), .B1(new_n902), .B2(new_n432), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n417), .B1(new_n439), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n704), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n479), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n474), .A2(new_n307), .A3(new_n438), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n909), .B(new_n417), .C1(new_n461), .C2(new_n462), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n456), .A2(new_n904), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n911), .A3(new_n906), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT102), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT37), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n440), .A2(new_n905), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT37), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n457), .A2(new_n915), .A3(new_n910), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n913), .B1(new_n912), .B2(KEYINPUT37), .ZN(new_n919));
  OAI211_X1 g0719(.A(KEYINPUT38), .B(new_n908), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n479), .A2(new_n440), .A3(new_n905), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n457), .A2(new_n915), .A3(new_n910), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT37), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n917), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT38), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n901), .B1(new_n921), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n284), .A2(new_n327), .A3(new_n297), .ZN(new_n928));
  OAI21_X1  g0728(.A(G169), .B1(new_n322), .B2(new_n323), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n331), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n329), .A2(KEYINPUT14), .A3(G169), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n932), .A2(new_n321), .A3(new_n706), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n908), .B1(new_n918), .B2(new_n919), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT38), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(KEYINPUT39), .A3(new_n920), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n927), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n695), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n537), .A2(new_n653), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT26), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n745), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n653), .B1(new_n539), .B2(new_n541), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n942), .B1(new_n943), .B2(new_n941), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n764), .B(new_n866), .C1(new_n939), .C2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n863), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n335), .A2(new_n706), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n932), .B2(new_n663), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n663), .B(new_n948), .C1(new_n932), .C2(new_n321), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT101), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT101), .B1(new_n336), .B2(new_n948), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n936), .A2(new_n920), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n947), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n704), .B1(new_n659), .B2(new_n660), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n938), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT103), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT103), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n938), .A2(new_n957), .A3(new_n961), .A4(new_n958), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n674), .B1(new_n750), .B2(new_n675), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n963), .B(new_n964), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n771), .A2(new_n772), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT93), .B1(new_n774), .B2(KEYINPUT30), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n966), .A2(new_n967), .A3(new_n760), .A4(new_n762), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n770), .A2(new_n777), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n970), .A2(new_n866), .A3(new_n955), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n906), .B1(new_n667), .B2(new_n661), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n914), .A2(new_n917), .ZN(new_n973));
  INV_X1    g0773(.A(new_n919), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n926), .B1(new_n975), .B2(KEYINPUT38), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT40), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT40), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n865), .A2(new_n369), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n946), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n951), .A2(new_n952), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n336), .A2(KEYINPUT101), .A3(new_n948), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n980), .B1(new_n983), .B2(new_n950), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n956), .A2(new_n978), .A3(new_n970), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n977), .A2(new_n985), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n480), .A2(new_n970), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n986), .A2(new_n987), .ZN(new_n990));
  INV_X1    g0790(.A(G330), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n900), .B1(new_n965), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n993), .B2(new_n965), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT35), .ZN(new_n996));
  OAI211_X1 g0796(.A(G116), .B(new_n231), .C1(new_n523), .C2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n996), .B2(new_n523), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT36), .Z(new_n999));
  NAND2_X1  g0799(.A1(new_n430), .A2(G77), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n245), .B1(new_n790), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1001), .A2(G1), .A3(new_n222), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n995), .A2(new_n999), .A3(new_n1002), .ZN(G367));
  INV_X1    g0803(.A(new_n797), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n290), .B1(new_n202), .B2(new_n834), .C1(new_n809), .C2(new_n207), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G143), .B2(new_n817), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n807), .A2(new_n887), .B1(new_n886), .B2(new_n812), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G77), .B2(new_n878), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n203), .B2(new_n825), .C1(new_n428), .C2(new_n882), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n807), .A2(new_n847), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n834), .A2(new_n600), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT46), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1011), .B(new_n1013), .C1(G283), .C2(new_n884), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n339), .B2(new_n825), .C1(new_n848), .C2(new_n875), .ZN(new_n1015));
  INV_X1    g0815(.A(G317), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n259), .B1(new_n812), .B2(new_n1016), .C1(new_n520), .C2(new_n837), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1017), .A2(KEYINPUT110), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(KEYINPUT110), .ZN(new_n1019));
  INV_X1    g0819(.A(G294), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1018), .B(new_n1019), .C1(new_n1020), .C2(new_n882), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1010), .B1(new_n1015), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT47), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1004), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n1023), .B2(new_n1022), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n789), .A2(new_n240), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n798), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n735), .B2(new_n358), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n787), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n652), .A2(new_n706), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n654), .A2(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n679), .A2(new_n1030), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1025), .B(new_n1029), .C1(new_n803), .C2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n1035));
  INV_X1    g0835(.A(KEYINPUT107), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n728), .A2(new_n536), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n539), .A2(new_n541), .A3(new_n547), .A4(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n540), .A2(new_n728), .A3(new_n511), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n731), .A2(new_n1036), .A3(new_n1040), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n718), .A2(new_n712), .A3(new_n719), .A4(new_n720), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n729), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(KEYINPUT107), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1035), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1036), .B1(new_n731), .B2(new_n1040), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1042), .A2(new_n1045), .A3(KEYINPUT107), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1035), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT45), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n731), .A2(KEYINPUT45), .A3(new_n1040), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1047), .A2(new_n1051), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n725), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n730), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n721), .A2(new_n722), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n1043), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n859), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n714), .A2(new_n1043), .A3(new_n1059), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n1063), .A2(new_n750), .A3(new_n779), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1047), .A2(new_n726), .A3(new_n1051), .A4(new_n1055), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1057), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT108), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT108), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1057), .A2(new_n1068), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n780), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n737), .B(KEYINPUT41), .Z(new_n1071));
  OAI21_X1  g0871(.A(new_n784), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1033), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT43), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1033), .A2(KEYINPUT43), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n689), .B1(new_n1042), .B2(new_n718), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n764), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1040), .A2(new_n597), .A3(new_n730), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(KEYINPUT42), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT104), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT105), .ZN(new_n1085));
  OR3_X1    g0885(.A1(new_n1079), .A2(new_n1085), .A3(KEYINPUT42), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1085), .B1(new_n1079), .B2(KEYINPUT42), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1075), .B(new_n1076), .C1(new_n1084), .C2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1081), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1090), .B1(new_n1091), .B2(KEYINPUT104), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1092), .A2(new_n1074), .A3(new_n1073), .A4(new_n1083), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n726), .A2(new_n1042), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1089), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1094), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1072), .A2(KEYINPUT109), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT109), .B1(new_n1072), .B2(new_n1097), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1034), .B1(new_n1098), .B2(new_n1099), .ZN(G387));
  NAND2_X1  g0900(.A1(new_n1063), .A2(new_n785), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(KEYINPUT111), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT111), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1063), .A2(new_n1103), .A3(new_n785), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n724), .A2(new_n796), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n789), .B1(new_n237), .B2(new_n272), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n224), .A2(new_n290), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n734), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n272), .B1(new_n203), .B2(new_n317), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n361), .A2(G50), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(KEYINPUT50), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1111), .B(new_n734), .C1(KEYINPUT50), .C2(new_n1110), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1108), .A2(new_n1112), .B1(new_n339), .B2(new_n735), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n786), .B1(new_n1113), .B2(new_n1027), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n825), .A2(new_n357), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n831), .A2(new_n389), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n809), .A2(new_n203), .B1(new_n887), .B2(new_n812), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G50), .B2(new_n877), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n290), .B1(new_n317), .B2(new_n834), .C1(new_n837), .C2(new_n520), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G159), .B2(new_n817), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1116), .A2(new_n1117), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n290), .B1(new_n813), .B2(G326), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n825), .A2(new_n845), .B1(new_n1020), .B2(new_n834), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n884), .A2(G303), .B1(new_n877), .B2(G317), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1125), .B1(new_n844), .B2(new_n875), .C1(new_n882), .C2(new_n848), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT48), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n1127), .B2(new_n1126), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT49), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1123), .B1(new_n600), .B2(new_n837), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1122), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1114), .B1(new_n1133), .B2(new_n797), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1102), .A2(new_n1104), .B1(new_n1105), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1064), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n737), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n781), .A2(new_n1063), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(G393));
  NAND2_X1  g0939(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1057), .A2(new_n1065), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n1136), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n737), .A3(new_n1142), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1141), .A2(KEYINPUT112), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n784), .B1(new_n1141), .B2(KEYINPUT112), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1042), .A2(new_n796), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n789), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n798), .B1(new_n520), .B2(new_n224), .C1(new_n1147), .C2(new_n244), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n786), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n290), .B1(new_n203), .B2(new_n834), .C1(new_n837), .C2(new_n571), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n361), .A2(new_n809), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(G143), .C2(new_n813), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n824), .A2(G77), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1152), .B(new_n1153), .C1(new_n207), .C2(new_n882), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n817), .A2(G150), .B1(new_n877), .B2(G159), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT51), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n259), .B1(new_n845), .B2(new_n834), .C1(new_n837), .C2(new_n339), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n809), .A2(new_n1020), .B1(new_n844), .B2(new_n812), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(G116), .C2(new_n824), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n847), .B2(new_n882), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n817), .A2(G317), .B1(new_n877), .B2(G311), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT52), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n1154), .A2(new_n1156), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1149), .B1(new_n1163), .B2(new_n797), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1144), .A2(new_n1145), .B1(new_n1146), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1143), .A2(new_n1165), .ZN(G390));
  AND2_X1   g0966(.A1(new_n970), .A2(G330), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n480), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1168), .B(new_n674), .C1(new_n675), .C2(new_n750), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT31), .B1(new_n968), .B2(new_n706), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1170), .A2(new_n767), .A3(new_n768), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n991), .B1(new_n1171), .B2(new_n770), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n955), .B1(new_n1172), .B2(new_n866), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n970), .A2(G330), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n949), .B1(new_n981), .B2(new_n982), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1174), .A2(new_n980), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n947), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1175), .B1(new_n1174), .B2(new_n980), .ZN(new_n1178));
  OAI21_X1  g0978(.A(KEYINPUT26), .B1(new_n537), .B2(new_n653), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n679), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n941), .B2(new_n943), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n718), .A2(new_n623), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n548), .A2(new_n694), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n706), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n863), .B1(new_n1184), .B2(new_n979), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n778), .A2(G330), .A3(new_n866), .A4(new_n955), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1178), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1169), .B1(new_n1177), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1186), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n933), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n863), .B1(new_n749), .B2(new_n866), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1191), .B1(new_n1192), .B2(new_n1175), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n927), .A2(new_n937), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT113), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n720), .B(new_n979), .C1(new_n744), .C2(new_n747), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1175), .B1(new_n1196), .B2(new_n946), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n924), .A2(new_n917), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n915), .B1(new_n667), .B2(new_n661), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n935), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n920), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1191), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1195), .B1(new_n1197), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n933), .B1(new_n1200), .B2(new_n920), .ZN(new_n1204));
  OAI211_X1 g1004(.A(KEYINPUT113), .B(new_n1204), .C1(new_n1185), .C2(new_n1175), .ZN(new_n1205));
  AOI221_X4 g1005(.A(new_n1190), .B1(new_n1193), .B2(new_n1194), .C1(new_n1203), .C2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1167), .A2(new_n984), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1205), .A2(new_n1203), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1207), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1189), .B1(new_n1206), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1186), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1188), .B(new_n1212), .C1(new_n1213), .C2(new_n1207), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1211), .A2(new_n1214), .A3(new_n737), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1206), .A2(new_n1210), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1194), .A2(new_n794), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n786), .B1(new_n872), .B2(new_n389), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT114), .Z(new_n1219));
  NOR2_X1   g1019(.A1(new_n834), .A2(new_n887), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT53), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n813), .A2(G125), .ZN(new_n1222));
  INV_X1    g1022(.A(G132), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1221), .B(new_n1222), .C1(new_n1223), .C2(new_n807), .ZN(new_n1224));
  INV_X1    g1024(.A(G128), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n290), .B1(new_n207), .B2(new_n837), .C1(new_n875), .C2(new_n1225), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G159), .C2(new_n824), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(KEYINPUT54), .B(G143), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n831), .A2(G137), .B1(new_n884), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1231), .A2(KEYINPUT115), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(KEYINPUT115), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1227), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1234), .A2(KEYINPUT116), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n875), .A2(new_n845), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n884), .A2(G97), .B1(G294), .B2(new_n813), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1237), .A2(new_n259), .A3(new_n836), .A4(new_n890), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1236), .B(new_n1238), .C1(G107), .C2(new_n831), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1153), .B1(new_n600), .B2(new_n807), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT117), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1234), .A2(KEYINPUT116), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1235), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1219), .B1(new_n1244), .B2(new_n797), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1216), .A2(new_n785), .B1(new_n1217), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1215), .A2(new_n1246), .ZN(G378));
  NOR3_X1   g1047(.A1(new_n797), .A2(G50), .A3(new_n794), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n736), .A2(new_n290), .ZN(new_n1249));
  AOI211_X1 g1049(.A(G50), .B(new_n1249), .C1(new_n255), .C2(new_n271), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n837), .A2(new_n202), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT118), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G68), .B2(new_n824), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n807), .A2(new_n339), .B1(new_n845), .B2(new_n812), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1249), .B1(new_n317), .B2(new_n834), .C1(new_n809), .C2(new_n357), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1255), .B(new_n1256), .C1(G116), .C2(new_n817), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1254), .B(new_n1257), .C1(new_n520), .C2(new_n882), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT58), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1250), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n835), .A2(new_n1229), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(KEYINPUT119), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n1262), .B1(new_n1225), .B2(new_n807), .C1(new_n886), .C2(new_n809), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(G125), .B2(new_n817), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1264), .B1(new_n1223), .B2(new_n882), .C1(new_n887), .C2(new_n825), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT59), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n255), .B(new_n271), .C1(new_n837), .C2(new_n428), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(G124), .B2(new_n813), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1265), .A2(KEYINPUT59), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1260), .B1(new_n1259), .B2(new_n1258), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n787), .B(new_n1248), .C1(new_n1271), .C2(new_n797), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n396), .A2(new_n704), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n413), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n398), .B1(new_n671), .B2(new_n672), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1273), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1274), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1278), .B1(new_n1274), .B2(new_n1277), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n794), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1272), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT120), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n984), .A2(new_n978), .A3(new_n970), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1201), .A2(new_n984), .A3(new_n970), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1286), .A2(new_n956), .B1(new_n1287), .B2(KEYINPUT40), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1281), .B1(new_n1288), .B2(new_n991), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1281), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n986), .A2(G330), .A3(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1289), .A2(new_n960), .A3(new_n1291), .A4(new_n962), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1289), .A2(new_n1291), .B1(new_n960), .B2(new_n962), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1285), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n959), .A2(KEYINPUT103), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n962), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1290), .B1(new_n986), .B2(G330), .ZN(new_n1298));
  AOI211_X1 g1098(.A(new_n991), .B(new_n1281), .C1(new_n977), .C2(new_n985), .ZN(new_n1299));
  OAI22_X1  g1099(.A1(new_n1296), .A2(new_n1297), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(KEYINPUT120), .A3(new_n1292), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1295), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1284), .B1(new_n1302), .B2(new_n785), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1169), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1214), .A2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT57), .B1(new_n1302), .B2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1169), .B1(new_n1216), .B2(new_n1188), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1300), .A2(KEYINPUT57), .A3(new_n1292), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n737), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1303), .B1(new_n1306), .B2(new_n1309), .ZN(G375));
  INV_X1    g1110(.A(new_n1187), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1175), .B1(new_n779), .B2(new_n980), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1192), .B1(new_n1312), .B2(new_n1207), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n785), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n786), .B1(new_n872), .B2(G68), .ZN(new_n1315));
  OAI22_X1  g1115(.A1(new_n875), .A2(new_n1223), .B1(new_n886), .B2(new_n807), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1316), .B1(new_n831), .B2(new_n1229), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1317), .B(KEYINPUT121), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n259), .B1(new_n835), .B2(G159), .ZN(new_n1319));
  OAI221_X1 g1119(.A(new_n1319), .B1(new_n1225), .B2(new_n812), .C1(new_n809), .C2(new_n887), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1321), .B(new_n1252), .C1(new_n207), .C2(new_n825), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n882), .A2(new_n600), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n290), .B1(new_n835), .B2(G97), .ZN(new_n1324));
  OAI221_X1 g1124(.A(new_n1324), .B1(new_n317), .B2(new_n837), .C1(new_n875), .C2(new_n1020), .ZN(new_n1325));
  AOI22_X1  g1125(.A1(new_n884), .A2(G107), .B1(new_n877), .B2(G283), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1326), .B1(new_n847), .B2(new_n812), .ZN(new_n1327));
  OR3_X1    g1127(.A1(new_n1325), .A2(new_n1327), .A3(new_n1115), .ZN(new_n1328));
  OAI22_X1  g1128(.A1(new_n1318), .A2(new_n1322), .B1(new_n1323), .B2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1315), .B1(new_n1329), .B2(new_n797), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1330), .B1(new_n795), .B2(new_n955), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1314), .A2(new_n1331), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1188), .A2(new_n1071), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1177), .A2(new_n1169), .A3(new_n1187), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1332), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(G381));
  INV_X1    g1136(.A(KEYINPUT122), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1099), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1072), .A2(KEYINPUT109), .A3(new_n1097), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  NOR3_X1   g1140(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1335), .ZN(new_n1342));
  NOR3_X1   g1142(.A1(G378), .A2(new_n1342), .A3(G390), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1340), .A2(new_n1343), .A3(new_n1034), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(G375), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1337), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1347));
  NOR3_X1   g1147(.A1(new_n1344), .A2(G375), .A3(KEYINPUT122), .ZN(new_n1348));
  OR2_X1    g1148(.A1(new_n1347), .A2(new_n1348), .ZN(G407));
  INV_X1    g1149(.A(G213), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n705), .A2(G213), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(new_n1351), .B(KEYINPUT123), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1352), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(G378), .A2(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1350), .B1(new_n1346), .B2(new_n1354), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1355), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT124), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  OAI211_X1 g1158(.A(KEYINPUT124), .B(new_n1355), .C1(new_n1347), .C2(new_n1348), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1358), .A2(new_n1359), .ZN(G409));
  AND3_X1   g1160(.A1(new_n1300), .A2(KEYINPUT120), .A3(new_n1292), .ZN(new_n1361));
  AOI21_X1  g1161(.A(KEYINPUT120), .B1(new_n1300), .B2(new_n1292), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1305), .B1(new_n1361), .B2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT57), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1309), .B1(new_n1363), .B2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(G378), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n785), .B1(new_n1361), .B2(new_n1362), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1367), .A2(new_n1283), .ZN(new_n1368));
  NOR3_X1   g1168(.A1(new_n1365), .A2(new_n1366), .A3(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1071), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1302), .A2(new_n1370), .A3(new_n1305), .ZN(new_n1371));
  NOR2_X1   g1171(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1284), .B1(new_n1372), .B2(new_n785), .ZN(new_n1373));
  AOI21_X1  g1173(.A(G378), .B1(new_n1371), .B2(new_n1373), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1353), .B1(new_n1369), .B2(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1352), .A2(G2897), .ZN(new_n1376));
  INV_X1    g1176(.A(new_n1376), .ZN(new_n1377));
  NAND4_X1  g1177(.A1(new_n1177), .A2(new_n1169), .A3(KEYINPUT60), .A4(new_n1187), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1378), .A2(new_n737), .ZN(new_n1379));
  INV_X1    g1179(.A(new_n1379), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT60), .ZN(new_n1381));
  OAI21_X1  g1181(.A(new_n1334), .B1(new_n1188), .B2(new_n1381), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1380), .A2(new_n1382), .ZN(new_n1383));
  INV_X1    g1183(.A(new_n1332), .ZN(new_n1384));
  AOI21_X1  g1184(.A(G384), .B1(new_n1383), .B2(new_n1384), .ZN(new_n1385));
  AOI211_X1 g1185(.A(new_n898), .B(new_n1332), .C1(new_n1380), .C2(new_n1382), .ZN(new_n1386));
  NOR2_X1   g1186(.A1(new_n1385), .A2(new_n1386), .ZN(new_n1387));
  INV_X1    g1187(.A(KEYINPUT125), .ZN(new_n1388));
  AOI21_X1  g1188(.A(new_n1377), .B1(new_n1387), .B2(new_n1388), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1383), .A2(new_n1384), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1390), .A2(new_n898), .ZN(new_n1391));
  NAND3_X1  g1191(.A1(new_n1383), .A2(G384), .A3(new_n1384), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1391), .A2(new_n1392), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1393), .A2(KEYINPUT125), .ZN(new_n1394));
  NAND2_X1  g1194(.A1(new_n1389), .A2(new_n1394), .ZN(new_n1395));
  NOR4_X1   g1195(.A1(new_n1385), .A2(new_n1386), .A3(KEYINPUT125), .A4(new_n1376), .ZN(new_n1396));
  INV_X1    g1196(.A(new_n1396), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1395), .A2(new_n1397), .ZN(new_n1398));
  AOI21_X1  g1198(.A(KEYINPUT61), .B1(new_n1375), .B2(new_n1398), .ZN(new_n1399));
  OAI211_X1 g1199(.A(new_n1353), .B(new_n1387), .C1(new_n1369), .C2(new_n1374), .ZN(new_n1400));
  INV_X1    g1200(.A(KEYINPUT63), .ZN(new_n1401));
  NAND2_X1  g1201(.A1(new_n1400), .A2(new_n1401), .ZN(new_n1402));
  INV_X1    g1202(.A(G390), .ZN(new_n1403));
  NAND2_X1  g1203(.A1(G387), .A2(new_n1403), .ZN(new_n1404));
  XNOR2_X1  g1204(.A(G393), .B(new_n861), .ZN(new_n1405));
  OAI211_X1 g1205(.A(new_n1034), .B(G390), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1406));
  AND3_X1   g1206(.A1(new_n1404), .A2(new_n1405), .A3(new_n1406), .ZN(new_n1407));
  AOI21_X1  g1207(.A(new_n1405), .B1(new_n1404), .B2(new_n1406), .ZN(new_n1408));
  NOR2_X1   g1208(.A1(new_n1407), .A2(new_n1408), .ZN(new_n1409));
  OAI211_X1 g1209(.A(G378), .B(new_n1303), .C1(new_n1306), .C2(new_n1309), .ZN(new_n1410));
  OAI21_X1  g1210(.A(new_n1373), .B1(new_n1363), .B2(new_n1071), .ZN(new_n1411));
  NAND2_X1  g1211(.A1(new_n1411), .A2(new_n1366), .ZN(new_n1412));
  AOI21_X1  g1212(.A(new_n1352), .B1(new_n1410), .B2(new_n1412), .ZN(new_n1413));
  NAND3_X1  g1213(.A1(new_n1413), .A2(KEYINPUT63), .A3(new_n1387), .ZN(new_n1414));
  NAND4_X1  g1214(.A1(new_n1399), .A2(new_n1402), .A3(new_n1409), .A4(new_n1414), .ZN(new_n1415));
  INV_X1    g1215(.A(KEYINPUT61), .ZN(new_n1416));
  AOI21_X1  g1216(.A(new_n1396), .B1(new_n1389), .B2(new_n1394), .ZN(new_n1417));
  OAI21_X1  g1217(.A(new_n1416), .B1(new_n1413), .B2(new_n1417), .ZN(new_n1418));
  INV_X1    g1218(.A(KEYINPUT62), .ZN(new_n1419));
  NAND2_X1  g1219(.A1(new_n1400), .A2(new_n1419), .ZN(new_n1420));
  NAND3_X1  g1220(.A1(new_n1413), .A2(KEYINPUT62), .A3(new_n1387), .ZN(new_n1421));
  AOI21_X1  g1221(.A(new_n1418), .B1(new_n1420), .B2(new_n1421), .ZN(new_n1422));
  INV_X1    g1222(.A(KEYINPUT126), .ZN(new_n1423));
  OAI21_X1  g1223(.A(new_n1423), .B1(new_n1407), .B2(new_n1408), .ZN(new_n1424));
  NAND2_X1  g1224(.A1(new_n1404), .A2(new_n1406), .ZN(new_n1425));
  INV_X1    g1225(.A(new_n1405), .ZN(new_n1426));
  NAND2_X1  g1226(.A1(new_n1425), .A2(new_n1426), .ZN(new_n1427));
  NAND3_X1  g1227(.A1(new_n1404), .A2(new_n1405), .A3(new_n1406), .ZN(new_n1428));
  NAND3_X1  g1228(.A1(new_n1427), .A2(KEYINPUT126), .A3(new_n1428), .ZN(new_n1429));
  NAND2_X1  g1229(.A1(new_n1424), .A2(new_n1429), .ZN(new_n1430));
  OAI21_X1  g1230(.A(new_n1415), .B1(new_n1422), .B2(new_n1430), .ZN(G405));
  OAI21_X1  g1231(.A(KEYINPUT127), .B1(new_n1407), .B2(new_n1408), .ZN(new_n1432));
  INV_X1    g1232(.A(KEYINPUT127), .ZN(new_n1433));
  NAND3_X1  g1233(.A1(new_n1427), .A2(new_n1433), .A3(new_n1428), .ZN(new_n1434));
  OAI21_X1  g1234(.A(new_n1366), .B1(new_n1365), .B2(new_n1368), .ZN(new_n1435));
  AND3_X1   g1235(.A1(new_n1435), .A2(new_n1393), .A3(new_n1410), .ZN(new_n1436));
  AOI21_X1  g1236(.A(new_n1393), .B1(new_n1435), .B2(new_n1410), .ZN(new_n1437));
  NOR2_X1   g1237(.A1(new_n1436), .A2(new_n1437), .ZN(new_n1438));
  NAND3_X1  g1238(.A1(new_n1432), .A2(new_n1434), .A3(new_n1438), .ZN(new_n1439));
  OAI221_X1 g1239(.A(KEYINPUT127), .B1(new_n1407), .B2(new_n1408), .C1(new_n1437), .C2(new_n1436), .ZN(new_n1440));
  NAND2_X1  g1240(.A1(new_n1439), .A2(new_n1440), .ZN(G402));
endmodule


