//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1050,
    new_n1051, new_n1052;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G43gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n204), .B2(KEYINPUT85), .ZN(new_n205));
  OR2_X1    g004(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n207));
  AOI21_X1  g006(.A(G36gat), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G29gat), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n209), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n205), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n208), .A2(new_n210), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n211), .A2(new_n213), .B1(new_n214), .B2(new_n202), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT17), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n205), .B(new_n212), .C1(new_n208), .C2(new_n210), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT86), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n215), .A2(KEYINPUT86), .A3(new_n216), .A4(new_n217), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n215), .A2(new_n217), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  INV_X1    g023(.A(G1gat), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(KEYINPUT16), .A3(new_n225), .ZN(new_n227));
  OR2_X1    g026(.A1(KEYINPUT87), .A2(G8gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(KEYINPUT87), .A3(G8gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT87), .A2(G8gat), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n226), .A2(new_n227), .A3(new_n231), .A4(new_n228), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n223), .A2(KEYINPUT17), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n222), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(new_n232), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(new_n223), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n234), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n234), .A2(KEYINPUT18), .A3(new_n235), .A4(new_n238), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n235), .B(KEYINPUT13), .Z(new_n243));
  AND2_X1   g042(.A1(new_n236), .A2(new_n223), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n243), .B1(new_n244), .B2(new_n237), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n241), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT84), .ZN(new_n248));
  XOR2_X1   g047(.A(G113gat), .B(G141gat), .Z(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(G169gat), .B(G197gat), .Z(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT12), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n246), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n253), .A2(new_n242), .A3(new_n245), .A4(new_n241), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT88), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n255), .A2(KEYINPUT88), .A3(new_n256), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G1gat), .B(G29gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT0), .ZN(new_n264));
  XNOR2_X1  g063(.A(G57gat), .B(G85gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n264), .B(new_n265), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  OR2_X1    g066(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(G134gat), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n268), .A2(KEYINPUT69), .A3(G134gat), .A4(new_n269), .ZN(new_n273));
  INV_X1    g072(.A(G134gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G127gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n272), .A2(new_n273), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G120gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G113gat), .ZN(new_n282));
  INV_X1    g081(.A(G113gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G120gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT1), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT70), .B1(new_n281), .B2(G113gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n281), .A2(G113gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n281), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT1), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G127gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G134gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n275), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n275), .A2(new_n295), .A3(KEYINPUT71), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G141gat), .ZN(new_n302));
  INV_X1    g101(.A(G148gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G162gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G155gat), .ZN(new_n306));
  INV_X1    g105(.A(G155gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G162gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n304), .A2(new_n306), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n313));
  OAI21_X1  g112(.A(G155gat), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT2), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n306), .A2(new_n308), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n304), .A2(new_n317), .A3(new_n309), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n311), .A2(new_n315), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n288), .A2(new_n301), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT4), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n280), .A2(new_n287), .B1(new_n293), .B2(new_n300), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n316), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT77), .B(G162gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n317), .B1(new_n324), .B2(G155gat), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n323), .B1(new_n325), .B2(new_n310), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT78), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT78), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n329), .B(new_n323), .C1(new_n325), .C2(new_n310), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n322), .A2(new_n327), .A3(new_n328), .A4(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT79), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n321), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n332), .B1(new_n321), .B2(new_n331), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n326), .A2(KEYINPUT3), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n336), .B(new_n323), .C1(new_n325), .C2(new_n310), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n275), .A2(new_n295), .A3(KEYINPUT71), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT71), .B1(new_n275), .B2(new_n295), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT70), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(new_n283), .B2(G120gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(new_n292), .A3(new_n284), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n286), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n270), .A2(new_n271), .B1(new_n277), .B2(new_n278), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n346), .A2(new_n273), .B1(new_n286), .B2(new_n285), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n335), .B(new_n337), .C1(new_n345), .C2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT5), .ZN(new_n349));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n333), .A2(new_n334), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n326), .B1(new_n347), .B2(new_n345), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n320), .ZN(new_n354));
  INV_X1    g153(.A(new_n350), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n349), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n320), .A2(new_n328), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n322), .A2(new_n327), .A3(KEYINPUT4), .A4(new_n330), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n357), .A2(new_n358), .A3(new_n348), .A4(new_n350), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n267), .B1(new_n352), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n356), .A2(new_n359), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n321), .A2(new_n331), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT79), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n321), .A2(new_n331), .A3(new_n332), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n363), .B(new_n266), .C1(new_n367), .C2(new_n351), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n361), .A2(new_n362), .A3(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(KEYINPUT6), .B(new_n267), .C1(new_n352), .C2(new_n360), .ZN(new_n370));
  NAND2_X1  g169(.A1(G211gat), .A2(G218gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT22), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT74), .ZN(new_n374));
  OR2_X1    g173(.A1(G197gat), .A2(G204gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(G197gat), .A2(G204gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT74), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n374), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G211gat), .B(G218gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n375), .A2(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n385), .A2(new_n382), .A3(new_n374), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388));
  INV_X1    g187(.A(G169gat), .ZN(new_n389));
  INV_X1    g188(.A(G176gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT23), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(G169gat), .B2(G176gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NOR3_X1   g196(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G183gat), .A2(G190gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT24), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT24), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(G183gat), .A3(G190gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n395), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(G183gat), .A2(G190gat), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n408), .B1(new_n401), .B2(new_n403), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n391), .A2(new_n393), .A3(KEYINPUT25), .A4(new_n394), .ZN(new_n410));
  OAI22_X1  g209(.A1(new_n405), .A2(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(G169gat), .A2(G176gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT26), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT26), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n394), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n413), .B(new_n400), .C1(new_n415), .C2(new_n412), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G183gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT27), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT27), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G183gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT66), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(G190gat), .B1(new_n419), .B2(KEYINPUT66), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT28), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT28), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n422), .A2(new_n427), .A3(G190gat), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n417), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n388), .B1(new_n411), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n411), .A2(new_n429), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT29), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n430), .B1(new_n433), .B2(new_n388), .ZN(new_n434));
  INV_X1    g233(.A(new_n388), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT76), .B(KEYINPUT29), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n411), .B2(new_n429), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n436), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT75), .ZN(new_n441));
  AND4_X1   g240(.A1(new_n382), .A2(new_n374), .A3(new_n377), .A4(new_n380), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n382), .B1(new_n385), .B2(new_n374), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n384), .A2(KEYINPUT75), .A3(new_n386), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n387), .A2(new_n434), .B1(new_n440), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT30), .ZN(new_n449));
  XNOR2_X1  g248(.A(G8gat), .B(G36gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(G64gat), .B(G92gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n450), .B(new_n451), .Z(new_n452));
  NAND3_X1  g251(.A1(new_n448), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n452), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT29), .B1(new_n411), .B2(new_n429), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n436), .B(new_n387), .C1(new_n435), .C2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n410), .A2(new_n409), .ZN(new_n458));
  INV_X1    g257(.A(new_n398), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n404), .A2(new_n459), .A3(new_n396), .ZN(new_n460));
  INV_X1    g259(.A(new_n395), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n458), .B1(new_n462), .B2(new_n406), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n419), .A2(KEYINPUT66), .ZN(new_n464));
  INV_X1    g263(.A(G190gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT66), .B1(new_n419), .B2(new_n421), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n427), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n422), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(KEYINPUT28), .A3(new_n465), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n416), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n463), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n388), .B1(new_n472), .B2(new_n438), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n446), .B1(new_n473), .B2(new_n436), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n454), .B1(new_n457), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n440), .A2(new_n447), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(new_n456), .A3(new_n452), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(KEYINPUT30), .A3(new_n477), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n369), .A2(new_n370), .B1(new_n453), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT35), .ZN(new_n480));
  NAND2_X1  g279(.A1(G228gat), .A2(G233gat), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n432), .B1(new_n442), .B2(new_n443), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n336), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n483), .B2(new_n326), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n337), .A2(new_n437), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(new_n444), .A3(new_n445), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT80), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n485), .A2(new_n444), .A3(KEYINPUT80), .A4(new_n445), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n484), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G22gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n387), .A2(new_n437), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n492), .A2(new_n336), .B1(new_n327), .B2(new_n330), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n387), .B1(new_n337), .B2(new_n437), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n481), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n490), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT81), .ZN(new_n497));
  XNOR2_X1  g296(.A(G78gat), .B(G106gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(KEYINPUT31), .B(G50gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n490), .A2(new_n495), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G22gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n496), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT81), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n503), .A2(new_n506), .A3(new_n496), .A4(new_n500), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n411), .B(new_n429), .C1(new_n345), .C2(new_n347), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n322), .B1(new_n463), .B2(new_n471), .ZN(new_n510));
  INV_X1    g309(.A(G227gat), .ZN(new_n511));
  INV_X1    g310(.A(G233gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(G71gat), .B(G99gat), .Z(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G43gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT33), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(KEYINPUT72), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n514), .A2(KEYINPUT32), .A3(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n509), .A2(new_n510), .A3(new_n513), .A4(new_n517), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT72), .B1(new_n521), .B2(new_n518), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n514), .A2(KEYINPUT32), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n510), .ZN(new_n525));
  INV_X1    g324(.A(new_n513), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT34), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT34), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n529), .A3(new_n526), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n524), .B(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n479), .A2(new_n480), .A3(new_n508), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n369), .A2(new_n370), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT73), .B1(new_n528), .B2(new_n530), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n524), .B(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n478), .A2(new_n453), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n508), .A2(new_n534), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n538), .A2(KEYINPUT82), .A3(KEYINPUT35), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT82), .B1(new_n538), .B2(KEYINPUT35), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n533), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n532), .A2(KEYINPUT36), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n536), .A2(KEYINPUT36), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n478), .A2(new_n361), .A3(new_n453), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT40), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n365), .A2(new_n366), .A3(new_n348), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT39), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n548), .A3(new_n355), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n266), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT39), .B1(new_n354), .B2(new_n355), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(new_n547), .B2(new_n355), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n546), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n552), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n554), .A2(KEYINPUT40), .A3(new_n266), .A4(new_n549), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n545), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT37), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n452), .B1(new_n448), .B2(new_n557), .ZN(new_n558));
  OAI22_X1  g357(.A1(new_n434), .A2(new_n387), .B1(new_n440), .B2(new_n447), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT38), .B1(new_n559), .B2(KEYINPUT37), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n558), .A2(new_n560), .B1(new_n448), .B2(new_n452), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n476), .A2(new_n456), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n454), .B1(new_n562), .B2(KEYINPUT37), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n448), .A2(new_n557), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT38), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n561), .A2(new_n565), .A3(new_n370), .A4(new_n369), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n556), .A2(new_n508), .A3(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n544), .B(new_n567), .C1(new_n479), .C2(new_n508), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n262), .B1(new_n541), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G57gat), .ZN(new_n570));
  OAI21_X1  g369(.A(G64gat), .B1(new_n570), .B2(KEYINPUT90), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT90), .ZN(new_n572));
  INV_X1    g371(.A(G64gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n573), .A3(G57gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(G71gat), .ZN(new_n577));
  INV_X1    g376(.A(G78gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT9), .ZN(new_n579));
  NAND2_X1  g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OR3_X1    g381(.A1(KEYINPUT89), .A2(G71gat), .A3(G78gat), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT89), .B1(G71gat), .B2(G78gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT9), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n573), .A2(G57gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n570), .A2(G64gat), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI22_X1  g388(.A1(new_n576), .A2(new_n582), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(new_n294), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n590), .A2(KEYINPUT91), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n590), .A2(KEYINPUT91), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n236), .B1(new_n598), .B2(new_n591), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n595), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G155gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n600), .A2(new_n604), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608));
  OR2_X1    g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(KEYINPUT92), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT92), .ZN(new_n612));
  AND2_X1   g411(.A1(G99gat), .A2(G106gat), .ZN(new_n613));
  NOR2_X1   g412(.A1(G99gat), .A2(G106gat), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT7), .ZN(new_n617));
  INV_X1    g416(.A(G85gat), .ZN(new_n618));
  INV_X1    g417(.A(G92gat), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n610), .A2(KEYINPUT8), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n619), .ZN(new_n622));
  NAND3_X1  g421(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n611), .A2(new_n615), .ZN(new_n626));
  AOI22_X1  g425(.A1(KEYINPUT8), .A2(new_n610), .B1(new_n618), .B2(new_n619), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n626), .A2(new_n627), .A3(new_n620), .A4(new_n623), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n629), .B1(new_n223), .B2(KEYINPUT17), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n222), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n223), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n632), .B1(new_n633), .B2(new_n629), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n631), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n637), .B1(new_n631), .B2(new_n634), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n608), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  INV_X1    g441(.A(new_n608), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n643), .A3(new_n638), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n641), .A2(new_n644), .A3(new_n646), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n607), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT10), .ZN(new_n652));
  INV_X1    g451(.A(new_n590), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n629), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT96), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(new_n616), .B2(new_n624), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n624), .A2(KEYINPUT95), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n627), .A2(new_n659), .A3(new_n620), .A4(new_n623), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n616), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n590), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT97), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n658), .A2(new_n616), .A3(new_n656), .A4(new_n660), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n662), .B2(new_n664), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n652), .B(new_n655), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n625), .A2(new_n628), .A3(KEYINPUT10), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT98), .B1(new_n598), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT98), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n668), .A2(new_n596), .A3(new_n671), .A4(new_n597), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(G230gat), .A2(G233gat), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n655), .B1(new_n665), .B2(new_n666), .ZN(new_n677));
  INV_X1    g476(.A(new_n675), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G120gat), .B(G148gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(G176gat), .B(G204gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n681), .B(new_n682), .Z(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n676), .A2(new_n679), .A3(new_n683), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n651), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n569), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n689), .A2(KEYINPUT99), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(KEYINPUT99), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n534), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(new_n225), .ZN(G1324gat));
  OAI21_X1  g493(.A(G8gat), .B1(new_n692), .B2(new_n537), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n692), .A2(new_n537), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT16), .B(G8gat), .Z(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n700), .A2(KEYINPUT100), .A3(KEYINPUT42), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n702), .B1(new_n699), .B2(new_n696), .ZN(new_n703));
  OAI221_X1 g502(.A(new_n695), .B1(new_n696), .B2(new_n699), .C1(new_n701), .C2(new_n703), .ZN(G1325gat));
  OAI21_X1  g503(.A(G15gat), .B1(new_n692), .B2(new_n544), .ZN(new_n705));
  INV_X1    g504(.A(G15gat), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n532), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n692), .B2(new_n707), .ZN(G1326gat));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n508), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT43), .B(G22gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n541), .A2(new_n568), .ZN(new_n713));
  INV_X1    g512(.A(new_n650), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n479), .B2(new_n508), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n534), .A2(new_n537), .ZN(new_n719));
  INV_X1    g518(.A(new_n508), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(new_n720), .A3(KEYINPUT101), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n544), .A2(new_n567), .A3(new_n718), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n541), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n723), .A2(KEYINPUT102), .A3(new_n712), .A4(new_n714), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n650), .B1(new_n541), .B2(new_n722), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT102), .B1(new_n726), .B2(new_n712), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n716), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n607), .A2(new_n687), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n257), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n728), .A2(KEYINPUT103), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n733));
  INV_X1    g532(.A(new_n533), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n535), .B(new_n520), .C1(new_n523), .C2(new_n522), .ZN(new_n735));
  INV_X1    g534(.A(new_n531), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n524), .B1(new_n736), .B2(KEYINPUT73), .ZN(new_n737));
  INV_X1    g536(.A(new_n507), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n497), .A2(new_n500), .B1(new_n503), .B2(new_n496), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n735), .B(new_n737), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT35), .B1(new_n719), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT82), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n538), .A2(KEYINPUT82), .A3(KEYINPUT35), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n734), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AND4_X1   g544(.A1(new_n544), .A2(new_n567), .A3(new_n721), .A4(new_n718), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n712), .B(new_n714), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n715), .B1(new_n749), .B2(new_n724), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n733), .B1(new_n750), .B2(new_n730), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n732), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G29gat), .B1(new_n752), .B2(new_n534), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n569), .A2(new_n714), .A3(new_n729), .ZN(new_n754));
  INV_X1    g553(.A(new_n534), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n209), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT45), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n753), .A2(new_n757), .ZN(G1328gat));
  OAI21_X1  g557(.A(G36gat), .B1(new_n752), .B2(new_n537), .ZN(new_n759));
  INV_X1    g558(.A(new_n537), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT104), .ZN(new_n761));
  AOI21_X1  g560(.A(G36gat), .B1(new_n761), .B2(KEYINPUT46), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n754), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n761), .A2(KEYINPUT46), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n759), .A2(new_n765), .ZN(G1329gat));
  INV_X1    g565(.A(G43gat), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n754), .A2(new_n767), .A3(new_n532), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n750), .A2(new_n544), .A3(new_n730), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n767), .ZN(new_n772));
  INV_X1    g571(.A(new_n544), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n732), .A2(new_n751), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n774), .A2(new_n775), .A3(G43gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n774), .B2(G43gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n776), .A2(new_n777), .A3(new_n768), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n772), .B1(new_n778), .B2(KEYINPUT47), .ZN(G1330gat));
  AND3_X1   g578(.A1(new_n754), .A2(new_n203), .A3(new_n720), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT48), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n750), .A2(new_n508), .A3(new_n730), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n203), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n732), .A2(new_n751), .A3(new_n720), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n780), .B1(new_n785), .B2(G50gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n786), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g586(.A(new_n687), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n651), .A2(new_n257), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n723), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n534), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(new_n570), .ZN(G1332gat));
  NOR2_X1   g591(.A1(new_n790), .A2(new_n537), .ZN(new_n793));
  NOR2_X1   g592(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n794));
  AND2_X1   g593(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n793), .B2(new_n794), .ZN(G1333gat));
  OAI21_X1  g596(.A(G71gat), .B1(new_n790), .B2(new_n544), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n532), .A2(new_n577), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n790), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g599(.A(new_n800), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g600(.A1(new_n790), .A2(new_n508), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(new_n578), .ZN(G1335gat));
  NOR2_X1   g602(.A1(new_n607), .A2(new_n257), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n726), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT106), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n806), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n807), .A2(KEYINPUT106), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n755), .A2(new_n618), .A3(new_n687), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n814), .B(KEYINPUT107), .Z(new_n815));
  NAND2_X1  g614(.A1(new_n804), .A2(new_n687), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n750), .A2(new_n534), .A3(new_n816), .ZN(new_n817));
  OAI22_X1  g616(.A1(new_n813), .A2(new_n815), .B1(new_n618), .B2(new_n817), .ZN(G1336gat));
  NOR2_X1   g617(.A1(new_n750), .A2(new_n816), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n760), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G92gat), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n807), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n809), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n788), .A2(G92gat), .A3(new_n537), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT109), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n821), .A2(new_n822), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT52), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(new_n812), .B2(new_n826), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n821), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1337gat));
  INV_X1    g633(.A(G99gat), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n812), .A2(new_n835), .A3(new_n532), .A4(new_n687), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n750), .A2(new_n544), .A3(new_n816), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT110), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n836), .B(KEYINPUT110), .C1(new_n835), .C2(new_n837), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1338gat));
  NOR2_X1   g641(.A1(new_n508), .A2(G106gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n812), .A2(new_n687), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n819), .A2(new_n720), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(G106gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n844), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n825), .A2(new_n687), .A3(new_n843), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n848), .B1(new_n850), .B2(new_n845), .ZN(G1339gat));
  INV_X1    g650(.A(new_n607), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n684), .B1(new_n676), .B2(KEYINPUT54), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n674), .B2(new_n675), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n667), .A2(new_n678), .A3(new_n673), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n857), .B1(new_n856), .B2(new_n858), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n854), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n854), .B(KEYINPUT55), .C1(new_n859), .C2(new_n860), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n863), .A2(new_n257), .A3(new_n686), .A4(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n235), .B1(new_n234), .B2(new_n238), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n866), .A2(KEYINPUT113), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(KEYINPUT113), .ZN(new_n868));
  OR3_X1    g667(.A1(new_n244), .A2(new_n237), .A3(new_n243), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n252), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n687), .A2(new_n871), .A3(new_n256), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n714), .B1(new_n865), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n860), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n853), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(KEYINPUT55), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n864), .A2(new_n686), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n648), .A2(new_n871), .A3(new_n256), .A4(new_n649), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n852), .B1(new_n873), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n257), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n607), .A2(new_n882), .A3(new_n650), .A4(new_n788), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT111), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n534), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n740), .A2(new_n760), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(G113gat), .B1(new_n887), .B2(new_n257), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n720), .B1(new_n881), .B2(new_n884), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n534), .A2(new_n760), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n894), .A2(new_n532), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n262), .A2(new_n283), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n888), .B1(new_n896), .B2(new_n897), .ZN(G1340gat));
  AOI21_X1  g697(.A(G120gat), .B1(new_n887), .B2(new_n687), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n788), .A2(new_n281), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n896), .B2(new_n900), .ZN(G1341gat));
  NAND2_X1  g700(.A1(new_n268), .A2(new_n269), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n893), .A2(new_n902), .A3(new_n607), .A4(new_n895), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT115), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n902), .B1(new_n887), .B2(new_n607), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(G1342gat));
  NAND3_X1  g707(.A1(new_n887), .A2(new_n274), .A3(new_n714), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n909), .A2(KEYINPUT56), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n714), .B(new_n895), .C1(new_n891), .C2(new_n892), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G134gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(KEYINPUT56), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT116), .Z(G1343gat));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n881), .A2(new_n884), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT119), .B1(new_n917), .B2(new_n755), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n919));
  AOI211_X1 g718(.A(new_n919), .B(new_n534), .C1(new_n881), .C2(new_n884), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n544), .A2(new_n720), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n760), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n302), .A3(new_n261), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT120), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n927));
  NOR4_X1   g726(.A1(new_n918), .A2(new_n920), .A3(new_n927), .A4(new_n924), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n544), .A2(new_n894), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT117), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT57), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n508), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n884), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n261), .A2(new_n863), .A3(new_n686), .A4(new_n864), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n714), .B1(new_n936), .B2(new_n872), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n852), .B1(new_n937), .B2(new_n880), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n935), .B1(new_n938), .B2(KEYINPUT118), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT118), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n940), .B(new_n852), .C1(new_n937), .C2(new_n880), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n934), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n508), .B1(new_n881), .B2(new_n884), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n943), .A2(KEYINPUT57), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n931), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(G141gat), .B1(new_n945), .B2(new_n882), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n916), .B1(new_n929), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(G141gat), .B1(new_n945), .B2(new_n262), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT58), .B1(new_n921), .B2(new_n925), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT121), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n918), .ZN(new_n952));
  INV_X1    g751(.A(new_n920), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(new_n953), .A3(new_n925), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n927), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n921), .A2(KEYINPUT120), .A3(new_n925), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(new_n931), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n255), .A2(KEYINPUT88), .A3(new_n256), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT88), .B1(new_n255), .B2(new_n256), .ZN(new_n960));
  OAI22_X1  g759(.A1(new_n876), .A2(KEYINPUT55), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n872), .B1(new_n961), .B2(new_n878), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n880), .B1(new_n962), .B2(new_n650), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT118), .B1(new_n963), .B2(new_n607), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n884), .A3(new_n941), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(new_n933), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n943), .A2(KEYINPUT57), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n958), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n302), .B1(new_n968), .B2(new_n257), .ZN(new_n969));
  OAI21_X1  g768(.A(KEYINPUT58), .B1(new_n957), .B2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT121), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n948), .A2(new_n916), .A3(new_n954), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n951), .A2(new_n973), .ZN(G1344gat));
  AND2_X1   g773(.A1(new_n921), .A2(new_n923), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n975), .A2(new_n303), .A3(new_n687), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT59), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n943), .A2(new_n932), .ZN(new_n978));
  INV_X1    g777(.A(new_n938), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n651), .A2(new_n261), .A3(new_n687), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n932), .B(new_n720), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n687), .B1(new_n931), .B2(KEYINPUT122), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n983), .B1(KEYINPUT122), .B2(new_n931), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n977), .B1(new_n985), .B2(G148gat), .ZN(new_n986));
  AOI211_X1 g785(.A(KEYINPUT59), .B(new_n303), .C1(new_n968), .C2(new_n687), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n976), .B1(new_n986), .B2(new_n987), .ZN(G1345gat));
  NAND3_X1  g787(.A1(new_n975), .A2(new_n307), .A3(new_n607), .ZN(new_n989));
  OAI21_X1  g788(.A(G155gat), .B1(new_n945), .B2(new_n852), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1346gat));
  INV_X1    g790(.A(new_n324), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n992), .A3(new_n714), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n968), .A2(new_n714), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n994), .A2(KEYINPUT123), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n324), .B1(new_n994), .B2(KEYINPUT123), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(G1347gat));
  NAND2_X1  g796(.A1(new_n917), .A2(new_n534), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n998), .B(KEYINPUT124), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n740), .A2(new_n537), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g800(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g801(.A(G169gat), .B1(new_n1002), .B2(new_n257), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n755), .A2(new_n537), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1004), .A2(new_n532), .ZN(new_n1005));
  XOR2_X1   g804(.A(new_n1005), .B(KEYINPUT125), .Z(new_n1006));
  AND2_X1   g805(.A1(new_n893), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n262), .A2(new_n389), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n1003), .B1(new_n1007), .B2(new_n1008), .ZN(G1348gat));
  NAND3_X1  g808(.A1(new_n1002), .A2(new_n390), .A3(new_n687), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1007), .A2(new_n687), .ZN(new_n1011));
  INV_X1    g810(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1010), .B1(new_n1012), .B2(new_n390), .ZN(G1349gat));
  NAND3_X1  g812(.A1(new_n893), .A2(new_n607), .A3(new_n1006), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1014), .A2(G183gat), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n607), .A2(new_n469), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1015), .B1(new_n1001), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1017), .A2(KEYINPUT60), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT60), .ZN(new_n1019));
  OAI211_X1 g818(.A(new_n1015), .B(new_n1019), .C1(new_n1001), .C2(new_n1016), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1018), .A2(new_n1020), .ZN(G1350gat));
  NAND3_X1  g820(.A1(new_n1002), .A2(new_n465), .A3(new_n714), .ZN(new_n1022));
  NAND3_X1  g821(.A1(new_n893), .A2(new_n714), .A3(new_n1006), .ZN(new_n1023));
  XNOR2_X1  g822(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1024));
  AND3_X1   g823(.A1(new_n1023), .A2(G190gat), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g824(.A(new_n1024), .B1(new_n1023), .B2(G190gat), .ZN(new_n1026));
  OAI21_X1  g825(.A(new_n1022), .B1(new_n1025), .B2(new_n1026), .ZN(G1351gat));
  NOR2_X1   g826(.A1(new_n922), .A2(new_n537), .ZN(new_n1028));
  AND2_X1   g827(.A1(new_n999), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g828(.A(G197gat), .B1(new_n1029), .B2(new_n257), .ZN(new_n1030));
  AND2_X1   g829(.A1(new_n544), .A2(new_n1004), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n982), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g831(.A(G197gat), .ZN(new_n1033));
  NOR3_X1   g832(.A1(new_n1032), .A2(new_n1033), .A3(new_n262), .ZN(new_n1034));
  NOR2_X1   g833(.A1(new_n1030), .A2(new_n1034), .ZN(G1352gat));
  XNOR2_X1  g834(.A(KEYINPUT127), .B(G204gat), .ZN(new_n1036));
  NOR2_X1   g835(.A1(new_n788), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n1029), .A2(new_n1037), .ZN(new_n1038));
  OR2_X1    g837(.A1(new_n1038), .A2(KEYINPUT62), .ZN(new_n1039));
  OAI21_X1  g838(.A(new_n1036), .B1(new_n1032), .B2(new_n788), .ZN(new_n1040));
  NAND2_X1  g839(.A1(new_n1038), .A2(KEYINPUT62), .ZN(new_n1041));
  NAND3_X1  g840(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(G1353gat));
  INV_X1    g841(.A(G211gat), .ZN(new_n1043));
  NAND3_X1  g842(.A1(new_n1029), .A2(new_n1043), .A3(new_n607), .ZN(new_n1044));
  NAND3_X1  g843(.A1(new_n982), .A2(new_n607), .A3(new_n1031), .ZN(new_n1045));
  NAND3_X1  g844(.A1(new_n1045), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1046));
  INV_X1    g845(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g846(.A(KEYINPUT63), .B1(new_n1045), .B2(G211gat), .ZN(new_n1048));
  OAI21_X1  g847(.A(new_n1044), .B1(new_n1047), .B2(new_n1048), .ZN(G1354gat));
  INV_X1    g848(.A(G218gat), .ZN(new_n1050));
  NAND3_X1  g849(.A1(new_n1029), .A2(new_n1050), .A3(new_n714), .ZN(new_n1051));
  OAI21_X1  g850(.A(G218gat), .B1(new_n1032), .B2(new_n650), .ZN(new_n1052));
  NAND2_X1  g851(.A1(new_n1051), .A2(new_n1052), .ZN(G1355gat));
endmodule


