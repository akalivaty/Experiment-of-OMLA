//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  AND2_X1   g0010(.A1(G116), .A2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n212), .A2(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n211), .B(new_n216), .C1(G87), .C2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G50), .A2(G226), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n203), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n210), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  OR3_X1    g0028(.A1(new_n210), .A2(KEYINPUT65), .A3(G13), .ZN(new_n229));
  OAI21_X1  g0029(.A(KEYINPUT65), .B1(new_n210), .B2(G13), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n231), .B(G250), .C1(G257), .C2(G264), .ZN(new_n232));
  INV_X1    g0032(.A(KEYINPUT0), .ZN(new_n233));
  OR2_X1    g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g0034(.A1(KEYINPUT66), .A2(G1), .A3(G13), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(KEYINPUT66), .B1(G1), .B2(G13), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(G20), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g0040(.A(G50), .ZN(new_n241));
  NOR2_X1   g0041(.A1(new_n206), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n232), .A2(new_n233), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n234), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n228), .A2(new_n246), .ZN(G361));
  XNOR2_X1  g0047(.A(G238), .B(G244), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G232), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT2), .B(G226), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G250), .B(G257), .Z(new_n252));
  XNOR2_X1  g0052(.A(G264), .B(G270), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G358));
  XOR2_X1   g0055(.A(G87), .B(G97), .Z(new_n256));
  XNOR2_X1  g0056(.A(G107), .B(G116), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XOR2_X1   g0058(.A(G68), .B(G77), .Z(new_n259));
  XNOR2_X1  g0059(.A(G50), .B(G58), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n258), .B(new_n261), .ZN(G351));
  OAI21_X1  g0062(.A(G20), .B1(new_n207), .B2(G50), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G20), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n265), .A2(new_n267), .B1(G150), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n237), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(new_n235), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G1), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G13), .A3(G20), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n270), .A2(new_n273), .B1(new_n241), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n273), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G1), .B2(new_n239), .ZN(new_n279));
  OR2_X1    g0079(.A1(new_n279), .A2(new_n241), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT9), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT9), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(new_n236), .B2(new_n237), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT3), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G33), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(G222), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT70), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(G1698), .ZN(new_n296));
  INV_X1    g0096(.A(G223), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n296), .A2(new_n297), .B1(new_n212), .B2(new_n292), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n288), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n274), .B1(G41), .B2(G45), .ZN(new_n300));
  INV_X1    g0100(.A(G274), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n286), .A2(KEYINPUT69), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT69), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(G33), .A3(G41), .ZN(new_n305));
  AND2_X1   g0105(.A1(G1), .A2(G13), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n300), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G226), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n299), .A2(G190), .A3(new_n302), .A4(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n283), .A2(new_n285), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G200), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n299), .A2(new_n302), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(new_n310), .ZN(new_n315));
  OR3_X1    g0115(.A1(new_n312), .A2(new_n315), .A3(KEYINPUT10), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT10), .B1(new_n312), .B2(new_n315), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT71), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n314), .A2(new_n310), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(G179), .ZN(new_n321));
  INV_X1    g0121(.A(G169), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n282), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G179), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n314), .A2(KEYINPUT71), .A3(new_n324), .A4(new_n310), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n321), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n276), .A2(new_n212), .ZN(new_n327));
  INV_X1    g0127(.A(new_n268), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n264), .A2(new_n328), .B1(new_n239), .B2(new_n212), .ZN(new_n329));
  XOR2_X1   g0129(.A(KEYINPUT15), .B(G87), .Z(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n267), .B2(new_n330), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n327), .B1(new_n279), .B2(new_n212), .C1(new_n331), .C2(new_n278), .ZN(new_n332));
  XOR2_X1   g0132(.A(new_n332), .B(KEYINPUT72), .Z(new_n333));
  OAI22_X1  g0133(.A1(new_n296), .A2(new_n224), .B1(new_n221), .B2(new_n292), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n289), .A2(new_n291), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n335), .A2(new_n220), .A3(G1698), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n288), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(new_n302), .C1(new_n213), .C2(new_n308), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G200), .ZN(new_n339));
  INV_X1    g0139(.A(G190), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n333), .B(new_n339), .C1(new_n340), .C2(new_n338), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n267), .A2(G77), .B1(new_n268), .B2(G50), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n203), .A2(G20), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n273), .ZN(new_n345));
  XOR2_X1   g0145(.A(new_n345), .B(KEYINPUT11), .Z(new_n346));
  INV_X1    g0146(.A(KEYINPUT74), .ZN(new_n347));
  INV_X1    g0147(.A(G13), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(G1), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n347), .B1(new_n350), .B2(new_n343), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n351), .A2(KEYINPUT12), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(KEYINPUT12), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n352), .B(new_n353), .C1(new_n279), .C2(new_n203), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n354), .A2(KEYINPUT75), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(KEYINPUT75), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n346), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT73), .ZN(new_n358));
  NOR2_X1   g0158(.A1(G226), .A2(G1698), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(new_n220), .B2(G1698), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n292), .A2(new_n360), .B1(G33), .B2(G97), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n302), .B1(new_n308), .B2(new_n224), .C1(new_n361), .C2(new_n287), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT13), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n361), .A2(new_n287), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n309), .A2(G238), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .A4(new_n302), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n358), .B1(new_n368), .B2(new_n340), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(G200), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n363), .A2(new_n367), .A3(KEYINPUT73), .A4(G190), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n357), .A2(new_n369), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n318), .A2(new_n326), .A3(new_n341), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n368), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT14), .B1(new_n374), .B2(new_n322), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(G179), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT14), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n368), .A2(new_n377), .A3(G169), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n355), .A2(new_n356), .ZN(new_n380));
  INV_X1    g0180(.A(new_n346), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n338), .A2(new_n322), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n384), .B(new_n332), .C1(G179), .C2(new_n338), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n202), .A2(new_n203), .ZN(new_n387));
  OAI21_X1  g0187(.A(G20), .B1(new_n206), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n268), .A2(G159), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT76), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n266), .B2(KEYINPUT3), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n289), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n266), .A3(KEYINPUT3), .ZN(new_n394));
  AOI21_X1  g0194(.A(G20), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  OAI21_X1  g0196(.A(G68), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT76), .B1(new_n290), .B2(G33), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n290), .A2(G33), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n394), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n239), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(KEYINPUT7), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n390), .B(KEYINPUT16), .C1(new_n397), .C2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n396), .B1(new_n292), .B2(G20), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n335), .A2(KEYINPUT7), .A3(new_n239), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n203), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n388), .A2(new_n389), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n404), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n403), .A2(new_n409), .A3(new_n273), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n265), .A2(new_n276), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n279), .B2(new_n265), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G87), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n297), .A2(new_n293), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n394), .B(new_n415), .C1(new_n398), .C2(new_n399), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n293), .A2(G226), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n288), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n307), .A2(G232), .A3(new_n300), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n420), .A2(new_n302), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n340), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n417), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n393), .A2(new_n394), .A3(new_n415), .A4(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n287), .B1(new_n424), .B2(new_n414), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n420), .A2(new_n302), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n313), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n410), .A2(new_n413), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT17), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n203), .B1(new_n401), .B2(KEYINPUT7), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n395), .A2(new_n396), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n408), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n278), .B1(new_n433), .B2(KEYINPUT16), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n412), .B1(new_n434), .B2(new_n409), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n419), .A2(new_n324), .A3(new_n421), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n322), .B1(new_n425), .B2(new_n426), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT77), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n438), .B1(new_n436), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT78), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(G169), .B1(new_n419), .B2(new_n421), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n425), .A2(G179), .A3(new_n426), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT77), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT78), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI211_X1 g0247(.A(KEYINPUT18), .B(new_n435), .C1(new_n441), .C2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT18), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n441), .A2(new_n447), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n410), .A2(new_n413), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n386), .A2(new_n430), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n373), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT79), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT79), .B1(new_n373), .B2(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT22), .ZN(new_n461));
  INV_X1    g0261(.A(G87), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n393), .A2(new_n239), .A3(new_n394), .A4(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n289), .A2(new_n291), .A3(new_n239), .A4(G87), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n461), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT87), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n239), .A2(G33), .A3(G116), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n221), .A2(G20), .ZN(new_n470));
  XOR2_X1   g0270(.A(new_n470), .B(KEYINPUT23), .Z(new_n471));
  NAND4_X1  g0271(.A1(new_n468), .A2(KEYINPUT24), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n467), .A2(KEYINPUT87), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT87), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(new_n464), .B2(new_n466), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n469), .B(new_n471), .C1(new_n473), .C2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT24), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n472), .A2(new_n478), .A3(new_n273), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n274), .A2(G33), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT80), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n275), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n266), .A2(G1), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(KEYINPUT80), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n273), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G107), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n350), .A2(new_n470), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n487), .B(KEYINPUT25), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n479), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n393), .B(new_n394), .C1(G250), .C2(G1698), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n293), .A2(G257), .ZN(new_n491));
  INV_X1    g0291(.A(G294), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n490), .A2(new_n491), .B1(new_n266), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n288), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT82), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT5), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(G41), .ZN(new_n497));
  INV_X1    g0297(.A(G41), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n274), .B(G45), .C1(new_n498), .C2(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n307), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G264), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n501), .A2(new_n301), .A3(new_n502), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n494), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(G169), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n509), .B1(new_n324), .B2(new_n508), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n489), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n493), .A2(new_n288), .B1(new_n504), .B2(G264), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n340), .A3(new_n507), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n508), .B2(G200), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n479), .A2(new_n514), .A3(new_n486), .A4(new_n488), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(G116), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G20), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n519), .B(new_n239), .C1(G33), .C2(new_n214), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n273), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT20), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n521), .B(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n350), .A2(new_n518), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n485), .A2(G116), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT21), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n215), .A2(new_n293), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n222), .A2(G1698), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n393), .A2(new_n394), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n335), .A2(G303), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT85), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n531), .A2(KEYINPUT85), .A3(new_n532), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n288), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n506), .B1(new_n504), .B2(G270), .ZN(new_n538));
  AOI211_X1 g0338(.A(new_n528), .B(new_n322), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(G179), .A3(new_n538), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n527), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n537), .A2(new_n538), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  INV_X1    g0344(.A(new_n527), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n544), .B(new_n545), .C1(new_n340), .C2(new_n543), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT86), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n322), .B1(new_n537), .B2(new_n538), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n527), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n549), .B2(new_n528), .ZN(new_n550));
  AOI211_X1 g0350(.A(KEYINPUT86), .B(KEYINPUT21), .C1(new_n548), .C2(new_n527), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n542), .B(new_n546), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n274), .A2(G45), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(new_n301), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n307), .A2(G250), .A3(new_n554), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n213), .A2(G1698), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(G238), .B2(G1698), .ZN(new_n558));
  OAI22_X1  g0358(.A1(new_n400), .A2(new_n558), .B1(new_n266), .B2(new_n517), .ZN(new_n559));
  AOI211_X1 g0359(.A(new_n555), .B(new_n556), .C1(new_n288), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n324), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n556), .B1(new_n559), .B2(new_n288), .ZN(new_n562));
  INV_X1    g0362(.A(new_n555), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n322), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n393), .A2(new_n239), .A3(G68), .A4(new_n394), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n267), .A2(G97), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT19), .ZN(new_n568));
  NAND3_X1  g0368(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n239), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G97), .A2(G107), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n462), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n567), .A2(new_n568), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n273), .ZN(new_n575));
  INV_X1    g0375(.A(new_n330), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n276), .ZN(new_n577));
  OR3_X1    g0377(.A1(new_n273), .A2(new_n482), .A3(new_n484), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n575), .B(new_n577), .C1(new_n576), .C2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n561), .A2(new_n565), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n564), .A2(new_n340), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n485), .A2(G87), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n575), .A2(new_n577), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n560), .B2(new_n313), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT83), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n584), .B(KEYINPUT83), .C1(new_n313), .C2(new_n560), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n581), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT7), .B1(new_n335), .B2(new_n239), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n396), .B(G20), .C1(new_n289), .C2(new_n291), .ZN(new_n591));
  OAI21_X1  g0391(.A(G107), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n328), .A2(new_n212), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT6), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n214), .A2(new_n221), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(new_n571), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n221), .A2(KEYINPUT6), .A3(G97), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n592), .B(new_n594), .C1(new_n239), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n273), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n275), .A2(G97), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n578), .A2(new_n214), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n601), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n289), .A2(new_n291), .A3(G250), .A4(G1698), .ZN(new_n607));
  AND2_X1   g0407(.A1(KEYINPUT4), .A2(G244), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n289), .A2(new_n291), .A3(new_n608), .A4(new_n293), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n609), .A3(new_n519), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT4), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n393), .A2(G244), .A3(new_n293), .A4(new_n394), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(new_n287), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n507), .B1(new_n503), .B2(new_n215), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n614), .A2(new_n615), .A3(new_n340), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n606), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n506), .B1(new_n504), .B2(G257), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n613), .A2(KEYINPUT81), .A3(new_n287), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT81), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n612), .A2(new_n611), .ZN(new_n621));
  INV_X1    g0421(.A(new_n610), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n620), .B1(new_n623), .B2(new_n288), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n618), .B1(new_n619), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G200), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n602), .B1(new_n600), .B2(new_n273), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n623), .A2(new_n288), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n618), .A2(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n627), .A2(new_n605), .B1(new_n629), .B2(new_n322), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n324), .B(new_n618), .C1(new_n619), .C2(new_n624), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n617), .A2(new_n626), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n589), .A2(new_n632), .A3(KEYINPUT84), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n614), .A2(new_n615), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G190), .ZN(new_n635));
  AOI211_X1 g0435(.A(new_n602), .B(new_n604), .C1(new_n600), .C2(new_n273), .ZN(new_n636));
  OAI21_X1  g0436(.A(KEYINPUT81), .B1(new_n613), .B2(new_n287), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n623), .A2(new_n620), .A3(new_n288), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n615), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n635), .B(new_n636), .C1(new_n313), .C2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n313), .B1(new_n562), .B2(new_n563), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n575), .A2(new_n577), .A3(new_n583), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n586), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n582), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n588), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n629), .A2(new_n322), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n631), .A2(new_n606), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n640), .A2(new_n645), .A3(new_n647), .A4(new_n580), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT84), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n516), .A2(new_n553), .A3(new_n633), .A4(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n460), .A2(new_n651), .ZN(G372));
  INV_X1    g0452(.A(new_n326), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n444), .A2(new_n446), .B1(new_n410), .B2(new_n413), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(new_n449), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n372), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n386), .A2(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n410), .A2(new_n413), .A3(new_n428), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT17), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n656), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n653), .B1(new_n661), .B2(new_n318), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n585), .A2(KEYINPUT88), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n582), .B1(new_n585), .B2(KEYINPUT88), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n581), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n515), .A2(new_n640), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n548), .A2(KEYINPUT21), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n545), .B1(new_n668), .B2(new_n540), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n549), .A2(new_n528), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT86), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n549), .A2(new_n547), .A3(new_n528), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n669), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n667), .B1(new_n673), .B2(new_n511), .ZN(new_n674));
  INV_X1    g0474(.A(new_n647), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n663), .B(new_n666), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  XOR2_X1   g0476(.A(new_n580), .B(KEYINPUT89), .Z(new_n677));
  NAND2_X1  g0477(.A1(new_n589), .A2(new_n675), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n677), .B1(new_n678), .B2(KEYINPUT26), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n662), .B1(new_n460), .B2(new_n681), .ZN(G369));
  NOR2_X1   g0482(.A1(new_n350), .A2(G20), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT27), .ZN(new_n684));
  OR3_X1    g0484(.A1(new_n683), .A2(KEYINPUT90), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G213), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n683), .B2(new_n684), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT90), .B1(new_n683), .B2(new_n684), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n685), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n489), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n516), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n691), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n511), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n542), .B1(new_n550), .B2(new_n551), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n545), .A2(new_n694), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n552), .B2(new_n697), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n695), .A2(G330), .A3(new_n699), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT91), .Z(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n673), .A2(new_n691), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n489), .A2(new_n510), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n703), .A2(new_n516), .B1(new_n704), .B2(new_n694), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n702), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n231), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n708), .A2(G116), .A3(new_n572), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n709), .A2(G1), .B1(new_n242), .B2(new_n708), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT92), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT28), .Z(new_n712));
  AOI211_X1 g0512(.A(KEYINPUT29), .B(new_n691), .C1(new_n676), .C2(new_n679), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT94), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n704), .B2(new_n696), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n673), .A2(KEYINPUT94), .A3(new_n511), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n666), .A2(new_n515), .A3(new_n632), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n589), .A2(new_n663), .A3(new_n675), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n666), .A2(new_n675), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT26), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT93), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n677), .B(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n719), .A2(new_n720), .A3(new_n722), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n714), .B1(new_n725), .B2(new_n694), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n512), .A2(new_n560), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n541), .A2(new_n727), .A3(new_n634), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n541), .A2(new_n727), .A3(KEYINPUT30), .A4(new_n634), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n512), .A2(new_n507), .B1(new_n537), .B2(new_n538), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(new_n625), .A3(new_n324), .A4(new_n564), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT31), .B1(new_n734), .B2(new_n691), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(new_n651), .B2(new_n691), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n713), .B(new_n726), .C1(G330), .C2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n712), .B1(new_n740), .B2(G1), .ZN(G364));
  NAND2_X1  g0541(.A1(new_n699), .A2(G330), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT95), .Z(new_n743));
  NOR2_X1   g0543(.A1(new_n348), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n274), .B1(new_n744), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n708), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n743), .B(new_n748), .C1(G330), .C2(new_n699), .ZN(new_n749));
  NOR3_X1   g0549(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT97), .Z(new_n751));
  OR2_X1    g0551(.A1(new_n699), .A2(new_n751), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n322), .A2(KEYINPUT98), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n322), .A2(KEYINPUT98), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n238), .B1(G20), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n239), .A2(new_n340), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n324), .A2(new_n313), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n239), .A2(G190), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n760), .A2(G326), .B1(new_n764), .B2(G329), .ZN(new_n765));
  INV_X1    g0565(.A(G303), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n313), .A2(G179), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n757), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n765), .B(new_n335), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(KEYINPUT101), .B(KEYINPUT33), .ZN(new_n770));
  INV_X1    g0570(.A(G317), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n758), .A2(new_n761), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n324), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n761), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n772), .A2(new_n774), .B1(G311), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G283), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n767), .A2(new_n761), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n239), .B1(new_n762), .B2(G190), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n778), .B1(new_n779), .B2(new_n780), .C1(new_n492), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n757), .A2(new_n775), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n769), .B(new_n782), .C1(G322), .C2(new_n788), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n776), .A2(KEYINPUT100), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n776), .A2(KEYINPUT100), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n781), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n793), .A2(G77), .B1(G97), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n202), .B2(new_n787), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n292), .B1(new_n780), .B2(new_n221), .ZN(new_n797));
  INV_X1    g0597(.A(new_n768), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G87), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n799), .B1(new_n773), .B2(new_n203), .C1(new_n241), .C2(new_n759), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n764), .A2(G159), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT32), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n796), .A2(new_n797), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n756), .B1(new_n789), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n400), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n707), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G45), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n242), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n806), .B(new_n808), .C1(new_n261), .C2(new_n807), .ZN(new_n809));
  INV_X1    g0609(.A(G355), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n231), .A2(new_n292), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n809), .B1(G116), .B2(new_n231), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT96), .Z(new_n813));
  INV_X1    g0613(.A(new_n751), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n756), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n752), .A2(new_n804), .A3(new_n747), .A4(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT102), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n749), .A2(new_n818), .ZN(G396));
  AOI21_X1  g0619(.A(new_n691), .B1(new_n676), .B2(new_n679), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n385), .A2(new_n691), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n332), .A2(new_n691), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n341), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n821), .B1(new_n823), .B2(new_n385), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n820), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n739), .A2(G330), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n748), .ZN(new_n829));
  NOR2_X1   g0629(.A1(G13), .A2(G33), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n748), .B1(new_n825), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n756), .A2(new_n830), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n212), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n788), .A2(G294), .B1(new_n793), .B2(G116), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n774), .A2(G283), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n335), .B1(new_n768), .B2(new_n221), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT103), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n759), .A2(new_n766), .B1(new_n780), .B2(new_n462), .ZN(new_n838));
  INV_X1    g0638(.A(G311), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n839), .A2(new_n763), .B1(new_n781), .B2(new_n214), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n834), .A2(new_n835), .A3(new_n837), .A4(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n788), .A2(G143), .B1(new_n793), .B2(G159), .ZN(new_n843));
  INV_X1    g0643(.A(G137), .ZN(new_n844));
  INV_X1    g0644(.A(G150), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n843), .B1(new_n844), .B2(new_n759), .C1(new_n845), .C2(new_n773), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT34), .Z(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n780), .A2(new_n203), .B1(new_n763), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n805), .B1(new_n241), .B2(new_n768), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n849), .B(new_n850), .C1(G58), .C2(new_n794), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT104), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n842), .B1(new_n847), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n756), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n831), .A2(new_n833), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n829), .A2(new_n855), .ZN(G384));
  NAND2_X1  g0656(.A1(new_n459), .A2(new_n739), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT111), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n379), .A2(new_n382), .A3(new_n694), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n382), .A2(new_n691), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n379), .A2(new_n382), .B1(new_n372), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT106), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n372), .A2(new_n860), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n383), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT106), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n379), .A2(new_n382), .A3(new_n694), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n511), .B(new_n515), .C1(new_n648), .C2(new_n649), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT84), .B1(new_n589), .B2(new_n632), .ZN(new_n870));
  NOR4_X1   g0670(.A1(new_n869), .A2(new_n870), .A3(new_n552), .A4(new_n691), .ZN(new_n871));
  INV_X1    g0671(.A(new_n737), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n735), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n868), .B(new_n824), .C1(new_n871), .C2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT110), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT108), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n390), .B1(new_n397), .B2(new_n402), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n404), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n412), .B1(new_n434), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(new_n689), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n453), .B2(new_n430), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n435), .B1(new_n441), .B2(new_n447), .ZN(new_n884));
  INV_X1    g0684(.A(new_n689), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n451), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT37), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(new_n887), .A3(new_n429), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT107), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n879), .A2(new_n273), .A3(new_n403), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n891), .A2(new_n413), .B1(new_n444), .B2(new_n446), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n890), .B1(new_n892), .B2(new_n659), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n439), .A2(new_n440), .ZN(new_n894));
  OAI211_X1 g0694(.A(KEYINPUT107), .B(new_n429), .C1(new_n894), .C2(new_n880), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n893), .A2(new_n882), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n889), .B1(new_n896), .B2(KEYINPUT37), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n876), .B(new_n877), .C1(new_n883), .C2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n877), .B1(new_n883), .B2(new_n897), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n900));
  INV_X1    g0700(.A(new_n889), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n439), .A2(new_n440), .A3(KEYINPUT78), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n445), .B1(new_n444), .B2(new_n446), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n451), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT18), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n884), .A2(new_n449), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n430), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n881), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n902), .A2(KEYINPUT38), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n899), .A2(KEYINPUT108), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT110), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n739), .A2(new_n824), .A3(new_n868), .A4(new_n913), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n875), .A2(new_n898), .A3(new_n911), .A4(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n886), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n655), .B2(new_n660), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n451), .B1(new_n440), .B2(new_n439), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(new_n429), .A3(new_n886), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT37), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n884), .B2(new_n888), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT38), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n900), .A2(new_n901), .B1(new_n908), .B2(new_n881), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n922), .B1(new_n923), .B2(KEYINPUT38), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT40), .B1(new_n874), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n915), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n858), .B(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(G330), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT112), .Z(new_n929));
  OAI21_X1  g0729(.A(new_n459), .B1(new_n726), .B2(new_n713), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n662), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT109), .B1(new_n924), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n917), .A2(new_n921), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n877), .ZN(new_n936));
  AND4_X1   g0736(.A1(KEYINPUT109), .A2(new_n910), .A3(new_n933), .A4(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n911), .A2(KEYINPUT39), .A3(new_n898), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n859), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n656), .A2(new_n885), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n680), .A2(new_n694), .A3(new_n824), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n821), .B(KEYINPUT105), .Z(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n946), .A2(new_n868), .A3(new_n898), .A4(new_n911), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n940), .A2(new_n942), .A3(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n932), .B(new_n948), .Z(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n274), .B2(new_n744), .ZN(new_n950));
  INV_X1    g0750(.A(new_n599), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n517), .B1(new_n951), .B2(KEYINPUT35), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n952), .B(new_n240), .C1(KEYINPUT35), .C2(new_n951), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT36), .ZN(new_n954));
  INV_X1    g0754(.A(new_n242), .ZN(new_n955));
  OAI21_X1  g0755(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n955), .A2(new_n956), .B1(G50), .B2(new_n203), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n957), .A2(G1), .A3(new_n348), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n950), .A2(new_n954), .A3(new_n958), .ZN(G367));
  INV_X1    g0759(.A(G159), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n792), .A2(new_n241), .B1(new_n960), .B2(new_n773), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT115), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n798), .A2(G58), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n292), .B1(new_n780), .B2(new_n212), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT116), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n964), .A2(new_n965), .B1(G143), .B2(new_n760), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n787), .A2(new_n845), .B1(new_n965), .B2(new_n964), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n844), .A2(new_n763), .B1(new_n781), .B2(new_n203), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n962), .A2(new_n963), .A3(new_n966), .A4(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n780), .A2(new_n214), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n971), .B(new_n805), .C1(G317), .C2(new_n764), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT114), .Z(new_n973));
  AOI22_X1  g0773(.A1(new_n788), .A2(G303), .B1(new_n793), .B2(G283), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n221), .B2(new_n781), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n976), .B1(new_n492), .B2(new_n773), .C1(new_n839), .C2(new_n759), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n768), .A2(new_n517), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT46), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n970), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT117), .Z(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT47), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n756), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n677), .A2(new_n642), .A3(new_n691), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n666), .B1(new_n584), .B2(new_n694), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n984), .A2(new_n814), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n806), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n815), .B1(new_n231), .B2(new_n576), .C1(new_n987), .C2(new_n254), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n983), .A2(new_n747), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n632), .B1(new_n636), .B2(new_n694), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT113), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n675), .A2(new_n691), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(new_n705), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT44), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n705), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT45), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n997), .B(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(new_n701), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n703), .A2(new_n516), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n695), .B2(new_n703), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n743), .A2(new_n1003), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n1004), .A2(new_n700), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n740), .A2(new_n1005), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n740), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n708), .B(KEYINPUT41), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n746), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n994), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1011), .A2(new_n1002), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT42), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n647), .B1(new_n992), .B2(new_n511), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n694), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n984), .A2(new_n985), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1013), .A2(new_n1015), .B1(KEYINPUT43), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(KEYINPUT43), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n702), .A2(new_n1011), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n989), .B1(new_n1010), .B2(new_n1021), .ZN(G387));
  OAI21_X1  g0822(.A(new_n806), .B1(new_n251), .B2(new_n807), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n572), .A2(G116), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1023), .B1(new_n1024), .B2(new_n811), .ZN(new_n1025));
  OR3_X1    g0825(.A1(new_n264), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1026));
  OAI21_X1  g0826(.A(KEYINPUT50), .B1(new_n264), .B2(G50), .ZN(new_n1027));
  AOI21_X1  g0827(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1024), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n707), .A2(new_n221), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n756), .B(new_n814), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n794), .A2(new_n330), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n845), .B2(new_n763), .C1(new_n264), .C2(new_n773), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n805), .B1(new_n214), .B2(new_n780), .C1(new_n787), .C2(new_n241), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(G77), .C2(new_n798), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n203), .B2(new_n776), .C1(new_n960), .C2(new_n759), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n788), .A2(G317), .B1(new_n793), .B2(G303), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n760), .A2(G322), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(new_n839), .C2(new_n773), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT48), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n779), .B2(new_n781), .C1(new_n492), .C2(new_n768), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT49), .Z(new_n1043));
  INV_X1    g0843(.A(new_n780), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G116), .A2(new_n1044), .B1(new_n764), .B2(G326), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n400), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1037), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n748), .B(new_n1032), .C1(new_n1047), .C2(new_n756), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n695), .A2(new_n751), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1005), .A2(new_n746), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1006), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n708), .B1(new_n740), .B2(new_n1005), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(G393));
  NAND3_X1  g0853(.A1(new_n1000), .A2(KEYINPUT118), .A3(new_n701), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n1001), .B2(KEYINPUT118), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1007), .B(new_n708), .C1(new_n1055), .C2(new_n1051), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n815), .B1(new_n214), .B2(new_n231), .C1(new_n987), .C2(new_n258), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n747), .B(new_n1057), .C1(new_n994), .C2(new_n751), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n788), .A2(G159), .B1(G150), .B2(new_n760), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n1059), .A2(KEYINPUT51), .B1(new_n241), .B2(new_n773), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n265), .B2(new_n793), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(KEYINPUT51), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n781), .A2(new_n212), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n400), .B(new_n1063), .C1(G87), .C2(new_n1044), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G68), .A2(new_n798), .B1(new_n764), .B2(G143), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n787), .A2(new_n839), .B1(new_n771), .B2(new_n759), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT52), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n292), .B1(new_n1044), .B2(G107), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n764), .A2(G322), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n773), .A2(new_n766), .B1(new_n776), .B2(new_n492), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G116), .B2(new_n794), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n768), .A2(new_n779), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1066), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1058), .B1(new_n756), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n1055), .B2(new_n746), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1056), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(KEYINPUT119), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT119), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1056), .A2(new_n1080), .A3(new_n1077), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1081), .ZN(G390));
  NOR2_X1   g0882(.A1(new_n924), .A2(new_n859), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n725), .A2(new_n694), .A3(new_n824), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1084), .A2(new_n945), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n868), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT109), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n910), .A2(new_n936), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1088), .B1(new_n1089), .B2(KEYINPUT39), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n924), .A2(KEYINPUT109), .A3(new_n933), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n911), .A2(KEYINPUT39), .A3(new_n898), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n859), .B1(new_n946), .B2(new_n868), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1087), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OR4_X1    g0896(.A1(new_n869), .A2(new_n870), .A3(new_n552), .A4(new_n691), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n825), .B1(new_n1097), .B2(new_n738), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT120), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1098), .A2(new_n1099), .A3(G330), .A4(new_n868), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n739), .A2(G330), .A3(new_n824), .A4(new_n868), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(KEYINPUT120), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1096), .A2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1087), .B(new_n1101), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n739), .A2(G330), .A3(new_n824), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n1086), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1100), .A2(new_n1102), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n946), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1085), .A2(new_n1101), .A3(new_n1108), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n459), .A2(G330), .A3(new_n739), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n930), .A2(new_n1113), .A3(new_n662), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1106), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1114), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1104), .A2(new_n1118), .A3(new_n1105), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n708), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1104), .A2(new_n746), .A3(new_n1105), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT123), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1092), .A2(new_n830), .A3(new_n1093), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n832), .A2(new_n264), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n792), .A2(new_n214), .B1(new_n221), .B2(new_n773), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT122), .Z(new_n1126));
  NAND2_X1  g0926(.A1(new_n788), .A2(G116), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n760), .A2(G283), .B1(new_n1044), .B2(G68), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1126), .A2(new_n799), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n763), .A2(new_n492), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n1129), .A2(new_n292), .A3(new_n1063), .A4(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n760), .A2(G128), .B1(new_n794), .B2(G159), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n335), .B1(new_n774), .B2(G137), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(new_n241), .C2(new_n780), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n768), .A2(new_n845), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT121), .Z(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1136), .B1(new_n787), .B2(new_n848), .C1(new_n1139), .C2(new_n792), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1134), .B(new_n1140), .C1(G125), .C2(new_n764), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n756), .B1(new_n1131), .B2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1123), .A2(new_n747), .A3(new_n1124), .A4(new_n1142), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1121), .A2(new_n1122), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1122), .B1(new_n1121), .B2(new_n1143), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1120), .B1(new_n1144), .B2(new_n1145), .ZN(G378));
  NAND2_X1  g0946(.A1(new_n318), .A2(new_n326), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n281), .A2(new_n885), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1147), .B(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n830), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n788), .A2(G128), .B1(G132), .B2(new_n774), .ZN(new_n1156));
  INV_X1    g0956(.A(G125), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n759), .A2(new_n1157), .B1(new_n781), .B2(new_n845), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G137), .B2(new_n777), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1156), .B(new_n1159), .C1(new_n768), .C2(new_n1139), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT59), .Z(new_n1161));
  OAI21_X1  g0961(.A(new_n266), .B1(new_n780), .B2(new_n960), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G124), .B2(new_n764), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1161), .A2(new_n498), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G41), .B1(new_n805), .B2(G33), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1164), .B1(G50), .B2(new_n1165), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n576), .A2(new_n776), .B1(new_n203), .B2(new_n781), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n805), .B(new_n1167), .C1(G77), .C2(new_n798), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n498), .B1(new_n780), .B2(new_n202), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n759), .A2(new_n517), .B1(new_n763), .B2(new_n779), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1169), .B(new_n1170), .C1(G97), .C2(new_n774), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1168), .B(new_n1171), .C1(new_n221), .C2(new_n787), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT58), .Z(new_n1173));
  OAI21_X1  g0973(.A(new_n756), .B1(new_n1166), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n832), .A2(new_n241), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1155), .A2(new_n747), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(G330), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n915), .B2(new_n925), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n948), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n926), .A2(G330), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1181), .A2(new_n942), .A3(new_n947), .A4(new_n940), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n1153), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n1182), .A3(new_n1154), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1177), .B1(new_n1186), .B2(new_n746), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1184), .A2(new_n1185), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n708), .B1(new_n1188), .B2(KEYINPUT57), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1119), .A2(new_n1115), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1180), .A2(new_n1154), .A3(new_n1182), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1154), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1190), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1187), .B1(new_n1189), .B2(new_n1195), .ZN(G375));
  AOI22_X1  g0996(.A1(new_n793), .A2(G107), .B1(G116), .B2(new_n774), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1197), .A2(KEYINPUT124), .B1(G283), .B2(new_n788), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n492), .B2(new_n759), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1197), .A2(KEYINPUT124), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n768), .A2(new_n214), .B1(new_n763), .B2(new_n766), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT126), .Z(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1033), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n335), .B1(new_n780), .B2(new_n212), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT125), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1199), .A2(new_n1200), .A3(new_n1203), .A4(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1138), .A2(new_n774), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n760), .A2(G132), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n764), .A2(G128), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G159), .A2(new_n798), .B1(new_n1044), .B2(G58), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n787), .A2(new_n844), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n781), .A2(new_n241), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n805), .B1(new_n845), .B2(new_n776), .ZN(new_n1214));
  NOR4_X1   g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n756), .B1(new_n1206), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n830), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n747), .B(new_n1216), .C1(new_n868), .C2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n203), .B2(new_n832), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1112), .B2(new_n746), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1110), .A2(new_n1114), .A3(new_n1111), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1009), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1220), .B1(new_n1222), .B2(new_n1118), .ZN(G381));
  OAI21_X1  g1023(.A(new_n746), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1176), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n708), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1188), .A2(KEYINPUT57), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1225), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1121), .A2(new_n1143), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1120), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1233), .A2(G384), .A3(G381), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(G390), .A2(G387), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(G393), .A2(G396), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(G407));
  OAI211_X1 g1037(.A(G407), .B(G213), .C1(G343), .C2(new_n1233), .ZN(G409));
  NAND2_X1  g1038(.A1(G390), .A2(G387), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  XOR2_X1   g1040(.A(G393), .B(G396), .Z(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1240), .A2(new_n1235), .A3(new_n1242), .ZN(new_n1243));
  OR2_X1    g1043(.A1(G390), .A2(G387), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1241), .B1(new_n1244), .B2(new_n1239), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n686), .A2(G343), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G378), .B(new_n1187), .C1(new_n1189), .C2(new_n1195), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1186), .A2(new_n1009), .A3(new_n1190), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1231), .B1(new_n1187), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1247), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT60), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1116), .B(new_n708), .C1(new_n1253), .C2(new_n1221), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1221), .A2(new_n1253), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1220), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(G384), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT62), .B1(new_n1252), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1250), .B1(new_n1229), .B2(G378), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT127), .B1(new_n1262), .B2(new_n1247), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT127), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1247), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1261), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1247), .A2(G2897), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1260), .A2(new_n1272), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1258), .A2(new_n1259), .A3(new_n1271), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1263), .A2(new_n1267), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1246), .B1(new_n1270), .B2(new_n1279), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1268), .A2(KEYINPUT63), .A3(new_n1260), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT63), .B1(new_n1252), .B2(new_n1275), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1252), .A2(new_n1260), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT61), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1281), .A2(new_n1282), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1280), .A2(new_n1286), .ZN(G405));
  OAI21_X1  g1087(.A(new_n1248), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1288), .B(new_n1260), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1246), .B(new_n1289), .ZN(G402));
endmodule


