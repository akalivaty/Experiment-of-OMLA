//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G128), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT93), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G128), .B(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT93), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n195), .A3(G134), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G116), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G122), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n201), .A2(G122), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT14), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n204), .B1(new_n203), .B2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n202), .A2(KEYINPUT94), .A3(KEYINPUT14), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT94), .B1(new_n202), .B2(KEYINPUT14), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G107), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n200), .A2(new_n207), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n205), .B(new_n206), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n194), .A2(KEYINPUT13), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n217), .B(G134), .C1(KEYINPUT13), .C2(new_n188), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n198), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT9), .B(G234), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n221), .B(KEYINPUT80), .ZN(new_n222));
  INV_X1    g036(.A(G217), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n222), .A2(new_n223), .A3(G953), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n215), .A2(new_n219), .A3(new_n224), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G902), .ZN(new_n229));
  INV_X1    g043(.A(G478), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT15), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n228), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT95), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(new_n228), .B2(new_n229), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n215), .A2(new_n219), .A3(new_n224), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n224), .B1(new_n215), .B2(new_n219), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n235), .B(new_n229), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n231), .B1(new_n236), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT96), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n234), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(G475), .A2(G902), .ZN(new_n244));
  INV_X1    g058(.A(G237), .ZN(new_n245));
  INV_X1    g059(.A(G953), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(G214), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(G143), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT18), .A2(G131), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT88), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n247), .B(new_n187), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT88), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT18), .A4(G131), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n250), .A2(new_n253), .B1(new_n248), .B2(new_n249), .ZN(new_n254));
  INV_X1    g068(.A(G140), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G125), .ZN(new_n256));
  INV_X1    g070(.A(G125), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G140), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT78), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(G125), .B(G140), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT78), .ZN(new_n263));
  INV_X1    g077(.A(G146), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n259), .A2(G146), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT89), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n266), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT89), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n254), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT91), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n262), .A2(KEYINPUT16), .ZN(new_n273));
  OR3_X1    g087(.A1(new_n257), .A2(KEYINPUT16), .A3(G140), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(G146), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(G146), .B1(new_n273), .B2(new_n274), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n272), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n277), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(KEYINPUT91), .A3(new_n275), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n251), .A2(G131), .ZN(new_n281));
  INV_X1    g095(.A(G131), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n248), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT17), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n281), .A2(KEYINPUT17), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n278), .B(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(G113), .B(G122), .ZN(new_n287));
  INV_X1    g101(.A(G104), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n287), .B(new_n288), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n271), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n276), .B1(new_n281), .B2(new_n283), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT19), .B1(new_n261), .B2(KEYINPUT90), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT78), .B1(KEYINPUT90), .B2(KEYINPUT19), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n259), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n264), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n289), .B1(new_n271), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n244), .B1(new_n290), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT92), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT20), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n289), .B1(new_n271), .B2(new_n286), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n229), .B1(new_n290), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G475), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n298), .A2(new_n299), .ZN(new_n306));
  OAI211_X1 g120(.A(KEYINPUT92), .B(new_n244), .C1(new_n290), .C2(new_n297), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(KEYINPUT20), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n229), .B1(new_n237), .B2(new_n238), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT95), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n239), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT96), .A3(new_n231), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n243), .A2(new_n305), .A3(new_n308), .A4(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n246), .A2(G952), .ZN(new_n314));
  INV_X1    g128(.A(G234), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(new_n245), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  AOI211_X1 g131(.A(new_n229), .B(new_n246), .C1(G234), .C2(G237), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT21), .B(G898), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT97), .B1(new_n313), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n241), .A2(new_n242), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n322), .A2(new_n312), .A3(new_n233), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT97), .ZN(new_n324));
  INV_X1    g138(.A(new_n320), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n307), .A2(KEYINPUT20), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n271), .A2(new_n286), .A3(new_n289), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n270), .A2(new_n267), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n328), .A2(new_n254), .B1(new_n295), .B2(new_n291), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n329), .B2(new_n289), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT92), .B1(new_n330), .B2(new_n244), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n304), .B(new_n301), .C1(new_n326), .C2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n323), .A2(new_n324), .A3(new_n325), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n321), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(G214), .B1(G237), .B2(G902), .ZN(new_n336));
  XNOR2_X1  g150(.A(G110), .B(G122), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(G116), .B(G119), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT5), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n201), .A2(KEYINPUT5), .A3(G119), .ZN(new_n341));
  INV_X1    g155(.A(G113), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT2), .B(G113), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n340), .A2(new_n343), .B1(new_n345), .B2(new_n339), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT83), .B1(new_n206), .B2(G104), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT83), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n288), .A3(G107), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n206), .A2(G104), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G101), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT3), .B1(new_n288), .B2(G107), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n206), .A3(G104), .ZN(new_n355));
  INV_X1    g169(.A(G101), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n288), .A2(G107), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n353), .A2(new_n355), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n352), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(KEYINPUT84), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(new_n352), .B2(new_n358), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n346), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT85), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT85), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n365), .B(new_n346), .C1(new_n360), .C2(new_n362), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n353), .A2(new_n355), .A3(new_n357), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G101), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(KEYINPUT4), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n344), .B(new_n339), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n358), .A2(KEYINPUT4), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n369), .A2(KEYINPUT81), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(new_n368), .B2(G101), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n375), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(KEYINPUT82), .B(new_n375), .C1(new_n376), .C2(new_n378), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n374), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n338), .B1(new_n367), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n364), .A2(new_n366), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n379), .A2(new_n380), .ZN(new_n386));
  INV_X1    g200(.A(new_n382), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n385), .B(new_n337), .C1(new_n388), .C2(new_n374), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n384), .A2(KEYINPUT6), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n264), .A2(G143), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n187), .A2(G146), .ZN(new_n392));
  NAND2_X1  g206(.A1(KEYINPUT0), .A2(G128), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  OR2_X1    g208(.A1(KEYINPUT0), .A2(G128), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n395), .A2(new_n393), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n391), .A2(new_n392), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OR3_X1    g212(.A1(new_n398), .A2(KEYINPUT86), .A3(new_n257), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT86), .B1(new_n398), .B2(new_n257), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n391), .A2(new_n392), .ZN(new_n401));
  OR3_X1    g215(.A1(new_n401), .A2(KEYINPUT1), .A3(new_n189), .ZN(new_n402));
  INV_X1    g216(.A(new_n392), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n401), .A2(new_n189), .B1(new_n403), .B2(KEYINPUT1), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n399), .B(new_n400), .C1(G125), .C2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G224), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(G953), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n406), .B(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n410), .B(new_n338), .C1(new_n367), .C2(new_n383), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n390), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(G210), .B1(G237), .B2(G902), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT87), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT7), .B1(new_n407), .B2(G953), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n406), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n414), .B1(new_n406), .B2(new_n415), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n406), .A2(new_n415), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n337), .B(KEYINPUT8), .Z(new_n419));
  INV_X1    g233(.A(new_n359), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n420), .A2(new_n346), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n419), .B1(new_n363), .B2(new_n421), .ZN(new_n422));
  NOR4_X1   g236(.A1(new_n416), .A2(new_n417), .A3(new_n418), .A4(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(G902), .B1(new_n423), .B2(new_n389), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n412), .A2(new_n413), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n413), .B1(new_n412), .B2(new_n424), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n336), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n335), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n391), .A2(new_n392), .B1(new_n395), .B2(new_n393), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT66), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT66), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n394), .B(new_n434), .C1(new_n396), .C2(new_n397), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G137), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT64), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT64), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G137), .ZN(new_n440));
  AND2_X1   g254(.A1(KEYINPUT11), .A2(G134), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(KEYINPUT11), .A2(G134), .ZN(new_n443));
  NOR2_X1   g257(.A1(KEYINPUT11), .A2(G134), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(G137), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G131), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT65), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n442), .A2(new_n282), .A3(new_n445), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n446), .A2(KEYINPUT65), .A3(G131), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n436), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT67), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n438), .A2(new_n440), .A3(new_n197), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n282), .B1(G134), .B2(G137), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n457), .A2(KEYINPUT68), .B1(new_n402), .B2(new_n404), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT68), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n449), .A2(new_n459), .A3(new_n456), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT67), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n436), .A2(new_n450), .A3(new_n462), .A4(new_n451), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n453), .A2(new_n372), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT70), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n450), .A2(new_n451), .A3(new_n398), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n405), .A2(new_n449), .A3(new_n456), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT30), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n373), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(new_n458), .B2(new_n460), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n453), .A2(new_n463), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT69), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT69), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n453), .A2(new_n472), .A3(new_n475), .A4(new_n463), .ZN(new_n476));
  AOI211_X1 g290(.A(new_n465), .B(new_n471), .C1(new_n474), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n476), .ZN(new_n478));
  INV_X1    g292(.A(new_n471), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT70), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n464), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT26), .B(G101), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n245), .A2(new_n246), .A3(G210), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT29), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n468), .A2(new_n373), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n464), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT28), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT28), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n461), .A2(new_n452), .A3(new_n372), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n492), .A2(KEYINPUT73), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT73), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n496), .A3(KEYINPUT28), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n495), .A2(KEYINPUT74), .A3(new_n486), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n492), .A2(KEYINPUT73), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n494), .A2(new_n493), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n499), .A2(new_n486), .A3(new_n497), .A4(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT74), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n488), .A2(new_n489), .A3(new_n498), .A4(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n453), .A2(new_n461), .A3(new_n463), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n373), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT75), .A3(new_n464), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT75), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n508), .A3(new_n373), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n507), .A2(KEYINPUT28), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n500), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n511), .A2(new_n489), .A3(new_n487), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(G902), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G472), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n464), .A2(new_n486), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT72), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n477), .B2(new_n480), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT31), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n495), .A2(new_n497), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n487), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT31), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n518), .B(new_n523), .C1(new_n477), .C2(new_n480), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n520), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(G472), .A2(G902), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT32), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n525), .A2(KEYINPUT32), .A3(new_n526), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n515), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  XOR2_X1   g345(.A(G119), .B(G128), .Z(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT24), .B(G110), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n189), .A2(KEYINPUT23), .A3(G119), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT76), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT77), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n538), .A2(KEYINPUT23), .B1(new_n189), .B2(G119), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n538), .B2(KEYINPUT23), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n537), .B(new_n540), .C1(G119), .C2(new_n189), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n534), .B1(new_n541), .B2(G110), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n277), .B2(new_n276), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n532), .A2(new_n533), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n541), .B2(G110), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n275), .A3(new_n265), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n246), .A2(G221), .A3(G234), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT22), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(G137), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n543), .A2(new_n546), .A3(new_n550), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n223), .B1(G234), .B2(new_n229), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(G902), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT79), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n552), .A2(new_n229), .A3(new_n553), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n560), .A2(KEYINPUT25), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(KEYINPUT25), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n555), .A3(new_n562), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G221), .B1(new_n222), .B2(G902), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n371), .A2(new_n436), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n381), .B2(new_n382), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n420), .A2(new_n405), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT10), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n360), .A2(new_n362), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n405), .A2(KEYINPUT10), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n450), .A2(new_n451), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n567), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(G110), .B(G140), .ZN(new_n577));
  INV_X1    g391(.A(G227), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(G953), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n577), .B(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n575), .B1(new_n567), .B2(new_n573), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OR2_X1    g397(.A1(new_n360), .A2(new_n362), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n568), .B1(new_n584), .B2(new_n405), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n575), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT12), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(KEYINPUT12), .A3(new_n575), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n576), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n580), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n583), .B(G469), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(G469), .A2(G902), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n588), .A2(new_n589), .ZN(new_n595));
  INV_X1    g409(.A(new_n566), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n386), .B2(new_n387), .ZN(new_n597));
  INV_X1    g411(.A(new_n572), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n584), .A2(new_n598), .B1(new_n569), .B2(new_n568), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n599), .A3(new_n574), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n582), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n595), .A2(new_n581), .B1(new_n601), .B2(new_n580), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n602), .A2(G469), .A3(G902), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n565), .B1(new_n594), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n430), .A2(new_n531), .A3(new_n564), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  INV_X1    g421(.A(new_n527), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n525), .A2(new_n229), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n525), .A2(KEYINPUT98), .A3(new_n229), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(G472), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n608), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n611), .A2(KEYINPUT99), .A3(G472), .A4(new_n612), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n605), .A2(new_n564), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n412), .A2(new_n424), .ZN(new_n620));
  INV_X1    g434(.A(new_n413), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n412), .A2(new_n424), .A3(new_n413), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n225), .B2(KEYINPUT100), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n228), .B(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n230), .A2(G902), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n311), .A2(new_n230), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n332), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n624), .A2(new_n633), .A3(new_n325), .A4(new_n336), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n619), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT34), .B(G104), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  AOI21_X1  g452(.A(new_n332), .B1(new_n243), .B2(new_n312), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n624), .A2(new_n325), .A3(new_n639), .A4(new_n336), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n617), .A2(new_n618), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT35), .B(G107), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NAND2_X1  g457(.A1(new_n613), .A2(new_n614), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n551), .A2(KEYINPUT36), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n547), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n556), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n563), .A2(new_n647), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n565), .B(new_n648), .C1(new_n594), .C2(new_n603), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n427), .B(new_n649), .C1(new_n321), .C2(new_n334), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n644), .A2(new_n527), .A3(new_n616), .A4(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT37), .B(G110), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  AND3_X1   g467(.A1(new_n525), .A2(KEYINPUT32), .A3(new_n526), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT32), .B1(new_n525), .B2(new_n526), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n649), .B1(new_n656), .B2(new_n515), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n428), .ZN(new_n658));
  INV_X1    g472(.A(new_n639), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n318), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n316), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n658), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n189), .ZN(G30));
  XNOR2_X1  g479(.A(new_n662), .B(KEYINPUT39), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n605), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n667), .B(KEYINPUT40), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n624), .B(KEYINPUT38), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n332), .A2(new_n336), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n243), .A2(new_n312), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n670), .A2(new_n648), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n519), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n507), .A2(new_n487), .A3(new_n509), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n229), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(G472), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n656), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n668), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G143), .ZN(G45));
  NOR2_X1   g496(.A1(new_n632), .A2(new_n663), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n658), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(new_n264), .ZN(G48));
  OAI21_X1  g500(.A(G469), .B1(new_n602), .B2(G902), .ZN(new_n687));
  INV_X1    g501(.A(G469), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n585), .A2(KEYINPUT12), .A3(new_n575), .ZN(new_n689));
  AOI21_X1  g503(.A(KEYINPUT12), .B1(new_n585), .B2(new_n575), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n600), .A2(new_n591), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n591), .B1(new_n600), .B2(new_n582), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n688), .B(new_n229), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n687), .A2(new_n695), .A3(new_n565), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT101), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n687), .A2(new_n695), .A3(new_n698), .A4(new_n565), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n634), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n531), .A2(new_n564), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT102), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT41), .B(G113), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NOR2_X1   g519(.A1(new_n700), .A2(new_n640), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n531), .A2(new_n564), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  NAND4_X1  g522(.A1(new_n648), .A2(new_n687), .A3(new_n695), .A4(new_n565), .ZN(new_n709));
  AOI211_X1 g523(.A(new_n709), .B(new_n427), .C1(new_n321), .C2(new_n334), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n531), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  NOR2_X1   g526(.A1(new_n425), .A2(new_n426), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n713), .A2(new_n674), .A3(new_n320), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n511), .A2(new_n487), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n520), .A2(new_n524), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n526), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(G472), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n525), .B2(new_n229), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n564), .B(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n700), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n714), .A2(new_n721), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  INV_X1    g540(.A(new_n648), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n718), .A2(new_n720), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n427), .A2(new_n696), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(KEYINPUT104), .A3(new_n683), .A4(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT104), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n609), .A2(G472), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n683), .A3(new_n648), .A4(new_n717), .ZN(new_n733));
  INV_X1    g547(.A(new_n729), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  NAND3_X1  g551(.A1(new_n605), .A2(new_n336), .A3(new_n713), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n531), .A2(new_n739), .A3(new_n564), .A4(new_n683), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT42), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n564), .B(KEYINPUT103), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n656), .B2(new_n515), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n738), .A2(new_n741), .A3(new_n684), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n740), .A2(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n282), .ZN(G33));
  NOR2_X1   g560(.A1(new_n659), .A2(new_n663), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n531), .A2(new_n739), .A3(new_n564), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  NAND2_X1  g563(.A1(new_n333), .A2(new_n631), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n750), .B1(KEYINPUT106), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n752), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n617), .A2(new_n648), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(KEYINPUT44), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n565), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n580), .B1(new_n691), .B2(new_n576), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(KEYINPUT45), .A3(new_n583), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(KEYINPUT105), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT45), .B1(new_n760), .B2(new_n583), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n762), .A2(new_n688), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(KEYINPUT105), .B2(new_n761), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT46), .B1(new_n765), .B2(new_n593), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n603), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(KEYINPUT46), .A3(new_n593), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n759), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n666), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n713), .A2(new_n336), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n755), .B2(KEYINPUT44), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n758), .B(new_n774), .C1(new_n773), .C2(new_n772), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  AND2_X1   g590(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n777));
  NOR2_X1   g591(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n769), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n777), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n769), .A2(new_n781), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n531), .A2(new_n564), .A3(new_n684), .A4(new_n771), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  OR2_X1    g599(.A1(new_n696), .A2(new_n336), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n669), .B1(KEYINPUT116), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n787), .B1(KEYINPUT116), .B2(new_n786), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n754), .A2(new_n317), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n723), .A3(new_n721), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT50), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n792), .A2(KEYINPUT117), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(KEYINPUT117), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n771), .A2(new_n696), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n789), .A2(new_n728), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n564), .A3(new_n317), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n680), .A2(new_n797), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n332), .A2(new_n631), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n796), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n793), .A2(new_n794), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n780), .A2(new_n782), .ZN(new_n802));
  INV_X1    g616(.A(new_n687), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n603), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n759), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n790), .A2(new_n771), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n802), .A2(new_n805), .B1(KEYINPUT114), .B2(new_n807), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n807), .A2(KEYINPUT114), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n801), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n657), .B(new_n428), .C1(new_n747), .C2(new_n683), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n674), .A2(new_n713), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n648), .A2(new_n663), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n680), .A2(new_n605), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n816), .A2(new_n736), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n816), .A2(new_n736), .A3(KEYINPUT52), .A4(new_n819), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT110), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n659), .A2(new_n632), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n826), .A2(new_n325), .A3(new_n428), .ZN(new_n827));
  INV_X1    g641(.A(new_n618), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n616), .A2(new_n615), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n651), .A2(new_n606), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n825), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n615), .A2(new_n827), .A3(new_n616), .A4(new_n828), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(KEYINPUT110), .A3(new_n606), .A4(new_n651), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n740), .A2(new_n741), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n743), .A2(new_n744), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n702), .A2(new_n707), .A3(new_n725), .A4(new_n711), .ZN(new_n838));
  OR3_X1    g652(.A1(new_n733), .A2(KEYINPUT111), .A3(new_n738), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT111), .B1(new_n733), .B2(new_n738), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n771), .A2(new_n313), .A3(new_n663), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n531), .A2(new_n842), .A3(new_n605), .A4(new_n648), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n748), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n837), .A2(new_n838), .A3(new_n841), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n824), .A2(new_n834), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n847), .B(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n849), .A2(KEYINPUT54), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n850), .A2(KEYINPUT112), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(KEYINPUT112), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n837), .A2(new_n838), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n702), .A2(new_n707), .A3(new_n725), .A4(new_n711), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT113), .B1(new_n745), .B2(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n822), .A2(new_n823), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n841), .A2(new_n844), .A3(KEYINPUT53), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n831), .B2(new_n833), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n847), .A2(new_n848), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n861), .A2(KEYINPUT54), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n851), .A2(new_n852), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n743), .A2(new_n789), .A3(new_n795), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n864), .B(KEYINPUT48), .Z(new_n865));
  OAI221_X1 g679(.A(new_n314), .B1(new_n790), .B2(new_n734), .C1(new_n798), .C2(new_n632), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n792), .ZN(new_n868));
  OR3_X1    g682(.A1(new_n868), .A2(new_n814), .A3(new_n800), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n867), .B1(new_n810), .B2(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n815), .A2(new_n863), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(G952), .A2(G953), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT118), .Z(new_n873));
  XOR2_X1   g687(.A(new_n804), .B(KEYINPUT49), .Z(new_n874));
  NAND3_X1  g688(.A1(new_n723), .A2(new_n565), .A3(new_n336), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n874), .A2(new_n750), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n670), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n871), .A2(new_n873), .B1(new_n680), .B2(new_n877), .ZN(G75));
  NOR2_X1   g692(.A1(new_n246), .A2(G952), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n860), .A2(new_n229), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT56), .B1(new_n881), .B2(G210), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n390), .A2(new_n411), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(new_n409), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT55), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n880), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n882), .A2(new_n885), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n887), .A2(KEYINPUT119), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(KEYINPUT119), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(G51));
  XOR2_X1   g704(.A(new_n860), .B(KEYINPUT54), .Z(new_n891));
  XOR2_X1   g705(.A(new_n593), .B(KEYINPUT57), .Z(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n694), .B2(new_n693), .ZN(new_n894));
  OR3_X1    g708(.A1(new_n860), .A2(new_n229), .A3(new_n765), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n879), .B1(new_n894), .B2(new_n895), .ZN(G54));
  NAND2_X1  g710(.A1(KEYINPUT58), .A2(G475), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT120), .Z(new_n898));
  NAND2_X1  g712(.A1(new_n881), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n330), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n880), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n900), .B2(new_n899), .ZN(G60));
  NAND2_X1  g716(.A1(G478), .A2(G902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT59), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n627), .B1(new_n863), .B2(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n891), .A2(new_n627), .A3(new_n904), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n905), .A2(new_n879), .A3(new_n906), .ZN(G63));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n908));
  XNOR2_X1  g722(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n223), .A2(new_n229), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n908), .B1(new_n860), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n845), .B1(new_n831), .B2(new_n833), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT53), .B1(new_n914), .B2(new_n824), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n854), .A2(new_n856), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n859), .A2(new_n824), .A3(new_n916), .ZN(new_n917));
  OAI211_X1 g731(.A(KEYINPUT122), .B(new_n911), .C1(new_n915), .C2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n646), .ZN(new_n920));
  INV_X1    g734(.A(new_n554), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n913), .A2(new_n921), .A3(new_n918), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n920), .A2(KEYINPUT61), .A3(new_n880), .A4(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n925), .A3(new_n880), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n920), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n925), .B1(new_n922), .B2(new_n880), .ZN(new_n928));
  OAI211_X1 g742(.A(KEYINPUT124), .B(new_n924), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n922), .A2(new_n880), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT123), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n926), .A3(new_n920), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT124), .B1(new_n933), .B2(new_n924), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n923), .B1(new_n930), .B2(new_n934), .ZN(G66));
  NOR3_X1   g749(.A1(new_n319), .A2(new_n407), .A3(new_n246), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n834), .A2(new_n838), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n936), .B1(new_n938), .B2(new_n246), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n883), .B1(G898), .B2(new_n246), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(G69));
  AND2_X1   g755(.A1(new_n816), .A2(new_n736), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n681), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n531), .A2(new_n564), .A3(new_n739), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n666), .A3(new_n826), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n784), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n775), .A2(new_n944), .A3(new_n945), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n478), .A2(new_n470), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n292), .A2(new_n294), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n950), .B(new_n951), .Z(new_n952));
  NAND3_X1  g766(.A1(new_n949), .A2(new_n246), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n660), .B1(new_n952), .B2(new_n578), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n769), .A2(new_n666), .A3(new_n817), .A4(new_n743), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT125), .Z(new_n956));
  NAND4_X1  g770(.A1(new_n775), .A2(new_n784), .A3(new_n942), .A4(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n745), .B1(new_n747), .B2(new_n946), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n959), .A2(new_n246), .ZN(new_n960));
  AOI22_X1  g774(.A1(new_n958), .A2(new_n960), .B1(G227), .B2(G953), .ZN(new_n961));
  OAI221_X1 g775(.A(new_n953), .B1(new_n246), .B2(new_n954), .C1(new_n961), .C2(new_n952), .ZN(G72));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  NAND2_X1  g778(.A1(new_n938), .A2(new_n959), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n957), .B2(new_n965), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n486), .B(new_n481), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n964), .B1(new_n949), .B2(new_n937), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n970), .A2(new_n486), .A3(new_n481), .ZN(new_n971));
  INV_X1    g785(.A(new_n488), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n964), .B1(new_n972), .B2(new_n676), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT127), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n879), .B1(new_n849), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n969), .A2(new_n976), .ZN(G57));
endmodule


