//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G231gat), .A2(G233gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  AND2_X1   g005(.A1(G15gat), .A2(G22gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G15gat), .A2(G22gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G1gat), .ZN(new_n210));
  INV_X1    g009(.A(G8gat), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n211), .B1(new_n209), .B2(new_n210), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n207), .A2(new_n208), .ZN(new_n214));
  OAI22_X1  g013(.A1(new_n212), .A2(new_n213), .B1(KEYINPUT81), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(new_n210), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G8gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n214), .A2(KEYINPUT81), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT21), .ZN(new_n222));
  NAND2_X1  g021(.A1(G71gat), .A2(G78gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT9), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT88), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT88), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n223), .A2(new_n227), .A3(new_n224), .ZN(new_n228));
  XNOR2_X1  g027(.A(G71gat), .B(G78gat), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G64gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G57gat), .ZN(new_n232));
  INV_X1    g031(.A(G57gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G64gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n235), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(G71gat), .A2(G78gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT87), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n221), .B1(new_n222), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G183gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n230), .A2(new_n235), .B1(new_n237), .B2(new_n240), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(KEYINPUT21), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n245), .A2(new_n248), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n205), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n251), .ZN(new_n253));
  INV_X1    g052(.A(new_n205), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(new_n249), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n204), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n252), .A2(new_n255), .A3(new_n204), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n259), .ZN(new_n261));
  INV_X1    g060(.A(new_n258), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n262), .B2(new_n256), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT82), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT17), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT14), .ZN(new_n266));
  INV_X1    g065(.A(G29gat), .ZN(new_n267));
  INV_X1    g066(.A(G36gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(KEYINPUT80), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G29gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n274), .A3(G36gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G43gat), .B(G50gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(KEYINPUT15), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(KEYINPUT15), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT15), .ZN(new_n280));
  INV_X1    g079(.A(G43gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n281), .A2(G50gat), .ZN(new_n282));
  INV_X1    g081(.A(G50gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(G43gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n280), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n279), .A2(new_n285), .A3(new_n271), .A4(new_n275), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n265), .B1(new_n278), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n278), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G85gat), .A2(G92gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT89), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(KEYINPUT89), .A2(G85gat), .A3(G92gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(KEYINPUT7), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT90), .ZN(new_n297));
  AND2_X1   g096(.A1(G85gat), .A2(G92gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT7), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT8), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n302), .B1(G99gat), .B2(G106gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT91), .B(G85gat), .ZN(new_n304));
  INV_X1    g103(.A(G92gat), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n294), .A2(new_n297), .A3(KEYINPUT7), .A4(new_n295), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n301), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  XOR2_X1   g107(.A(G99gat), .B(G106gat), .Z(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n309), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n301), .A2(new_n306), .A3(new_n311), .A4(new_n307), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n310), .A2(KEYINPUT92), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT92), .B1(new_n310), .B2(new_n312), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n291), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(G232gat), .A2(G233gat), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n315), .A2(KEYINPUT93), .B1(KEYINPUT41), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n310), .A2(new_n312), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT92), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n278), .A2(new_n286), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n310), .A2(KEYINPUT92), .A3(new_n312), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT93), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n291), .B(new_n324), .C1(new_n313), .C2(new_n314), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n317), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G190gat), .B(G218gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n327), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n317), .A2(new_n325), .A3(new_n329), .A4(new_n323), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n316), .A2(KEYINPUT41), .ZN(new_n332));
  XNOR2_X1  g131(.A(G134gat), .B(G162gat), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n332), .B(new_n333), .Z(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n328), .A2(new_n334), .A3(new_n330), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n260), .A2(new_n263), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G230gat), .A2(G233gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n310), .A2(new_n246), .A3(new_n312), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n246), .B1(new_n310), .B2(new_n312), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT10), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n246), .A2(KEYINPUT10), .ZN(new_n346));
  NOR3_X1   g145(.A1(new_n313), .A2(new_n314), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n341), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n341), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(new_n343), .B2(new_n344), .ZN(new_n350));
  XNOR2_X1  g149(.A(G120gat), .B(G148gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(G176gat), .B(G204gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n348), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT94), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n348), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n318), .A2(new_n242), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT10), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n359), .A3(new_n342), .ZN(new_n360));
  INV_X1    g159(.A(new_n346), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n320), .A2(new_n322), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n349), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT94), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n357), .A2(new_n350), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n355), .B1(new_n365), .B2(new_n353), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n340), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT95), .ZN(new_n368));
  NAND2_X1  g167(.A1(G226gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(G169gat), .A2(G176gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n371), .A2(KEYINPUT23), .ZN(new_n372));
  INV_X1    g171(.A(G169gat), .ZN(new_n373));
  INV_X1    g172(.A(G176gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G190gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n244), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(KEYINPUT24), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT24), .B1(new_n244), .B2(new_n378), .ZN(new_n382));
  NOR2_X1   g181(.A1(G183gat), .A2(G190gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n377), .B1(new_n385), .B2(KEYINPUT66), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT66), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n381), .B2(new_n384), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n371), .B(KEYINPUT65), .Z(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT23), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n386), .A2(KEYINPUT25), .A3(new_n388), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n371), .A2(KEYINPUT23), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n385), .A2(new_n376), .A3(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT26), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n375), .B1(new_n389), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n398), .B1(new_n397), .B2(new_n371), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT27), .B(G183gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n401));
  OR2_X1    g200(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n402));
  AND4_X1   g201(.A1(new_n378), .A2(new_n400), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n400), .B2(new_n378), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n403), .A2(new_n379), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n396), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n370), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(G197gat), .A2(G204gat), .ZN(new_n411));
  AND2_X1   g210(.A1(G197gat), .A2(G204gat), .ZN(new_n412));
  AND2_X1   g211(.A1(G211gat), .A2(G218gat), .ZN(new_n413));
  OAI22_X1  g212(.A1(new_n411), .A2(new_n412), .B1(new_n413), .B2(KEYINPUT22), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n414), .A2(KEYINPUT73), .ZN(new_n415));
  NOR2_X1   g214(.A1(G211gat), .A2(G218gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n415), .B(new_n417), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n391), .A2(new_n395), .B1(new_n399), .B2(new_n405), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(new_n369), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n420), .A2(KEYINPUT75), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n407), .A2(KEYINPUT75), .A3(new_n370), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n410), .B(new_n418), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(new_n418), .B(KEYINPUT74), .Z(new_n424));
  OAI21_X1  g223(.A(new_n424), .B1(new_n409), .B2(new_n420), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G8gat), .B(G36gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(G64gat), .B(G92gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n427), .A2(KEYINPUT30), .A3(new_n430), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n423), .A2(KEYINPUT30), .A3(new_n425), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT30), .B1(new_n423), .B2(new_n425), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n432), .A2(new_n433), .A3(new_n430), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(G141gat), .B(G148gat), .Z(new_n436));
  INV_X1    g235(.A(G155gat), .ZN(new_n437));
  INV_X1    g236(.A(G162gat), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT2), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G155gat), .B(G162gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT3), .ZN(new_n444));
  XNOR2_X1  g243(.A(G127gat), .B(G134gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(G113gat), .B(G120gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n446), .A2(KEYINPUT1), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n445), .B1(new_n447), .B2(KEYINPUT68), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT68), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n449), .B1(new_n446), .B2(KEYINPUT1), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n449), .B(new_n445), .C1(new_n446), .C2(KEYINPUT1), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT3), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n442), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n444), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n453), .A2(new_n442), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n458), .A2(KEYINPUT4), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(KEYINPUT4), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G225gat), .A2(G233gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n453), .B(new_n442), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n464), .B(KEYINPUT39), .C1(new_n463), .C2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G1gat), .B(G29gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(G85gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT0), .B(G57gat), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n468), .B(new_n469), .Z(new_n470));
  XOR2_X1   g269(.A(KEYINPUT79), .B(KEYINPUT39), .Z(new_n471));
  OAI211_X1 g270(.A(new_n466), .B(new_n470), .C1(new_n464), .C2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n470), .ZN(new_n475));
  OR3_X1    g274(.A1(new_n461), .A2(KEYINPUT5), .A3(new_n463), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n462), .B1(new_n453), .B2(new_n442), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n461), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT76), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n463), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT5), .A4(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(KEYINPUT5), .B(new_n481), .C1(new_n461), .C2(new_n478), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT76), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n477), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n474), .B1(new_n475), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n473), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n435), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n456), .A2(new_n408), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n424), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n418), .A2(new_n408), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n442), .B1(new_n492), .B2(new_n455), .ZN(new_n493));
  OAI211_X1 g292(.A(G228gat), .B(G233gat), .C1(new_n491), .C2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n417), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT29), .B1(new_n495), .B2(new_n414), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n443), .B(new_n496), .C1(new_n495), .C2(new_n414), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n497), .A2(new_n444), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n498), .A2(KEYINPUT78), .ZN(new_n499));
  NAND2_X1  g298(.A1(G228gat), .A2(G233gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n418), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n490), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n498), .A2(KEYINPUT78), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n499), .A2(new_n500), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n494), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G22gat), .ZN(new_n506));
  INV_X1    g305(.A(G22gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n494), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(KEYINPUT77), .A3(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G78gat), .B(G106gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT31), .B(G50gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n509), .B(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n427), .A2(KEYINPUT38), .A3(new_n430), .ZN(new_n514));
  INV_X1    g313(.A(new_n430), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n426), .A2(KEYINPUT37), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT37), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n423), .A2(new_n517), .A3(new_n425), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n515), .B1(new_n519), .B2(KEYINPUT38), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT38), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n409), .A2(new_n424), .A3(new_n420), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n410), .B1(new_n421), .B2(new_n422), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(new_n501), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n518), .B(new_n521), .C1(new_n524), .C2(new_n517), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n514), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT6), .B1(new_n485), .B2(new_n470), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(new_n470), .B2(new_n485), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n486), .A2(KEYINPUT6), .A3(new_n475), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n489), .B(new_n513), .C1(new_n526), .C2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n435), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n513), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT69), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n407), .A2(new_n536), .A3(new_n454), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT69), .B1(new_n419), .B2(new_n453), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n419), .A2(new_n453), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G227gat), .ZN(new_n541));
  INV_X1    g340(.A(G233gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT33), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G15gat), .B(G43gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(G71gat), .B(G99gat), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n545), .B(new_n546), .Z(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT32), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n550), .B1(new_n540), .B2(new_n543), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n551), .B1(new_n544), .B2(new_n548), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT72), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n553), .A2(KEYINPUT72), .A3(new_n554), .ZN(new_n558));
  NOR3_X1   g357(.A1(new_n540), .A2(KEYINPUT34), .A3(new_n543), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT71), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT70), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n540), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n543), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n540), .A2(new_n563), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n561), .A2(new_n562), .B1(new_n567), .B2(KEYINPUT34), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n557), .A2(new_n558), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n561), .A2(new_n562), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(KEYINPUT34), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n572), .A2(KEYINPUT72), .A3(new_n554), .A4(new_n553), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT36), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n569), .A2(new_n573), .A3(KEYINPUT36), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n531), .A2(new_n535), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT35), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n574), .A2(new_n513), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(new_n533), .ZN(new_n581));
  INV_X1    g380(.A(new_n533), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n582), .A2(KEYINPUT35), .A3(new_n574), .A4(new_n513), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT86), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT83), .ZN(new_n586));
  INV_X1    g385(.A(new_n290), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n221), .B1(new_n587), .B2(new_n287), .ZN(new_n588));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n215), .A2(new_n321), .A3(new_n220), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT18), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n586), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n215), .A2(new_n321), .A3(new_n220), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n594), .B1(new_n291), .B2(new_n221), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n595), .A2(KEYINPUT83), .A3(KEYINPUT18), .A4(new_n589), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n221), .A2(new_n278), .A3(new_n286), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(KEYINPUT84), .A3(new_n590), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n589), .B(KEYINPUT13), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT84), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n215), .A2(new_n321), .A3(new_n220), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n598), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n591), .A2(new_n592), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n593), .A2(new_n596), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G197gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT11), .B(G169gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n605), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT85), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n584), .A2(new_n585), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n585), .B1(new_n584), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n368), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT96), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT96), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n618), .B(new_n368), .C1(new_n614), .C2(new_n615), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n530), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g422(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n206), .A2(new_n211), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n620), .A2(new_n435), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT42), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n620), .A2(new_n435), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(G8gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n627), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n630), .A3(new_n631), .ZN(G1325gat));
  AOI21_X1  g431(.A(G15gat), .B1(new_n620), .B2(new_n574), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n576), .A2(new_n577), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(G15gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(KEYINPUT97), .Z(new_n636));
  AOI21_X1  g435(.A(new_n633), .B1(new_n620), .B2(new_n636), .ZN(G1326gat));
  AOI21_X1  g436(.A(new_n507), .B1(new_n620), .B2(new_n534), .ZN(new_n638));
  AOI211_X1 g437(.A(G22gat), .B(new_n513), .C1(new_n617), .C2(new_n619), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT98), .B(KEYINPUT43), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n584), .A2(new_n613), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT86), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n584), .A2(new_n585), .A3(new_n613), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n618), .B1(new_n646), .B2(new_n368), .ZN(new_n647));
  INV_X1    g446(.A(new_n619), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n534), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(G22gat), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n620), .A2(new_n507), .A3(new_n534), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n640), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n642), .A2(new_n652), .ZN(G1327gat));
  INV_X1    g452(.A(new_n338), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n260), .A2(new_n263), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n366), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n646), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n272), .A2(new_n274), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OR3_X1    g460(.A1(new_n659), .A2(new_n530), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(KEYINPUT45), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT45), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n584), .A2(new_n654), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT99), .B(KEYINPUT44), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n605), .B(new_n610), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n584), .A2(new_n654), .ZN(new_n669));
  NOR2_X1   g468(.A1(KEYINPUT99), .A2(KEYINPUT44), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n667), .A2(new_n668), .A3(new_n671), .A4(new_n658), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n672), .A2(new_n530), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n664), .B1(new_n673), .B2(new_n661), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n663), .B1(new_n674), .B2(new_n662), .ZN(G1328gat));
  NOR3_X1   g474(.A1(new_n659), .A2(G36gat), .A3(new_n532), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT46), .ZN(new_n677));
  OAI21_X1  g476(.A(G36gat), .B1(new_n672), .B2(new_n532), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1329gat));
  INV_X1    g478(.A(new_n634), .ZN(new_n680));
  OAI21_X1  g479(.A(G43gat), .B1(new_n672), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n574), .A2(new_n281), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n659), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n683), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n659), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n646), .A2(KEYINPUT100), .A3(new_n654), .A4(new_n658), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n686), .A2(new_n283), .A3(new_n534), .A4(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT48), .ZN(new_n689));
  OAI21_X1  g488(.A(G50gat), .B1(new_n672), .B2(new_n513), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n689), .B1(new_n688), .B2(new_n690), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(G1331gat));
  NAND4_X1  g492(.A1(new_n584), .A2(new_n612), .A3(new_n340), .A4(new_n657), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n530), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT101), .B(G57gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1332gat));
  NOR2_X1   g496(.A1(new_n694), .A2(new_n532), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT49), .B(G64gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n698), .B2(new_n701), .ZN(G1333gat));
  OAI21_X1  g501(.A(G71gat), .B1(new_n694), .B2(new_n680), .ZN(new_n703));
  INV_X1    g502(.A(new_n574), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n704), .A2(G71gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n694), .B2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g506(.A1(new_n694), .A2(new_n513), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g508(.A1(new_n655), .A2(new_n612), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT102), .Z(new_n711));
  NAND2_X1  g510(.A1(new_n665), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT51), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n657), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n621), .A2(new_n304), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n667), .A2(new_n657), .A3(new_n671), .A4(new_n711), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n530), .ZN(new_n718));
  OAI22_X1  g517(.A1(new_n715), .A2(new_n716), .B1(new_n304), .B2(new_n718), .ZN(G1336gat));
  NAND3_X1  g518(.A1(new_n435), .A2(new_n305), .A3(new_n657), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT103), .Z(new_n721));
  NAND2_X1  g520(.A1(new_n714), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G92gat), .B1(new_n717), .B2(new_n532), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT52), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n723), .B2(KEYINPUT104), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n724), .B(new_n726), .ZN(G1337gat));
  OAI21_X1  g526(.A(G99gat), .B1(new_n717), .B2(new_n680), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n704), .A2(G99gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n715), .B2(new_n729), .ZN(G1338gat));
  NOR3_X1   g529(.A1(new_n513), .A2(G106gat), .A3(new_n366), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT105), .Z(new_n732));
  AOI21_X1  g531(.A(KEYINPUT106), .B1(new_n714), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G106gat), .B1(new_n717), .B2(new_n513), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT53), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n733), .A2(new_n737), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1339gat));
  NOR3_X1   g538(.A1(new_n339), .A2(new_n668), .A3(new_n657), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT54), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n363), .A2(KEYINPUT94), .ZN(new_n743));
  AOI211_X1 g542(.A(new_n356), .B(new_n349), .C1(new_n360), .C2(new_n362), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n360), .A2(new_n362), .A3(new_n349), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT107), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n360), .A2(new_n362), .A3(new_n748), .A4(new_n349), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n747), .A2(KEYINPUT54), .A3(new_n348), .A4(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n745), .A2(KEYINPUT55), .A3(new_n353), .A4(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n355), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n348), .A2(new_n749), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n742), .B1(new_n746), .B2(KEYINPUT107), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n354), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT55), .B1(new_n756), .B2(new_n745), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n753), .A2(new_n757), .A3(new_n612), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n600), .B1(new_n598), .B2(new_n602), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n595), .A2(new_n589), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n609), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AND4_X1   g561(.A1(new_n603), .A2(new_n593), .A3(new_n596), .A4(new_n604), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(new_n611), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n743), .A2(new_n744), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n354), .B1(new_n765), .B2(new_n350), .ZN(new_n766));
  OAI211_X1 g565(.A(KEYINPUT108), .B(new_n764), .C1(new_n766), .C2(new_n355), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n595), .A2(new_n589), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n759), .A2(new_n769), .ZN(new_n770));
  OAI22_X1  g569(.A1(new_n605), .A2(new_n610), .B1(new_n770), .B2(new_n609), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n768), .B1(new_n366), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n338), .B1(new_n758), .B2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n336), .A2(new_n337), .A3(new_n764), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n776), .A2(new_n753), .A3(new_n757), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n774), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n655), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n750), .A2(new_n353), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT54), .B1(new_n357), .B2(new_n364), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n668), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n772), .B(new_n767), .C1(new_n785), .C2(new_n753), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n777), .B1(new_n786), .B2(new_n338), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n775), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n741), .B1(new_n780), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT110), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n656), .B1(new_n787), .B2(new_n775), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n778), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT109), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n795), .A3(new_n741), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n790), .A2(new_n513), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT111), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n530), .A2(new_n435), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n790), .A2(new_n800), .A3(new_n796), .A4(new_n513), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n798), .A2(new_n574), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n613), .A3(new_n805), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n806), .A2(KEYINPUT113), .A3(G113gat), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT113), .B1(new_n806), .B2(G113gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n790), .A2(new_n796), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n580), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n799), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n612), .A2(G113gat), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT114), .ZN(new_n813));
  OAI22_X1  g612(.A1(new_n807), .A2(new_n808), .B1(new_n811), .B2(new_n813), .ZN(G1340gat));
  XNOR2_X1  g613(.A(new_n802), .B(KEYINPUT112), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n657), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G120gat), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n366), .A2(G120gat), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n811), .B2(new_n818), .ZN(G1341gat));
  NOR2_X1   g618(.A1(new_n811), .A2(new_n655), .ZN(new_n820));
  XOR2_X1   g619(.A(new_n820), .B(KEYINPUT115), .Z(new_n821));
  INV_X1    g620(.A(G127gat), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n655), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n821), .A2(new_n822), .B1(new_n815), .B2(new_n823), .ZN(G1342gat));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825));
  INV_X1    g624(.A(G134gat), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(new_n815), .B2(new_n654), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n811), .A2(G134gat), .A3(new_n338), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n828), .B(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n825), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n828), .B(KEYINPUT56), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n804), .A2(new_n654), .A3(new_n805), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n832), .B(KEYINPUT116), .C1(new_n833), .C2(new_n826), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n834), .ZN(G1343gat));
  AOI21_X1  g634(.A(new_n795), .B1(new_n794), .B2(new_n741), .ZN(new_n836));
  AOI211_X1 g635(.A(KEYINPUT110), .B(new_n740), .C1(new_n791), .C2(new_n793), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n839), .A3(new_n534), .ZN(new_n840));
  INV_X1    g639(.A(new_n799), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n634), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT118), .B1(new_n782), .B2(new_n783), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n756), .A2(new_n844), .A3(new_n745), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n845), .A3(new_n781), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT119), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n843), .A2(new_n845), .A3(new_n848), .A4(new_n781), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n753), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT120), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(KEYINPUT120), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n613), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n366), .A2(new_n771), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT117), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n654), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n655), .B1(new_n856), .B2(new_n777), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n513), .B1(new_n857), .B2(new_n741), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n840), .B(new_n842), .C1(new_n858), .C2(new_n839), .ZN(new_n859));
  INV_X1    g658(.A(new_n613), .ZN(new_n860));
  OAI21_X1  g659(.A(G141gat), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g660(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n680), .A2(new_n534), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n809), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n863), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n841), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n860), .A2(G141gat), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT122), .Z(new_n870));
  OAI211_X1 g669(.A(new_n861), .B(new_n862), .C1(new_n868), .C2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n868), .A2(new_n870), .ZN(new_n872));
  INV_X1    g671(.A(new_n859), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n668), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n872), .B1(new_n874), .B2(G141gat), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(G1344gat));
  NOR2_X1   g676(.A1(new_n513), .A2(KEYINPUT57), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n368), .A2(new_n860), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n857), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n839), .B1(new_n838), .B2(new_n534), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n883), .A2(G148gat), .A3(new_n657), .A4(new_n842), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n366), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(G148gat), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT59), .B1(new_n873), .B2(new_n657), .ZN(new_n887));
  AOI22_X1  g686(.A1(KEYINPUT59), .A2(new_n886), .B1(new_n887), .B2(G148gat), .ZN(G1345gat));
  NOR2_X1   g687(.A1(new_n868), .A2(new_n655), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT124), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n656), .A2(G155gat), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n890), .A2(G155gat), .B1(new_n859), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(G1346gat));
  NAND3_X1  g692(.A1(new_n873), .A2(G162gat), .A3(new_n654), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n438), .B1(new_n868), .B2(new_n338), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n621), .A2(new_n532), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n798), .A2(new_n574), .A3(new_n801), .A4(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G169gat), .B1(new_n898), .B2(new_n860), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n810), .A2(new_n897), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n373), .A3(new_n668), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1348gat));
  NOR3_X1   g701(.A1(new_n898), .A2(new_n374), .A3(new_n366), .ZN(new_n903));
  AOI21_X1  g702(.A(G176gat), .B1(new_n900), .B2(new_n657), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(G1349gat));
  OAI21_X1  g704(.A(G183gat), .B1(new_n898), .B2(new_n655), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n900), .A2(new_n400), .A3(new_n656), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g708(.A1(new_n900), .A2(new_n378), .A3(new_n654), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n898), .A2(new_n338), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n912), .A3(G190gat), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n911), .B2(G190gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n910), .B1(new_n914), .B2(new_n915), .ZN(G1351gat));
  OAI21_X1  g715(.A(KEYINPUT57), .B1(new_n809), .B2(new_n513), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n857), .A2(new_n880), .ZN(new_n918));
  OAI211_X1 g717(.A(KEYINPUT125), .B(new_n917), .C1(new_n918), .C2(new_n879), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n881), .B2(new_n882), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n634), .A2(new_n621), .A3(new_n532), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G197gat), .B1(new_n923), .B2(new_n860), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n838), .A2(new_n680), .A3(new_n534), .A4(new_n897), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n612), .A2(G197gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(G1352gat));
  OAI21_X1  g726(.A(G204gat), .B1(new_n923), .B2(new_n366), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n925), .A2(G204gat), .A3(new_n366), .ZN(new_n929));
  XNOR2_X1  g728(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n929), .B(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(new_n931), .ZN(G1353gat));
  OR3_X1    g731(.A1(new_n925), .A2(G211gat), .A3(new_n655), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n883), .A2(new_n656), .A3(new_n922), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n934), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT63), .B1(new_n934), .B2(G211gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(G1354gat));
  INV_X1    g736(.A(KEYINPUT127), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n919), .A2(new_n921), .A3(KEYINPUT127), .A4(new_n922), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n654), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G218gat), .ZN(new_n942));
  OR3_X1    g741(.A1(new_n925), .A2(G218gat), .A3(new_n338), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1355gat));
endmodule


