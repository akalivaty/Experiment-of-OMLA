//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n203), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT64), .B(G238), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n202), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n211), .B(new_n217), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT65), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n202), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n239), .B(new_n245), .Z(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n214), .ZN(new_n248));
  OR2_X1    g0048(.A1(new_n248), .A2(KEYINPUT66), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(KEYINPUT66), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(G20), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G50), .A3(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n258));
  INV_X1    g0058(.A(G150), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT8), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(new_n201), .B2(KEYINPUT67), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT67), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(KEYINPUT8), .A3(G58), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n215), .A2(G33), .ZN(new_n267));
  OAI221_X1 g0067(.A(new_n258), .B1(new_n259), .B2(new_n261), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n268), .A2(new_n251), .B1(new_n240), .B2(new_n254), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n257), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT9), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT72), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AND3_X1   g0079(.A1(new_n275), .A2(G226), .A3(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n214), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n278), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT3), .B(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G222), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G77), .ZN(new_n290));
  INV_X1    g0090(.A(G223), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(G1698), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n289), .B1(new_n290), .B2(new_n287), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  AOI211_X1 g0093(.A(new_n280), .B(new_n286), .C1(new_n293), .C2(new_n282), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G190), .ZN(new_n295));
  INV_X1    g0095(.A(G200), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n295), .B1(new_n271), .B2(new_n270), .C1(new_n296), .C2(new_n294), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n273), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g0098(.A(new_n298), .B(KEYINPUT10), .Z(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n270), .B1(new_n294), .B2(G169), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n287), .A2(G20), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT7), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n308), .B(G68), .C1(new_n306), .C2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G58), .A2(G68), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n203), .A2(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n312), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n310), .A2(KEYINPUT16), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n248), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT76), .ZN(new_n316));
  INV_X1    g0116(.A(new_n307), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n306), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G33), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT74), .B1(new_n319), .B2(KEYINPUT3), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT74), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT3), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(new_n322), .A3(G33), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n320), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n309), .A2(G20), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT75), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT75), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n325), .A2(new_n329), .A3(new_n326), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n318), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n316), .B1(new_n331), .B2(new_n202), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n325), .A2(new_n329), .A3(new_n326), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n329), .B1(new_n325), .B2(new_n326), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n333), .A2(new_n334), .B1(new_n306), .B2(new_n317), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(KEYINPUT76), .A3(G68), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n332), .A2(new_n336), .A3(new_n313), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT16), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n315), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G232), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n279), .A2(new_n275), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n285), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n291), .A2(new_n288), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n287), .B(new_n343), .C1(G226), .C2(new_n288), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G87), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n275), .B1(new_n346), .B2(KEYINPUT77), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT77), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n344), .A2(new_n348), .A3(new_n345), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n342), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(G200), .ZN(new_n351));
  AOI211_X1 g0151(.A(G190), .B(new_n342), .C1(new_n347), .C2(new_n349), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n266), .B1(new_n252), .B2(G20), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n255), .A2(new_n354), .B1(new_n254), .B2(new_n266), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n339), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT17), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n350), .A2(G179), .ZN(new_n359));
  INV_X1    g0159(.A(G169), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(new_n360), .B2(new_n350), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n339), .B2(new_n356), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT18), .ZN(new_n363));
  INV_X1    g0163(.A(G190), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n350), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(G200), .B2(new_n350), .ZN(new_n366));
  INV_X1    g0166(.A(new_n313), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n335), .A2(G68), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n367), .B1(new_n368), .B2(new_n316), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT16), .B1(new_n369), .B2(new_n336), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n355), .B(new_n366), .C1(new_n370), .C2(new_n315), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT17), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT18), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n374), .B(new_n361), .C1(new_n339), .C2(new_n356), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n358), .A2(new_n363), .A3(new_n373), .A4(new_n375), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT8), .B(G58), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n377), .A2(new_n261), .B1(new_n215), .B2(new_n290), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT15), .B(G87), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n267), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n248), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT70), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n254), .A2(new_n248), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(G77), .A3(new_n256), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(G77), .B2(new_n253), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G244), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n285), .B1(new_n387), .B2(new_n341), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT68), .ZN(new_n389));
  XNOR2_X1  g0189(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n287), .A2(G232), .A3(new_n288), .ZN(new_n391));
  INV_X1    g0191(.A(G107), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(new_n287), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n292), .A2(new_n218), .ZN(new_n394));
  OR3_X1    g0194(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT69), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT69), .B1(new_n393), .B2(new_n394), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n282), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OAI211_X1 g0199(.A(KEYINPUT71), .B(new_n386), .C1(new_n399), .C2(new_n296), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT71), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n296), .B1(new_n390), .B2(new_n397), .ZN(new_n402));
  INV_X1    g0202(.A(new_n386), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n399), .A2(G190), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n400), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT14), .ZN(new_n407));
  INV_X1    g0207(.A(G238), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n285), .B1(new_n408), .B2(new_n341), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n340), .A2(G1698), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n287), .B(new_n410), .C1(G226), .C2(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G97), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n275), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OR3_X1    g0213(.A1(new_n409), .A2(KEYINPUT13), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT13), .B1(new_n409), .B2(new_n413), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n407), .B1(new_n416), .B2(G169), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n414), .A2(G179), .A3(new_n415), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(new_n407), .A3(G169), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n254), .A2(new_n202), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n422), .B(KEYINPUT12), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n260), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n290), .B2(new_n267), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n251), .A2(KEYINPUT11), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n383), .A2(G68), .A3(new_n256), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT11), .B1(new_n251), .B2(new_n425), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n421), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n430), .B1(new_n416), .B2(new_n364), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n296), .B1(new_n414), .B2(new_n415), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n398), .A2(new_n360), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n390), .A2(new_n397), .A3(new_n300), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(new_n403), .A3(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n406), .A2(new_n432), .A3(new_n436), .A4(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n305), .A2(new_n376), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n322), .A2(G33), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n442), .A2(new_n324), .A3(G238), .A4(new_n288), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n442), .A2(new_n324), .A3(G244), .A4(G1698), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G116), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n282), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n277), .A2(G1), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n275), .A2(G274), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT79), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n252), .A2(G45), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n451), .B(G250), .C1(new_n281), .C2(new_n214), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n450), .B1(new_n449), .B2(new_n452), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n447), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(KEYINPUT80), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT80), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n449), .A2(new_n452), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT79), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n453), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n458), .B1(new_n461), .B2(new_n447), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n360), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n456), .A2(KEYINPUT80), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(new_n458), .A3(new_n447), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n300), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n287), .A2(new_n215), .A3(G68), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT19), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n215), .B1(new_n412), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(G87), .B2(new_n206), .ZN(new_n470));
  INV_X1    g0270(.A(G97), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n267), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n467), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n248), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n379), .A2(new_n254), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n252), .A2(G33), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n249), .A2(new_n253), .A3(new_n250), .A4(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n474), .B(new_n475), .C1(new_n379), .C2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n463), .A2(new_n466), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(G200), .B1(new_n457), .B2(new_n462), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n464), .A2(G190), .A3(new_n465), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n474), .A2(new_n475), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT81), .ZN(new_n483));
  INV_X1    g0283(.A(G87), .ZN(new_n484));
  OR3_X1    g0284(.A1(new_n477), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n477), .B2(new_n484), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n480), .A2(new_n481), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n479), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT82), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n322), .A2(G33), .ZN(new_n493));
  OAI21_X1  g0293(.A(G303), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n442), .A2(new_n324), .A3(G264), .A4(G1698), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n442), .A2(new_n324), .A3(G257), .A4(new_n288), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n282), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT83), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n497), .A2(KEYINPUT83), .A3(new_n282), .ZN(new_n501));
  XNOR2_X1  g0301(.A(KEYINPUT5), .B(G41), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n282), .B1(new_n448), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n502), .A2(new_n448), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n503), .A2(G270), .B1(new_n504), .B2(new_n284), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n500), .A2(new_n501), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G283), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n507), .B(new_n215), .C1(G33), .C2(new_n471), .ZN(new_n508));
  INV_X1    g0308(.A(G116), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G20), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n248), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT20), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(G13), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n510), .A2(G1), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n509), .B1(new_n252), .B2(G33), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(new_n383), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n360), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n506), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT21), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n506), .A2(new_n518), .A3(KEYINPUT21), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n505), .A2(new_n501), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n513), .A2(new_n517), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n523), .A2(G179), .A3(new_n524), .A4(new_n500), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n521), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n524), .B1(new_n506), .B2(G200), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT84), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n506), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n527), .A2(new_n528), .B1(G190), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n526), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n479), .A2(new_n488), .A3(KEYINPUT82), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n335), .A2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n392), .A2(KEYINPUT6), .A3(G97), .ZN(new_n535));
  XOR2_X1   g0335(.A(G97), .B(G107), .Z(new_n536));
  OAI21_X1  g0336(.A(new_n535), .B1(new_n536), .B2(KEYINPUT6), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n537), .A2(G20), .B1(G77), .B2(new_n260), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n248), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n477), .A2(new_n471), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n253), .A2(G97), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n287), .A2(G250), .A3(G1698), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n287), .A2(G244), .A3(new_n288), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT4), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n507), .B(new_n544), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n282), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND4_X1   g0349(.A1(G274), .A2(new_n502), .A3(new_n275), .A4(new_n448), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n503), .A2(G257), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(KEYINPUT78), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT78), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n503), .A2(new_n553), .A3(G257), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n549), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G200), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n549), .A2(new_n552), .A3(G190), .A4(new_n554), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n540), .A2(new_n543), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n555), .A2(new_n360), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n549), .A2(new_n552), .A3(new_n300), .A4(new_n554), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n534), .A2(new_n538), .B1(new_n214), .B2(new_n247), .ZN(new_n561));
  INV_X1    g0361(.A(new_n543), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n559), .B(new_n560), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n491), .A2(new_n532), .A3(new_n533), .A4(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT87), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n442), .A2(new_n324), .A3(G257), .A4(G1698), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n442), .A2(new_n324), .A3(G250), .A4(new_n288), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G33), .A2(G294), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n282), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n503), .A2(G264), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n566), .B1(new_n573), .B2(new_n550), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n282), .A2(new_n570), .B1(new_n503), .B2(G264), .ZN(new_n575));
  INV_X1    g0375(.A(new_n550), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(KEYINPUT87), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n364), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT89), .ZN(new_n579));
  OR2_X1    g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT88), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n573), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n575), .A2(KEYINPUT88), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n576), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n578), .A2(new_n579), .B1(new_n584), .B2(new_n296), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n442), .A2(new_n324), .A3(new_n215), .A4(G87), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT22), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT22), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n287), .A2(new_n589), .A3(new_n215), .A4(G87), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n445), .A2(G20), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT23), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n215), .B2(G107), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n392), .A2(KEYINPUT23), .A3(G20), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT24), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(KEYINPUT85), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n596), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n588), .B2(new_n590), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT85), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT24), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n597), .A2(KEYINPUT85), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n248), .B(new_n599), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n253), .A2(G107), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n606), .B(KEYINPUT25), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n477), .B2(new_n392), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT86), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n607), .B(KEYINPUT86), .C1(new_n477), .C2(new_n392), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n586), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n577), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT87), .B1(new_n575), .B2(new_n576), .ZN(new_n617));
  OAI21_X1  g0417(.A(G169), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n582), .A2(new_n583), .A3(G179), .A4(new_n576), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n613), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n565), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n441), .A2(new_n623), .ZN(G372));
  INV_X1    g0424(.A(new_n563), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n491), .A2(KEYINPUT26), .A3(new_n533), .A4(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n456), .A2(G200), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n481), .A2(new_n487), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n456), .A2(new_n360), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n466), .A2(new_n478), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n627), .B1(new_n632), .B2(new_n563), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT90), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(KEYINPUT90), .B(new_n627), .C1(new_n632), .C2(new_n563), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n626), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n631), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n558), .A2(new_n563), .A3(new_n631), .A4(new_n629), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n613), .B1(new_n580), .B2(new_n585), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n526), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n621), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n638), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n441), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT91), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n355), .B1(new_n370), .B2(new_n315), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n374), .B1(new_n648), .B2(new_n361), .ZN(new_n649));
  INV_X1    g0449(.A(new_n375), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n363), .A2(KEYINPUT91), .A3(new_n375), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n358), .A2(new_n373), .ZN(new_n654));
  INV_X1    g0454(.A(new_n439), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n436), .A2(new_n655), .B1(new_n421), .B2(new_n431), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n653), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n303), .B1(new_n657), .B2(new_n299), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n646), .A2(new_n658), .ZN(G369));
  NAND3_X1  g0459(.A1(new_n252), .A2(new_n215), .A3(G13), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT92), .ZN(new_n662));
  INV_X1    g0462(.A(G213), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n660), .B2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n524), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n642), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n532), .B2(new_n668), .ZN(new_n670));
  INV_X1    g0470(.A(G330), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n618), .A2(new_n619), .B1(new_n605), .B2(new_n612), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n640), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n667), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n614), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n667), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n642), .A2(new_n667), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n674), .A2(new_n680), .B1(new_n673), .B2(new_n675), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(G399));
  INV_X1    g0482(.A(KEYINPUT93), .ZN(new_n683));
  INV_X1    g0483(.A(new_n209), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n683), .B1(new_n684), .B2(G41), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n209), .A2(KEYINPUT93), .A3(new_n276), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n212), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n639), .A2(new_n640), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT97), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n642), .A2(new_n621), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT97), .B1(new_n673), .B2(new_n526), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n631), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n632), .A2(new_n563), .A3(new_n627), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n491), .A2(new_n533), .A3(new_n625), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n627), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n675), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT29), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n667), .B1(new_n637), .B2(new_n644), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n702), .B1(KEYINPUT29), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT96), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n457), .A2(new_n462), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n500), .A2(G179), .A3(new_n501), .A4(new_n505), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT94), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n582), .A2(new_n583), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n549), .A2(new_n552), .A3(new_n554), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n708), .A2(new_n710), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n709), .A2(KEYINPUT94), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n707), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n464), .A2(new_n465), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n582), .A2(new_n583), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n716), .A2(new_n717), .A3(new_n555), .ZN(new_n718));
  INV_X1    g0518(.A(new_n714), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n719), .A4(new_n710), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n584), .A2(new_n555), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT95), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n584), .A2(KEYINPUT95), .A3(new_n555), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n506), .A2(new_n300), .A3(new_n456), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n715), .A2(new_n720), .A3(new_n726), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT31), .B1(new_n727), .B2(new_n667), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n706), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n727), .A2(new_n667), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(KEYINPUT96), .A3(new_n734), .ZN(new_n735));
  OR3_X1    g0535(.A1(new_n565), .A2(new_n622), .A3(new_n667), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n730), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n705), .B1(G330), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n691), .B1(new_n738), .B2(G1), .ZN(G364));
  XNOR2_X1  g0539(.A(new_n672), .B(KEYINPUT98), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n514), .A2(G20), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G45), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(KEYINPUT99), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n252), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(KEYINPUT99), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n687), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n670), .B2(new_n671), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n740), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n215), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT100), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n670), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n748), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n214), .B1(G20), .B2(new_n360), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n215), .A2(G179), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(new_n364), .A3(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n392), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n215), .A2(new_n300), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n763), .A2(new_n296), .A3(G190), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n759), .A2(G190), .A3(G200), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n765), .A2(new_n202), .B1(new_n766), .B2(new_n484), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n763), .A2(new_n364), .A3(new_n296), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n761), .B(new_n767), .C1(G50), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n296), .A2(G190), .ZN(new_n770));
  OAI21_X1  g0570(.A(G20), .B1(new_n770), .B2(G179), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT101), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G97), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G190), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n759), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT32), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n763), .A2(new_n770), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n287), .B1(new_n785), .B2(new_n201), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n762), .A2(new_n779), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n786), .B1(G77), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n769), .A2(new_n778), .A3(new_n783), .A4(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G322), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n785), .A2(new_n791), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n780), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n287), .B(new_n793), .C1(G329), .C2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n768), .ZN(new_n796));
  INV_X1    g0596(.A(G326), .ZN(new_n797));
  INV_X1    g0597(.A(G303), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n796), .A2(new_n797), .B1(new_n766), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(KEYINPUT33), .B(G317), .Z(new_n800));
  INV_X1    g0600(.A(G283), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n765), .A2(new_n800), .B1(new_n760), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G294), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n795), .B(new_n803), .C1(new_n804), .C2(new_n776), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n758), .B1(new_n790), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n754), .A2(new_n757), .ZN(new_n807));
  NAND3_X1  g0607(.A1(G355), .A2(new_n287), .A3(new_n209), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n245), .A2(new_n277), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n684), .A2(new_n287), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(G45), .B2(new_n212), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n808), .B1(G116), .B2(new_n209), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n756), .B(new_n806), .C1(new_n807), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n755), .A2(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n750), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  NAND2_X1  g0616(.A1(new_n439), .A2(KEYINPUT105), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT105), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n437), .A2(new_n818), .A3(new_n403), .A4(new_n438), .ZN(new_n819));
  AND3_X1   g0619(.A1(new_n406), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n645), .A2(new_n675), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n403), .A2(new_n667), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n406), .A2(new_n817), .A3(new_n822), .A4(new_n819), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n655), .A2(new_n667), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n821), .B1(new_n703), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n737), .A2(G330), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n748), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n827), .B2(new_n826), .ZN(new_n829));
  INV_X1    g0629(.A(new_n751), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n758), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n748), .B1(G77), .B2(new_n831), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n785), .A2(new_n804), .B1(new_n787), .B2(new_n509), .ZN(new_n833));
  INV_X1    g0633(.A(new_n760), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(G87), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n835), .B1(new_n796), .B2(new_n798), .C1(new_n801), .C2(new_n765), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n833), .B(new_n836), .C1(G311), .C2(new_n794), .ZN(new_n837));
  INV_X1    g0637(.A(new_n287), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n766), .B2(new_n392), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT102), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n837), .A2(new_n778), .A3(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G143), .A2(new_n784), .B1(new_n788), .B2(G159), .ZN(new_n842));
  INV_X1    g0642(.A(G137), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n842), .B1(new_n796), .B2(new_n843), .C1(new_n259), .C2(new_n765), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT34), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(KEYINPUT103), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n760), .A2(new_n202), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n838), .B1(new_n794), .B2(G132), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n240), .B2(new_n766), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n847), .B(new_n849), .C1(new_n777), .C2(G58), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n845), .A2(KEYINPUT103), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n841), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n832), .B1(new_n853), .B2(new_n757), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT104), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n830), .B2(new_n825), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n829), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  NAND2_X1  g0658(.A1(new_n314), .A2(new_n251), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT16), .B1(new_n310), .B2(new_n313), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n355), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n665), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT107), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n863), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n376), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n361), .A2(new_n861), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT108), .B1(new_n371), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(new_n865), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n371), .A2(KEYINPUT108), .A3(new_n868), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n862), .B1(new_n339), .B2(new_n356), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n362), .A2(new_n873), .A3(new_n371), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n874), .A2(KEYINPUT37), .ZN(new_n875));
  OAI211_X1 g0675(.A(KEYINPUT38), .B(new_n866), .C1(new_n872), .C2(new_n875), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n874), .B(new_n867), .ZN(new_n877));
  INV_X1    g0677(.A(new_n654), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n363), .A2(KEYINPUT91), .A3(new_n375), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT91), .B1(new_n363), .B2(new_n375), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n873), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n877), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n876), .B1(new_n883), .B2(KEYINPUT38), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n728), .A2(new_n729), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n736), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n431), .A2(new_n667), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n432), .A2(new_n436), .A3(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n431), .B(new_n667), .C1(new_n421), .C2(new_n435), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n890), .A2(new_n825), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n886), .A2(new_n891), .A3(KEYINPUT40), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT109), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n884), .A2(new_n892), .A3(KEYINPUT109), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT40), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT108), .ZN(new_n899));
  INV_X1    g0699(.A(new_n868), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n899), .B1(new_n357), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n863), .B(KEYINPUT107), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n871), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n875), .B1(new_n903), .B2(KEYINPUT37), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n376), .A2(new_n865), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n898), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n876), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n886), .A2(new_n891), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n895), .A2(new_n896), .B1(new_n897), .B2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n441), .A2(new_n886), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n910), .A2(new_n911), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n913), .A2(new_n671), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n873), .B1(new_n653), .B2(new_n878), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n898), .B1(new_n916), .B2(new_n877), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT39), .B1(new_n917), .B2(new_n876), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n906), .A2(new_n876), .A3(KEYINPUT39), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n421), .A2(new_n431), .A3(new_n675), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n667), .B1(new_n817), .B2(new_n819), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT106), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n703), .B2(new_n820), .ZN(new_n924));
  INV_X1    g0724(.A(new_n890), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n907), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n653), .B2(new_n862), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n705), .A2(new_n441), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n658), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n915), .A2(new_n932), .B1(new_n252), .B2(new_n741), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n932), .B2(new_n915), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n537), .A2(KEYINPUT35), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n537), .A2(KEYINPUT35), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n935), .A2(G116), .A3(new_n216), .A4(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT36), .Z(new_n938));
  NAND3_X1  g0738(.A1(new_n213), .A2(G77), .A3(new_n311), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n252), .B(G13), .C1(new_n939), .C2(new_n241), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n934), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT110), .Z(G367));
  OAI21_X1  g0742(.A(new_n807), .B1(new_n209), .B2(new_n379), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n235), .A2(new_n810), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n748), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n287), .B1(new_n788), .B2(G283), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n768), .A2(G311), .B1(G97), .B2(new_n834), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n784), .A2(G303), .B1(new_n794), .B2(G317), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n764), .A2(G294), .ZN(new_n949));
  AND4_X1   g0749(.A1(new_n946), .A2(new_n947), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n766), .ZN(new_n951));
  OAI21_X1  g0751(.A(G116), .B1(KEYINPUT114), .B2(KEYINPUT46), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(KEYINPUT114), .A2(KEYINPUT46), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n954), .B1(new_n951), .B2(new_n953), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n950), .B1(new_n392), .B2(new_n776), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT115), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n785), .A2(new_n259), .B1(new_n787), .B2(new_n240), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n838), .B(new_n959), .C1(G137), .C2(new_n794), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n777), .A2(G68), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n760), .A2(new_n290), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n764), .B2(G159), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n768), .A2(G143), .B1(G58), .B2(new_n951), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n960), .A2(new_n961), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n958), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT47), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n945), .B1(new_n967), .B2(new_n757), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n487), .A2(new_n675), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n632), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n638), .A2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n754), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n968), .A2(new_n974), .ZN(new_n975));
  OR3_X1    g0775(.A1(new_n563), .A2(KEYINPUT111), .A3(new_n675), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT111), .B1(new_n563), .B2(new_n675), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n667), .B1(new_n561), .B2(new_n562), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n564), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n674), .A3(new_n680), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT42), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n978), .A2(KEYINPUT112), .A3(new_n980), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT112), .B1(new_n978), .B2(new_n980), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n673), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n667), .B1(new_n986), .B2(new_n563), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT43), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n988), .A2(new_n989), .A3(new_n973), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n973), .A2(new_n989), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n991), .B(new_n992), .C1(new_n983), .C2(new_n987), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n984), .A2(new_n985), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n995), .A2(new_n679), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(KEYINPUT113), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n994), .A2(new_n997), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT113), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n990), .A2(new_n993), .A3(new_n1000), .A4(new_n996), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n674), .A2(new_n680), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n678), .B2(new_n680), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n1004), .A2(new_n671), .A3(new_n670), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n740), .B2(new_n1004), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n705), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1006), .A2(new_n1007), .A3(new_n827), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n681), .A2(new_n981), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(KEYINPUT44), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT44), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n681), .A2(new_n981), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n681), .A2(new_n981), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT45), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT45), .B1(new_n681), .B2(new_n981), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n1010), .A2(new_n1012), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n679), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n738), .B1(new_n1008), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n687), .B(KEYINPUT41), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n746), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n975), .B1(new_n1002), .B2(new_n1023), .ZN(G387));
  NAND2_X1  g0824(.A1(new_n1008), .A2(new_n747), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT117), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OR3_X1    g0827(.A1(new_n738), .A2(KEYINPUT118), .A3(new_n1006), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1008), .A2(KEYINPUT117), .A3(new_n747), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT118), .B1(new_n738), .B2(new_n1006), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1006), .A2(new_n746), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n838), .B1(new_n780), .B2(new_n797), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G317), .A2(new_n784), .B1(new_n788), .B2(G303), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n796), .B2(new_n791), .C1(new_n792), .C2(new_n765), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n777), .A2(G283), .B1(G294), .B2(new_n951), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT49), .Z(new_n1041));
  AOI211_X1 g0841(.A(new_n1033), .B(new_n1041), .C1(G116), .C2(new_n834), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n784), .A2(G50), .B1(new_n794), .B2(G150), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1043), .B(new_n287), .C1(new_n202), .C2(new_n787), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n776), .A2(new_n379), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n796), .A2(new_n781), .B1(new_n760), .B2(new_n471), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n765), .A2(new_n266), .B1(new_n766), .B2(new_n290), .ZN(new_n1047));
  NOR4_X1   g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n757), .B1(new_n1042), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n232), .A2(G45), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n377), .A2(G50), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT50), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n277), .B1(new_n202), .B2(new_n290), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n688), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT116), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1052), .B(new_n1056), .C1(new_n1055), .C2(new_n1054), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1050), .A2(new_n810), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n287), .A2(new_n209), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1058), .B1(G107), .B2(new_n209), .C1(new_n688), .C2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n756), .B1(new_n1060), .B2(new_n807), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1049), .B(new_n1061), .C1(new_n678), .C2(new_n753), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1032), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1031), .A2(new_n1063), .ZN(G393));
  INV_X1    g0864(.A(new_n1008), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1019), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n687), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n1008), .A2(new_n1019), .A3(KEYINPUT120), .ZN(new_n1068));
  AOI21_X1  g0868(.A(KEYINPUT120), .B1(new_n1008), .B2(new_n1019), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n239), .A2(new_n810), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n807), .B1(new_n471), .B2(new_n209), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n768), .A2(G317), .B1(new_n784), .B2(G311), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT119), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT52), .Z(new_n1075));
  OAI221_X1 g0875(.A(new_n838), .B1(new_n780), .B2(new_n791), .C1(new_n804), .C2(new_n787), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n761), .B1(new_n764), .B2(G303), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n801), .B2(new_n766), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1076), .B(new_n1078), .C1(G116), .C2(new_n777), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n768), .A2(G150), .B1(new_n784), .B2(G159), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT51), .Z(new_n1081));
  INV_X1    g0881(.A(G143), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n287), .B1(new_n780), .B2(new_n1082), .C1(new_n377), .C2(new_n787), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n835), .B1(new_n202), .B2(new_n766), .C1(new_n765), .C2(new_n240), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(G77), .C2(new_n777), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1075), .A2(new_n1079), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n748), .B1(new_n1071), .B2(new_n1072), .C1(new_n1086), .C2(new_n758), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n995), .B2(new_n754), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n1066), .B2(new_n746), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1070), .A2(new_n1089), .ZN(G390));
  AND3_X1   g0890(.A1(new_n886), .A2(new_n891), .A3(G330), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n920), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n922), .B(KEYINPUT106), .Z(new_n1093));
  NAND2_X1  g0893(.A1(new_n821), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1092), .B1(new_n1094), .B2(new_n890), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT39), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n884), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n906), .A2(new_n876), .A3(KEYINPUT39), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n675), .B(new_n820), .C1(new_n697), .C2(new_n700), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n1093), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1092), .B1(new_n1101), .B2(new_n890), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n884), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1091), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n918), .A2(new_n919), .B1(new_n1092), .B2(new_n926), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n737), .A2(G330), .A3(new_n891), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n1107), .A3(new_n1103), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n733), .A2(new_n734), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n565), .A2(new_n622), .A3(new_n667), .ZN(new_n1111));
  OAI211_X1 g0911(.A(G330), .B(new_n825), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n925), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1100), .A2(new_n1093), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1107), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT121), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1107), .A2(new_n1113), .A3(new_n1114), .A4(KEYINPUT121), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n737), .A2(G330), .A3(new_n825), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1091), .B1(new_n925), .B2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1117), .B(new_n1118), .C1(new_n924), .C2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n441), .A2(G330), .A3(new_n886), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n930), .A2(new_n658), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1109), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1105), .A2(new_n1108), .A3(new_n1121), .A4(new_n1124), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n747), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1105), .A2(new_n1108), .A3(new_n746), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n751), .B1(new_n918), .B2(new_n919), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n392), .A2(new_n765), .B1(new_n796), .B2(new_n801), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n847), .B(new_n1131), .C1(G87), .C2(new_n951), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n785), .A2(new_n509), .B1(new_n787), .B2(new_n471), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n287), .B(new_n1133), .C1(G294), .C2(new_n794), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1132), .B(new_n1134), .C1(new_n290), .C2(new_n776), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n838), .B1(new_n794), .B2(G125), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n240), .B2(new_n760), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT122), .Z(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G132), .A2(new_n784), .B1(new_n788), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(G128), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(new_n1142), .B2(new_n796), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G137), .B2(new_n764), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n766), .A2(new_n259), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT53), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(new_n781), .C2(new_n776), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1135), .B1(new_n1138), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n757), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n758), .A2(new_n266), .A3(new_n830), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1130), .A2(new_n748), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1128), .A2(new_n1129), .A3(new_n1151), .ZN(G378));
  AOI21_X1  g0952(.A(new_n671), .B1(new_n909), .B2(new_n897), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n270), .A2(new_n862), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n299), .A2(new_n304), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1154), .B1(new_n299), .B2(new_n304), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  OR3_X1    g0958(.A1(new_n1155), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1158), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n896), .ZN(new_n1162));
  AOI21_X1  g0962(.A(KEYINPUT109), .B1(new_n884), .B2(new_n892), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1153), .B(new_n1161), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n895), .A2(new_n896), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1161), .B1(new_n1166), .B2(new_n1153), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n1165), .A2(new_n1167), .B1(new_n921), .B2(new_n928), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1153), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1161), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1171), .A2(new_n929), .A3(new_n1164), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n746), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1170), .A2(new_n751), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n748), .B1(G50), .B2(new_n831), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n240), .B1(G33), .B2(G41), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n838), .B2(new_n276), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n785), .A2(new_n392), .B1(new_n379), .B2(new_n787), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n838), .B(new_n276), .C1(new_n801), .C2(new_n780), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n760), .A2(new_n201), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G77), .B2(new_n951), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n764), .A2(G97), .B1(new_n768), .B2(G116), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n961), .A2(new_n1181), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1178), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n785), .A2(new_n1142), .B1(new_n787), .B2(new_n843), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G132), .B2(new_n764), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n768), .A2(G125), .B1(new_n951), .B2(new_n1140), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n259), .C2(new_n776), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n834), .A2(G159), .ZN(new_n1193));
  AOI211_X1 g0993(.A(G33), .B(G41), .C1(new_n794), .C2(G124), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1187), .B1(new_n1186), .B2(new_n1185), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1176), .B1(new_n1197), .B2(new_n757), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1175), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1174), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1127), .A2(new_n1124), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1171), .A2(new_n929), .A3(new_n1164), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n929), .B1(new_n1171), .B2(new_n1164), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1201), .B(KEYINPUT57), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1204), .A2(new_n747), .ZN(new_n1205));
  AOI21_X1  g1005(.A(KEYINPUT57), .B1(new_n1173), .B2(new_n1201), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1200), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(G375));
  NAND2_X1  g1009(.A1(new_n1119), .A2(new_n925), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1091), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1094), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1213), .A2(new_n1117), .A3(new_n1118), .A4(new_n1123), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1125), .A2(new_n1022), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n925), .A2(new_n751), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n748), .B1(G68), .B2(new_n831), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n765), .A2(new_n1139), .B1(new_n781), .B2(new_n766), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1182), .B(new_n1218), .C1(G132), .C2(new_n768), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n787), .A2(new_n259), .B1(new_n780), .B2(new_n1142), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n838), .B(new_n1220), .C1(G137), .C2(new_n784), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(new_n240), .C2(new_n776), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n785), .A2(new_n801), .B1(new_n787), .B2(new_n392), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n287), .B(new_n1223), .C1(G303), .C2(new_n794), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n962), .B1(new_n764), .B2(G116), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n768), .A2(G294), .B1(G97), .B2(new_n951), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1222), .B1(new_n1045), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1217), .B1(new_n1228), .B2(new_n757), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1121), .A2(new_n746), .B1(new_n1216), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1215), .A2(new_n1230), .ZN(G381));
  NAND3_X1  g1031(.A1(new_n1070), .A2(new_n857), .A3(new_n1089), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1232), .A2(G387), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1031), .A2(new_n815), .A3(new_n1063), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(new_n1233), .A2(G378), .A3(G381), .A4(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1208), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT123), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1236), .B(new_n1237), .ZN(G407));
  INV_X1    g1038(.A(G378), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n663), .A2(G343), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT124), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n663), .B1(new_n1208), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(G407), .A2(KEYINPUT125), .A3(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT123), .B1(new_n1235), .B2(new_n1208), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1243), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT125), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1244), .A2(new_n1249), .ZN(G409));
  INV_X1    g1050(.A(new_n1234), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1070), .A2(new_n1089), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n815), .B1(new_n1031), .B2(new_n1063), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G393), .A2(G396), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G390), .B1(new_n1255), .B2(new_n1234), .ZN(new_n1256));
  OAI21_X1  g1056(.A(G387), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1252), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1258));
  INV_X1    g1058(.A(G387), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1255), .A2(G390), .A3(new_n1234), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1257), .A2(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT127), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1173), .A2(new_n746), .B1(new_n1175), .B2(new_n1198), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1204), .A2(new_n747), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G378), .B(new_n1264), .C1(new_n1265), .C2(new_n1206), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1201), .B(new_n1022), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1174), .A2(new_n1267), .A3(new_n1199), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1239), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1240), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1214), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n747), .A3(new_n1125), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1121), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT126), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1275), .A2(new_n1276), .A3(KEYINPUT60), .A4(new_n1123), .ZN(new_n1277));
  OAI21_X1  g1077(.A(KEYINPUT126), .B1(new_n1214), .B2(new_n1272), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1274), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1230), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n857), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1274), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1284), .A2(G384), .A3(new_n1230), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1270), .A2(new_n1271), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1241), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n1288), .A2(new_n1289), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1241), .A2(G2897), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1240), .A2(G2897), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1295), .B1(new_n1287), .B2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1293), .B1(new_n1298), .B2(new_n1290), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1263), .B1(new_n1292), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1286), .A2(new_n1296), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1301), .B1(new_n1295), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1288), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1290), .A2(KEYINPUT63), .A3(new_n1287), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1262), .A2(KEYINPUT61), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1303), .A2(new_n1305), .A3(new_n1306), .A4(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1300), .A2(new_n1308), .ZN(G405));
  NAND2_X1  g1109(.A1(G375), .A2(new_n1239), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(new_n1266), .A3(new_n1286), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1208), .A2(G378), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1266), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1287), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1311), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1262), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1311), .A2(new_n1314), .A3(new_n1261), .A4(new_n1257), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(G402));
endmodule


