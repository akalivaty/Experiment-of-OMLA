//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  INV_X1    g004(.A(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(KEYINPUT26), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT71), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(G169gat), .A3(G176gat), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n212), .A2(new_n214), .B1(new_n207), .B2(KEYINPUT26), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n204), .B1(new_n210), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT28), .ZN(new_n218));
  NOR2_X1   g017(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n219));
  INV_X1    g018(.A(G183gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT69), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT69), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G183gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n219), .B1(new_n224), .B2(KEYINPUT27), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n218), .B1(new_n225), .B2(G190gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT27), .B(G183gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n218), .A2(G190gat), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n226), .A2(KEYINPUT70), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n219), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT69), .B(G183gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT27), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G190gat), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT28), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n217), .B1(new_n229), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT23), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n212), .A2(new_n214), .B1(new_n207), .B2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT23), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(KEYINPUT25), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT68), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n245), .B1(new_n231), .B2(new_n234), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n242), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n212), .A2(new_n214), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n207), .A2(new_n239), .ZN(new_n251));
  NOR2_X1   g050(.A1(G169gat), .A2(G176gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n249), .A2(new_n250), .A3(new_n251), .A4(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n240), .A2(KEYINPUT67), .A3(new_n249), .A4(new_n253), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n245), .B1(new_n220), .B2(new_n234), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n243), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n259), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n256), .A2(new_n257), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT25), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n247), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G113gat), .B(G120gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(KEYINPUT1), .ZN(new_n267));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n268), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n270), .B1(KEYINPUT1), .B2(new_n266), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n238), .A2(new_n265), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n269), .A2(new_n271), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n263), .A2(new_n264), .ZN(new_n275));
  INV_X1    g074(.A(new_n247), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n208), .B(KEYINPUT71), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n278), .A2(new_n215), .B1(G183gat), .B2(G190gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n227), .A2(new_n228), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n280), .B1(new_n235), .B2(new_n236), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n226), .A2(KEYINPUT70), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n279), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n274), .B1(new_n277), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n203), .B1(new_n273), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT32), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT33), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(G15gat), .B(G43gat), .Z(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT72), .ZN(new_n290));
  XNOR2_X1  g089(.A(G71gat), .B(G99gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT73), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n290), .B(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n286), .A2(new_n288), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n272), .B1(new_n238), .B2(new_n265), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n274), .A3(new_n283), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n202), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n293), .B1(new_n297), .B2(KEYINPUT33), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT32), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT34), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n295), .A2(new_n296), .A3(new_n303), .A4(new_n202), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT75), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n295), .A2(new_n296), .A3(new_n202), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT34), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n304), .A2(new_n305), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT74), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n302), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n273), .A2(new_n284), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n313), .A2(KEYINPUT75), .A3(new_n303), .A4(new_n202), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(new_n308), .A3(new_n306), .ZN(new_n315));
  AOI22_X1  g114(.A1(KEYINPUT74), .A2(new_n315), .B1(new_n294), .B2(new_n301), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT36), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n306), .A2(new_n308), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n294), .A2(new_n318), .A3(new_n301), .A4(new_n314), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n298), .A2(new_n300), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n295), .A2(new_n296), .ZN(new_n321));
  AOI221_X4 g120(.A(new_n299), .B1(KEYINPUT33), .B2(new_n293), .C1(new_n321), .C2(new_n203), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n315), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n317), .A2(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(G8gat), .B(G36gat), .Z(new_n328));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(new_n238), .B2(new_n265), .ZN(new_n333));
  XOR2_X1   g132(.A(G211gat), .B(G218gat), .Z(new_n334));
  XNOR2_X1  g133(.A(G197gat), .B(G204gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT22), .ZN(new_n336));
  INV_X1    g135(.A(G211gat), .ZN(new_n337));
  INV_X1    g136(.A(G218gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n334), .B1(new_n341), .B2(KEYINPUT77), .ZN(new_n342));
  INV_X1    g141(.A(new_n334), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n344), .A3(new_n340), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT29), .B1(new_n277), .B2(new_n283), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n333), .B(new_n346), .C1(new_n347), .C2(new_n332), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n350), .B1(new_n238), .B2(new_n265), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n331), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n346), .B1(new_n352), .B2(new_n333), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n330), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT30), .ZN(new_n355));
  INV_X1    g154(.A(new_n346), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n347), .A2(new_n332), .ZN(new_n357));
  INV_X1    g156(.A(new_n333), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n348), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT30), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n361), .A3(new_n330), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(G1gat), .B(G29gat), .Z(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(KEYINPUT0), .ZN(new_n365));
  XNOR2_X1  g164(.A(G57gat), .B(G85gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT81), .ZN(new_n370));
  INV_X1    g169(.A(G148gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G141gat), .ZN(new_n372));
  INV_X1    g171(.A(G141gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G148gat), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT80), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G155gat), .B(G162gat), .ZN(new_n376));
  INV_X1    g175(.A(G155gat), .ZN(new_n377));
  INV_X1    g176(.A(G162gat), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT2), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n375), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n376), .B1(new_n375), .B2(new_n379), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(new_n274), .ZN(new_n384));
  INV_X1    g183(.A(new_n382), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n385), .A2(new_n380), .A3(new_n269), .A4(new_n271), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n370), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT5), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT3), .B1(new_n381), .B2(new_n382), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n385), .A2(new_n391), .A3(new_n380), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n392), .A3(new_n272), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n383), .A2(new_n274), .A3(KEYINPUT4), .ZN(new_n396));
  INV_X1    g195(.A(new_n370), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n393), .A2(new_n395), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n389), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT5), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n368), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(KEYINPUT6), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n401), .A3(new_n368), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AND4_X1   g204(.A1(KEYINPUT6), .A2(new_n399), .A3(new_n401), .A4(new_n368), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n349), .B2(new_n353), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n359), .A2(KEYINPUT78), .A3(new_n348), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n330), .B(KEYINPUT79), .Z(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n363), .A2(new_n408), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n342), .A2(new_n350), .A3(new_n345), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n383), .B1(new_n415), .B2(new_n391), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n392), .A2(new_n350), .B1(new_n345), .B2(new_n342), .ZN(new_n417));
  NAND2_X1  g216(.A1(G228gat), .A2(G233gat), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT82), .B1(new_n335), .B2(new_n339), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n335), .A2(KEYINPUT82), .A3(new_n339), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n334), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT29), .B1(new_n420), .B2(new_n343), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n391), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT83), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n385), .A2(new_n380), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n417), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT3), .B1(new_n423), .B2(new_n424), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT83), .B1(new_n431), .B2(new_n383), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n419), .B1(new_n433), .B2(new_n418), .ZN(new_n434));
  OR2_X1    g233(.A1(KEYINPUT84), .A2(G22gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(KEYINPUT84), .A2(G22gat), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(G78gat), .B(G106gat), .Z(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT31), .B(G50gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n437), .B(new_n440), .C1(new_n434), .C2(new_n435), .ZN(new_n441));
  INV_X1    g240(.A(G22gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(KEYINPUT85), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n440), .B1(new_n434), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(new_n434), .B2(new_n444), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n414), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n441), .A2(new_n446), .ZN(new_n449));
  NOR3_X1   g248(.A1(new_n349), .A2(new_n353), .A3(new_n409), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT78), .B1(new_n359), .B2(new_n348), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n452), .A2(new_n412), .B1(new_n355), .B2(new_n362), .ZN(new_n453));
  INV_X1    g252(.A(new_n404), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n370), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n384), .A2(new_n387), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n456), .B(KEYINPUT39), .C1(new_n370), .C2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT39), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n455), .A2(new_n459), .A3(new_n370), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n460), .A2(new_n461), .A3(new_n367), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n461), .B1(new_n460), .B2(new_n367), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n458), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT40), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n454), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(KEYINPUT40), .B(new_n458), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n467), .A2(KEYINPUT87), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(KEYINPUT87), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n449), .B1(new_n453), .B2(new_n470), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n454), .A2(new_n402), .A3(KEYINPUT6), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(new_n406), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n349), .B2(new_n353), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n359), .A2(KEYINPUT37), .A3(new_n348), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT38), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .A4(new_n412), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n478), .A3(new_n354), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT37), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n330), .B1(new_n360), .B2(new_n474), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n327), .B(new_n448), .C1(new_n471), .C2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n449), .B1(new_n312), .B2(new_n316), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT35), .B1(new_n485), .B2(new_n414), .ZN(new_n486));
  INV_X1    g285(.A(new_n324), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n447), .A2(KEYINPUT35), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n487), .A2(new_n488), .A3(new_n408), .A4(new_n453), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G229gat), .A2(G233gat), .ZN(new_n492));
  XOR2_X1   g291(.A(new_n492), .B(KEYINPUT13), .Z(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G43gat), .B(G50gat), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n495), .A2(KEYINPUT15), .ZN(new_n496));
  NOR3_X1   g295(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(G29gat), .A2(G36gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n495), .A2(KEYINPUT15), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n496), .A2(new_n500), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT89), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n497), .B1(new_n504), .B2(new_n499), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n504), .B2(new_n499), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n502), .B1(new_n506), .B2(new_n501), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT90), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n507), .A2(new_n508), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT91), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n507), .B(new_n508), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n514), .A3(new_n503), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G15gat), .B(G22gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT16), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(G1gat), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(G1gat), .B2(new_n517), .ZN(new_n520));
  INV_X1    g319(.A(G8gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n522), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n512), .A2(new_n515), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n494), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT92), .B(KEYINPUT17), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n515), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n513), .A2(KEYINPUT17), .A3(new_n503), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n530), .A3(new_n522), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(new_n492), .A3(new_n525), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT18), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n526), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n531), .A2(KEYINPUT18), .A3(new_n492), .A4(new_n525), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G113gat), .B(G141gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT88), .B(G197gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(KEYINPUT11), .B(G169gat), .Z(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT12), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n536), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n534), .A2(new_n535), .A3(new_n542), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(G71gat), .A2(G78gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G57gat), .B(G64gat), .Z(new_n550));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(KEYINPUT9), .B2(new_n547), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n552), .B(new_n553), .Z(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(KEYINPUT21), .ZN(new_n556));
  NAND2_X1  g355(.A1(G231gat), .A2(G233gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G127gat), .B(G155gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT20), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n558), .B(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n524), .B1(KEYINPUT21), .B2(new_n555), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n562), .B(KEYINPUT95), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n561), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G183gat), .B(G211gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n564), .B(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G190gat), .B(G218gat), .Z(new_n569));
  NAND2_X1  g368(.A1(G85gat), .A2(G92gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT7), .ZN(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  INV_X1    g371(.A(G85gat), .ZN(new_n573));
  INV_X1    g372(.A(G92gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(KEYINPUT8), .A2(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G99gat), .B(G106gat), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n576), .B(KEYINPUT96), .ZN(new_n581));
  INV_X1    g380(.A(new_n579), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n529), .A2(new_n530), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT41), .ZN(new_n588));
  NAND2_X1  g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589));
  OAI22_X1  g388(.A1(new_n516), .A2(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n569), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n588), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  NOR2_X1   g393(.A1(new_n589), .A2(new_n588), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n512), .A2(new_n515), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n595), .B1(new_n596), .B2(new_n584), .ZN(new_n597));
  INV_X1    g396(.A(new_n569), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n598), .A3(new_n586), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n591), .A2(new_n594), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n594), .B1(new_n591), .B2(new_n599), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n568), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n584), .A2(new_n555), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT97), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n580), .A2(new_n583), .A3(new_n554), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n585), .A2(KEYINPUT97), .A3(new_n554), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT10), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n604), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n604), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n608), .A2(new_n614), .A3(new_n609), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n615), .A2(new_n622), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n623), .A2(new_n613), .A3(new_n619), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n491), .A2(new_n546), .A3(new_n603), .A4(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(new_n408), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(G1gat), .Z(G1324gat));
  INV_X1    g429(.A(new_n628), .ZN(new_n631));
  INV_X1    g430(.A(new_n453), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n521), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT16), .B(G8gat), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n628), .A2(new_n453), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT42), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n636), .B1(KEYINPUT42), .B2(new_n635), .ZN(G1325gat));
  OAI21_X1  g436(.A(G15gat), .B1(new_n628), .B2(new_n327), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n324), .A2(G15gat), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n638), .B1(new_n628), .B2(new_n639), .ZN(G1326gat));
  NOR2_X1   g439(.A1(new_n628), .A2(new_n449), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT43), .B(G22gat), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(G1327gat));
  INV_X1    g442(.A(new_n568), .ZN(new_n644));
  INV_X1    g443(.A(new_n545), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n542), .B1(new_n534), .B2(new_n535), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n644), .A2(new_n647), .A3(new_n626), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n600), .A2(new_n601), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n484), .B2(new_n490), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n654), .A2(G29gat), .A3(new_n408), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n655), .B(KEYINPUT45), .Z(new_n656));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n491), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n484), .A2(new_n490), .A3(KEYINPUT99), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n602), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n658), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n652), .A2(KEYINPUT44), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n649), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(G29gat), .B1(new_n666), .B2(new_n408), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n656), .A2(new_n667), .ZN(G1328gat));
  NOR3_X1   g467(.A1(new_n654), .A2(G36gat), .A3(new_n453), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT100), .B(KEYINPUT46), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(G36gat), .B1(new_n666), .B2(new_n453), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(G1329gat));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT101), .B(KEYINPUT47), .Z(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n324), .A2(G43gat), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n648), .A2(new_n651), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n327), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n484), .A2(new_n490), .A3(KEYINPUT99), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT99), .B1(new_n484), .B2(new_n490), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n681), .A2(new_n682), .A3(new_n661), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n651), .A2(new_n660), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n680), .B(new_n648), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G43gat), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n679), .B1(new_n686), .B2(KEYINPUT102), .ZN(new_n687));
  INV_X1    g486(.A(G43gat), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(new_n665), .B2(new_n680), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n676), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT47), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n686), .B2(new_n695), .ZN(new_n696));
  AOI211_X1 g495(.A(KEYINPUT103), .B(new_n694), .C1(new_n685), .C2(G43gat), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n674), .B1(new_n692), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n678), .B1(new_n689), .B2(new_n690), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n686), .A2(KEYINPUT102), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n675), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT103), .B1(new_n689), .B2(new_n694), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n686), .A2(new_n693), .A3(new_n695), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n702), .A2(KEYINPUT104), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n699), .A2(new_n706), .ZN(G1330gat));
  OAI21_X1  g506(.A(G50gat), .B1(new_n666), .B2(new_n449), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n654), .A2(G50gat), .A3(new_n449), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT48), .B1(new_n709), .B2(KEYINPUT105), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1331gat));
  INV_X1    g511(.A(new_n603), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n546), .A2(new_n627), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR4_X1   g514(.A1(new_n681), .A2(new_n682), .A3(new_n713), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n473), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n632), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT49), .B(G64gat), .Z(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n719), .B2(new_n721), .ZN(G1333gat));
  AND2_X1   g521(.A1(new_n716), .A2(new_n487), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n723), .A2(G71gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n716), .A2(G71gat), .A3(new_n680), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(KEYINPUT106), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(KEYINPUT106), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n724), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g528(.A1(new_n716), .A2(new_n447), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT107), .B(G78gat), .Z(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1335gat));
  NAND3_X1  g531(.A1(new_n651), .A2(new_n647), .A3(new_n568), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT51), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n626), .B1(new_n734), .B2(KEYINPUT108), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n735), .B1(KEYINPUT108), .B2(new_n734), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(new_n573), .A3(new_n473), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n663), .A2(new_n664), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n715), .A2(new_n644), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741), .B2(new_n408), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n737), .A2(new_n742), .ZN(G1336gat));
  NOR2_X1   g542(.A1(new_n734), .A2(new_n627), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n574), .A3(new_n632), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n746));
  NAND2_X1  g545(.A1(new_n740), .A2(new_n632), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G92gat), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n747), .A2(new_n748), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n745), .B(new_n746), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n745), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n574), .B1(new_n740), .B2(new_n632), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT52), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(G1337gat));
  INV_X1    g555(.A(G99gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n736), .A2(new_n757), .A3(new_n487), .ZN(new_n758));
  OAI21_X1  g557(.A(G99gat), .B1(new_n741), .B2(new_n327), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(G1338gat));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761));
  INV_X1    g560(.A(G106gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n744), .A2(new_n762), .A3(new_n447), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n740), .A2(new_n447), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT111), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G106gat), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n764), .A2(KEYINPUT111), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n761), .B(new_n763), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n763), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n762), .B1(new_n740), .B2(new_n447), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT53), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(G1339gat));
  NAND3_X1  g571(.A1(new_n603), .A2(new_n647), .A3(new_n627), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n492), .B1(new_n531), .B2(new_n525), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n523), .A2(new_n525), .A3(new_n494), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n541), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n626), .A2(new_n545), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n608), .A2(new_n609), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n611), .ZN(new_n780));
  INV_X1    g579(.A(new_n612), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n780), .A2(new_n614), .A3(new_n781), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n782), .A2(KEYINPUT54), .A3(new_n613), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n620), .B1(new_n613), .B2(KEYINPUT54), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n778), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n614), .B1(new_n780), .B2(new_n781), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n619), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n782), .A2(KEYINPUT54), .A3(new_n613), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(KEYINPUT55), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n785), .A2(new_n625), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n777), .B1(new_n791), .B2(new_n647), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n650), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n545), .A2(new_n776), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n792), .A2(new_n650), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n773), .B1(new_n795), .B2(new_n644), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n797), .A2(new_n408), .A3(new_n485), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(new_n453), .ZN(new_n799));
  INV_X1    g598(.A(G113gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n800), .A3(new_n546), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n449), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n324), .B1(new_n802), .B2(KEYINPUT112), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n453), .A2(new_n473), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n796), .A2(new_n806), .A3(new_n449), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n803), .A2(new_n546), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n808), .A2(KEYINPUT113), .A3(G113gat), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT113), .B1(new_n808), .B2(G113gat), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n801), .B1(new_n809), .B2(new_n810), .ZN(G1340gat));
  INV_X1    g610(.A(G120gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n799), .A2(new_n812), .A3(new_n626), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n803), .A2(new_n626), .A3(new_n805), .A4(new_n807), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n814), .A2(new_n815), .A3(G120gat), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n814), .B2(G120gat), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n813), .B1(new_n816), .B2(new_n817), .ZN(G1341gat));
  INV_X1    g617(.A(G127gat), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n799), .A2(new_n819), .A3(new_n644), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n803), .A2(new_n805), .A3(new_n807), .ZN(new_n821));
  OAI21_X1  g620(.A(G127gat), .B1(new_n821), .B2(new_n568), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(G1342gat));
  INV_X1    g622(.A(G134gat), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n602), .A2(new_n453), .ZN(new_n825));
  XOR2_X1   g624(.A(new_n825), .B(KEYINPUT115), .Z(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n798), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT56), .Z(new_n829));
  OAI21_X1  g628(.A(G134gat), .B1(new_n821), .B2(new_n650), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(G1343gat));
  INV_X1    g630(.A(new_n625), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n788), .A2(new_n789), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n833), .B2(new_n778), .ZN(new_n834));
  AND4_X1   g633(.A1(new_n602), .A2(new_n834), .A3(new_n790), .A4(new_n794), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n792), .A2(new_n650), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n834), .A2(new_n546), .A3(new_n790), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n602), .B1(new_n839), .B2(new_n777), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT117), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n644), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n773), .ZN(new_n843));
  OAI211_X1 g642(.A(KEYINPUT57), .B(new_n447), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g643(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n845), .B1(new_n797), .B2(new_n449), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n680), .A2(new_n804), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G141gat), .B1(new_n849), .B2(new_n647), .ZN(new_n850));
  NAND2_X1  g649(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n797), .A2(new_n408), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n680), .A2(new_n449), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n453), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n647), .A2(G141gat), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT119), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n850), .A2(new_n851), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n859), .ZN(new_n861));
  INV_X1    g660(.A(new_n848), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n862), .B1(new_n844), .B2(new_n846), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n373), .B1(new_n863), .B2(new_n546), .ZN(new_n864));
  INV_X1    g663(.A(new_n856), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n851), .B1(new_n854), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n861), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n860), .A2(new_n867), .ZN(G1344gat));
  NAND3_X1  g667(.A1(new_n855), .A2(new_n371), .A3(new_n626), .ZN(new_n869));
  AOI211_X1 g668(.A(KEYINPUT59), .B(new_n371), .C1(new_n863), .C2(new_n626), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871));
  INV_X1    g670(.A(new_n845), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n796), .A2(new_n447), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n568), .B1(new_n840), .B2(new_n835), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n449), .B1(new_n874), .B2(new_n773), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n873), .B1(KEYINPUT57), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n626), .A3(new_n848), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n871), .B1(new_n877), .B2(G148gat), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n869), .B1(new_n870), .B2(new_n878), .ZN(G1345gat));
  OAI21_X1  g678(.A(G155gat), .B1(new_n849), .B2(new_n568), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n855), .A2(new_n377), .A3(new_n644), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1346gat));
  OAI21_X1  g681(.A(G162gat), .B1(new_n849), .B2(new_n650), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n852), .A2(new_n853), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n827), .A2(new_n378), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(G1347gat));
  NAND2_X1  g685(.A1(new_n632), .A2(new_n408), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT120), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n803), .A2(new_n807), .A3(new_n888), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(new_n205), .A3(new_n647), .ZN(new_n890));
  NOR4_X1   g689(.A1(new_n797), .A2(new_n473), .A3(new_n453), .A4(new_n485), .ZN(new_n891));
  AOI21_X1  g690(.A(G169gat), .B1(new_n891), .B2(new_n546), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n890), .A2(new_n892), .ZN(G1348gat));
  OAI21_X1  g692(.A(G176gat), .B1(new_n889), .B2(new_n627), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n891), .A2(new_n206), .A3(new_n626), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT121), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n894), .A2(new_n898), .A3(new_n895), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1349gat));
  OAI21_X1  g699(.A(new_n224), .B1(new_n889), .B2(new_n568), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n891), .A2(new_n227), .A3(new_n644), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT60), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n901), .A2(new_n905), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1350gat));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n234), .A3(new_n602), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n803), .A2(new_n602), .A3(new_n807), .A4(new_n888), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n910));
  AND4_X1   g709(.A1(KEYINPUT122), .A2(new_n909), .A3(new_n910), .A4(G190gat), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n234), .B1(new_n912), .B2(KEYINPUT61), .ZN(new_n913));
  AOI22_X1  g712(.A1(new_n909), .A2(new_n913), .B1(KEYINPUT122), .B2(new_n910), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n908), .B1(new_n911), .B2(new_n914), .ZN(G1351gat));
  NAND4_X1  g714(.A1(new_n796), .A2(new_n408), .A3(new_n632), .A4(new_n853), .ZN(new_n916));
  OR3_X1    g715(.A1(new_n916), .A2(G197gat), .A3(new_n647), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n888), .A2(new_n327), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n876), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n546), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT123), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G197gat), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n920), .A2(KEYINPUT123), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n917), .B1(new_n922), .B2(new_n923), .ZN(G1352gat));
  NAND2_X1  g723(.A1(new_n919), .A2(new_n626), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(G204gat), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n916), .A2(G204gat), .A3(new_n627), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT62), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(G1353gat));
  INV_X1    g728(.A(new_n916), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n337), .A3(new_n644), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT63), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n932), .A2(KEYINPUT125), .ZN(new_n933));
  AOI211_X1 g732(.A(new_n449), .B(new_n845), .C1(new_n874), .C2(new_n773), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT57), .B1(new_n796), .B2(new_n447), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n644), .B(new_n918), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT124), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n876), .A2(new_n938), .A3(new_n644), .A4(new_n918), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n337), .B1(KEYINPUT125), .B2(new_n932), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n933), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n933), .ZN(new_n943));
  INV_X1    g742(.A(new_n941), .ZN(new_n944));
  AOI211_X1 g743(.A(new_n943), .B(new_n944), .C1(new_n937), .C2(new_n939), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n931), .B1(new_n942), .B2(new_n945), .ZN(G1354gat));
  NOR3_X1   g745(.A1(new_n916), .A2(G218gat), .A3(new_n650), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n919), .A2(new_n602), .ZN(new_n949));
  OAI211_X1 g748(.A(KEYINPUT126), .B(new_n948), .C1(new_n949), .C2(new_n338), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n338), .B1(new_n919), .B2(new_n602), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(new_n947), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(new_n953), .ZN(G1355gat));
endmodule


