//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n214, new_n215,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298;
  INV_X1    g0000(.A(KEYINPUT65), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G50), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(G58), .A2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n201), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT64), .B(G50), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n211), .A2(KEYINPUT65), .A3(new_n207), .ZN(new_n212));
  AND3_X1   g0012(.A1(new_n209), .A2(new_n210), .A3(new_n212), .ZN(G353));
  NOR2_X1   g0013(.A1(G97), .A2(G107), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G87), .ZN(G355));
  INV_X1    g0016(.A(G1), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT0), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n208), .A2(G50), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n218), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n229));
  INV_X1    g0029(.A(G58), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  INV_X1    g0031(.A(G97), .ZN(new_n232));
  INV_X1    g0032(.A(G257), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n229), .B1(new_n230), .B2(new_n231), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  AOI22_X1  g0034(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n235));
  AOI22_X1  g0035(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g0037(.A(new_n220), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  OAI211_X1 g0038(.A(new_n223), .B(new_n228), .C1(KEYINPUT1), .C2(new_n238), .ZN(new_n239));
  AOI21_X1  g0039(.A(new_n239), .B1(KEYINPUT1), .B2(new_n238), .ZN(G361));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n231), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT66), .ZN(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G68), .B(G77), .Z(new_n253));
  XOR2_X1   g0053(.A(G50), .B(G58), .Z(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  INV_X1    g0056(.A(KEYINPUT10), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(new_n262), .A3(G274), .ZN(new_n263));
  INV_X1    g0063(.A(new_n262), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n260), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G226), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n263), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  OR2_X1    g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT67), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n273), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(G223), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n275), .A2(new_n276), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G1698), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n281), .A2(G222), .B1(new_n280), .B2(G77), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n268), .B1(new_n283), .B2(new_n264), .ZN(new_n284));
  INV_X1    g0084(.A(G200), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n257), .B1(new_n286), .B2(KEYINPUT72), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n226), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT68), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n218), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n230), .A2(KEYINPUT8), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT8), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G58), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G150), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n290), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT8), .B(G58), .ZN(new_n300));
  OAI211_X1 g0100(.A(KEYINPUT68), .B(new_n297), .C1(new_n300), .C2(new_n291), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n218), .B1(new_n209), .B2(new_n212), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n289), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n217), .A2(G20), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G50), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT71), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n217), .A2(G13), .A3(G20), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT69), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT69), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n310), .A2(new_n217), .A3(G13), .A4(G20), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n289), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT70), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT70), .ZN(new_n315));
  AOI211_X1 g0115(.A(new_n315), .B(new_n289), .C1(new_n309), .C2(new_n311), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n307), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n309), .A2(new_n311), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n202), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n304), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT9), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n320), .A2(new_n321), .B1(new_n284), .B2(G190), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n304), .A2(KEYINPUT9), .A3(new_n317), .A4(new_n319), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT72), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(KEYINPUT73), .A3(KEYINPUT10), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n287), .A2(new_n322), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n320), .A2(new_n321), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n284), .A2(G190), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n286), .B1(new_n329), .B2(KEYINPUT73), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n326), .B1(new_n330), .B2(new_n257), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n284), .A2(G169), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n284), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n320), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g0136(.A(G223), .B(new_n269), .C1(new_n275), .C2(new_n276), .ZN(new_n337));
  OAI211_X1 g0137(.A(G226), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G33), .A2(G87), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n264), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n217), .B1(G41), .B2(G45), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n262), .A2(G232), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n263), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT76), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT76), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n263), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n341), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n285), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n263), .A2(new_n343), .A3(new_n346), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n346), .B1(new_n263), .B2(new_n343), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G190), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(new_n353), .A3(new_n341), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  INV_X1    g0156(.A(G68), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT3), .B(G33), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n359), .B2(G20), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n280), .A2(KEYINPUT7), .A3(new_n218), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n230), .A2(new_n357), .ZN(new_n363));
  OAI21_X1  g0163(.A(G20), .B1(new_n363), .B2(new_n207), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n296), .A2(G159), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n356), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT7), .B1(new_n280), .B2(new_n218), .ZN(new_n368));
  NOR4_X1   g0168(.A1(new_n275), .A2(new_n276), .A3(new_n358), .A4(G20), .ZN(new_n369));
  OAI21_X1  g0169(.A(G68), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n366), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(KEYINPUT16), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n367), .A2(new_n372), .A3(new_n289), .ZN(new_n373));
  INV_X1    g0173(.A(new_n305), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n300), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n314), .B2(new_n316), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n318), .A2(new_n300), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n355), .A2(KEYINPUT77), .A3(new_n373), .A4(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT17), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n376), .A2(new_n377), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n370), .A2(new_n371), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n313), .B1(new_n383), .B2(new_n356), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n382), .B1(new_n384), .B2(new_n372), .ZN(new_n385));
  INV_X1    g0185(.A(G169), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n348), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(G179), .B2(new_n348), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT18), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n385), .A2(KEYINPUT77), .A3(KEYINPUT17), .A4(new_n355), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n378), .A2(new_n373), .ZN(new_n391));
  AOI21_X1  g0191(.A(G169), .B1(new_n352), .B2(new_n341), .ZN(new_n392));
  AND4_X1   g0192(.A1(new_n333), .A2(new_n341), .A3(new_n345), .A4(new_n347), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT18), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n391), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n381), .A2(new_n389), .A3(new_n390), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n312), .A2(new_n313), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n398), .A2(new_n210), .A3(new_n374), .ZN(new_n399));
  INV_X1    g0199(.A(new_n300), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n400), .A2(new_n296), .B1(G20), .B2(G77), .ZN(new_n401));
  XNOR2_X1  g0201(.A(KEYINPUT15), .B(G87), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G33), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(G20), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n313), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n312), .A2(G77), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n399), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n263), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(G244), .B2(new_n265), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n359), .A2(G232), .A3(new_n269), .ZN(new_n412));
  INV_X1    g0212(.A(G107), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(new_n359), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT67), .B1(new_n280), .B2(new_n269), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n277), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n416), .B2(G238), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n411), .B1(new_n417), .B2(new_n262), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n409), .B1(new_n418), .B2(new_n386), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(G179), .B2(new_n418), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n418), .A2(G200), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n409), .B1(new_n418), .B2(new_n353), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n397), .A2(new_n423), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n405), .A2(G77), .B1(G20), .B2(new_n357), .ZN(new_n425));
  INV_X1    g0225(.A(new_n296), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n425), .B1(new_n202), .B2(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n427), .A2(KEYINPUT11), .A3(new_n289), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT11), .B1(new_n427), .B2(new_n289), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT12), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n318), .A2(new_n431), .A3(new_n357), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT12), .B1(new_n312), .B2(G68), .ZN(new_n433));
  INV_X1    g0233(.A(new_n398), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n374), .A2(new_n357), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n432), .A2(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT75), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n430), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n432), .A2(new_n433), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(new_n435), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n439), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT13), .ZN(new_n445));
  OAI211_X1 g0245(.A(G232), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n446));
  OAI211_X1 g0246(.A(G226), .B(new_n269), .C1(new_n275), .C2(new_n276), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G97), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n264), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT74), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT74), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n452), .A3(new_n264), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n410), .B1(G238), .B2(new_n265), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n445), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n449), .A2(new_n452), .A3(new_n264), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n452), .B1(new_n449), .B2(new_n264), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n445), .B(new_n455), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n444), .B(G169), .C1(new_n456), .C2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT13), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(G179), .A3(new_n459), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n459), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n444), .B1(new_n466), .B2(G169), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n443), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n463), .A2(G190), .A3(new_n459), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n442), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n285), .B1(new_n463), .B2(new_n459), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n336), .A2(new_n424), .A3(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G244), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n476));
  OAI211_X1 g0276(.A(G238), .B(new_n269), .C1(new_n275), .C2(new_n276), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n476), .B(new_n477), .C1(new_n404), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n264), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n217), .A2(G45), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(new_n262), .A3(G274), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n262), .A2(G250), .A3(new_n481), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT79), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT79), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n480), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(new_n353), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(G200), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n312), .A2(new_n403), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n215), .A2(G87), .ZN(new_n494));
  INV_X1    g0294(.A(new_n448), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT81), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(KEYINPUT19), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(KEYINPUT81), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n494), .B1(new_n500), .B2(new_n218), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n359), .A2(new_n218), .A3(G68), .ZN(new_n502));
  XNOR2_X1  g0302(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n218), .A2(G33), .A3(G97), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT82), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(G20), .B1(new_n270), .B2(new_n271), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n508), .A2(G68), .B1(new_n503), .B2(new_n504), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n498), .A2(KEYINPUT81), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n496), .A2(KEYINPUT19), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n448), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n512), .A2(G20), .B1(G87), .B2(new_n215), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT82), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n509), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n507), .A2(new_n289), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n217), .A2(G33), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n312), .A2(new_n313), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G87), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n491), .A2(new_n493), .A3(new_n516), .A4(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT83), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n490), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n509), .A2(new_n513), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n313), .B1(new_n523), .B2(KEYINPUT82), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n492), .B1(new_n524), .B2(new_n515), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n525), .A2(KEYINPUT83), .A3(new_n491), .A4(new_n519), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n518), .A2(new_n403), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n525), .A2(new_n527), .B1(new_n386), .B2(new_n489), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n480), .A2(new_n333), .A3(new_n487), .A4(new_n488), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT80), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n529), .B(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n522), .A2(new_n526), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(G244), .B(new_n269), .C1(new_n275), .C2(new_n276), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(G33), .B2(G283), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n359), .A2(KEYINPUT4), .A3(G244), .A4(new_n269), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT78), .B1(new_n272), .B2(G250), .ZN(new_n537));
  OAI211_X1 g0337(.A(G250), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT78), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n535), .B(new_n536), .C1(new_n537), .C2(new_n540), .ZN(new_n541));
  XNOR2_X1  g0341(.A(KEYINPUT5), .B(G41), .ZN(new_n542));
  INV_X1    g0342(.A(new_n226), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n542), .A2(new_n482), .B1(new_n543), .B2(new_n261), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n541), .A2(new_n264), .B1(G257), .B2(new_n544), .ZN(new_n545));
  OR2_X1    g0345(.A1(KEYINPUT5), .A2(G41), .ZN(new_n546));
  NAND2_X1  g0346(.A1(KEYINPUT5), .A2(G41), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n481), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(G274), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n543), .B2(new_n261), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n545), .A2(G190), .A3(new_n551), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n413), .A2(KEYINPUT6), .A3(G97), .ZN(new_n553));
  XNOR2_X1  g0353(.A(G97), .B(G107), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT6), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI22_X1  g0356(.A1(new_n556), .A2(new_n218), .B1(new_n210), .B2(new_n426), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n413), .B1(new_n360), .B2(new_n361), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n289), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n318), .A2(new_n232), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n312), .A2(new_n313), .A3(G97), .A4(new_n517), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g0364(.A(new_n538), .B(KEYINPUT78), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n533), .A2(new_n534), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G283), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n536), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n264), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n544), .A2(G257), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n551), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n564), .B1(new_n571), .B2(G200), .ZN(new_n572));
  OAI21_X1  g0372(.A(G107), .B1(new_n368), .B2(new_n369), .ZN(new_n573));
  AND2_X1   g0373(.A1(G97), .A2(G107), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n555), .B1(new_n574), .B2(new_n214), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n413), .A2(KEYINPUT6), .A3(G97), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(G20), .B1(G77), .B2(new_n296), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n562), .B1(new_n579), .B2(new_n289), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n571), .B2(new_n386), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n545), .A2(new_n333), .A3(new_n551), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n552), .A2(new_n572), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(G264), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n584));
  OAI211_X1 g0384(.A(G257), .B(new_n269), .C1(new_n275), .C2(new_n276), .ZN(new_n585));
  INV_X1    g0385(.A(G303), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n584), .B(new_n585), .C1(new_n586), .C2(new_n359), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n264), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n544), .A2(G270), .B1(new_n550), .B2(new_n548), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n312), .A2(new_n313), .A3(G116), .A4(new_n517), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n567), .B(new_n218), .C1(G33), .C2(new_n232), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n478), .A2(G20), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n289), .A3(new_n593), .ZN(new_n594));
  XOR2_X1   g0394(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n309), .A2(new_n478), .A3(new_n311), .ZN(new_n597));
  NOR2_X1   g0397(.A1(KEYINPUT84), .A2(KEYINPUT20), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n592), .A2(new_n289), .A3(new_n593), .A4(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n591), .A2(new_n596), .A3(new_n597), .A4(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n590), .A2(new_n600), .A3(KEYINPUT21), .A4(G169), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n600), .A2(G179), .A3(new_n588), .A4(new_n589), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n386), .B1(new_n588), .B2(new_n589), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT21), .B1(new_n604), .B2(new_n600), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(G257), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n607));
  OAI211_X1 g0407(.A(G250), .B(new_n269), .C1(new_n275), .C2(new_n276), .ZN(new_n608));
  INV_X1    g0408(.A(G294), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n607), .B(new_n608), .C1(new_n404), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n264), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n544), .A2(G264), .B1(new_n550), .B2(new_n548), .ZN(new_n612));
  AOI21_X1  g0412(.A(G169), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n333), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT24), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n218), .B(G87), .C1(new_n275), .C2(new_n276), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT22), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT22), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n359), .A2(new_n619), .A3(new_n218), .A4(G87), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n413), .A2(KEYINPUT23), .A3(G20), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT23), .B1(new_n413), .B2(G20), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n622), .A2(new_n623), .B1(new_n478), .B2(new_n291), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n616), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n621), .A2(new_n616), .A3(new_n625), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n313), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n309), .A2(new_n413), .A3(new_n311), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT25), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n518), .A2(G107), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n615), .B1(new_n629), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n600), .B1(new_n590), .B2(G200), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n353), .B2(new_n590), .ZN(new_n637));
  AOI211_X1 g0437(.A(KEYINPUT24), .B(new_n624), .C1(new_n618), .C2(new_n620), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n289), .B1(new_n638), .B2(new_n626), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n632), .A2(new_n633), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n611), .A2(new_n612), .A3(G190), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n611), .A2(new_n612), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G200), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n639), .A2(new_n640), .A3(new_n641), .A4(new_n643), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n606), .A2(new_n635), .A3(new_n637), .A4(new_n644), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n475), .A2(new_n532), .A3(new_n583), .A4(new_n645), .ZN(G372));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n571), .A2(new_n386), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n582), .A3(new_n564), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n647), .B1(new_n532), .B2(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n639), .A2(new_n640), .A3(new_n641), .A4(new_n643), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n606), .B2(new_n635), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n480), .A2(G190), .A3(new_n487), .A4(new_n488), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n525), .A2(new_n491), .A3(new_n519), .A4(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n516), .A2(new_n527), .A3(new_n493), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n489), .A2(new_n386), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(new_n529), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n653), .A2(new_n583), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n647), .A3(new_n650), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n475), .B1(new_n651), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n335), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n389), .A2(new_n396), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n468), .A2(new_n420), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n473), .A2(new_n381), .A3(new_n390), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n664), .B1(new_n668), .B2(new_n331), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n663), .A2(new_n669), .ZN(G369));
  NAND3_X1  g0470(.A1(new_n217), .A2(new_n218), .A3(G13), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G343), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n600), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n606), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n637), .ZN(new_n679));
  XNOR2_X1  g0479(.A(KEYINPUT85), .B(G330), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n676), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n683), .B1(new_n639), .B2(new_n640), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n635), .B1(new_n652), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n635), .B2(new_n676), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n606), .A2(new_n676), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n635), .A2(new_n676), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n688), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n221), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n215), .A2(G87), .A3(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n699), .A2(KEYINPUT86), .B1(new_n224), .B2(new_n697), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(KEYINPUT86), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g0501(.A(new_n701), .B(KEYINPUT28), .Z(new_n702));
  NAND4_X1  g0502(.A1(new_n655), .A2(new_n658), .A3(new_n582), .A4(new_n581), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT88), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n658), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n656), .A2(KEYINPUT88), .A3(new_n657), .A4(new_n529), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n703), .A2(KEYINPUT26), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n520), .A2(new_n521), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(new_n526), .A3(new_n654), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n528), .A2(new_n531), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(new_n647), .A3(new_n650), .A4(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(new_n660), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(KEYINPUT29), .A3(new_n683), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n660), .A2(new_n658), .A3(new_n661), .ZN(new_n714));
  INV_X1    g0514(.A(new_n651), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n676), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n713), .B1(new_n716), .B2(KEYINPUT29), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n588), .A2(new_n589), .A3(G179), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n718), .A2(new_n489), .A3(new_n642), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n545), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n571), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n489), .A2(new_n590), .A3(new_n642), .A4(new_n333), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT87), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n722), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT30), .B1(new_n719), .B2(new_n545), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n723), .A2(new_n724), .ZN(new_n729));
  OAI21_X1  g0529(.A(KEYINPUT87), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n719), .A2(KEYINPUT30), .A3(new_n545), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n683), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n722), .A2(new_n725), .A3(new_n731), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n676), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n732), .A2(new_n734), .B1(new_n736), .B2(new_n733), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n645), .A2(new_n532), .A3(new_n583), .A4(new_n683), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n680), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n717), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n702), .B1(new_n741), .B2(G1), .ZN(G364));
  NAND2_X1  g0542(.A1(new_n679), .A2(new_n680), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n218), .A2(G13), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n217), .B1(new_n744), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n682), .B(new_n743), .C1(new_n696), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n679), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n696), .A2(new_n746), .ZN(new_n752));
  XOR2_X1   g0552(.A(new_n752), .B(KEYINPUT89), .Z(new_n753));
  INV_X1    g0553(.A(KEYINPUT90), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n221), .B(new_n359), .C1(new_n754), .C2(G355), .ZN(new_n755));
  AOI21_X1  g0555(.A(KEYINPUT90), .B1(new_n215), .B2(G87), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n756), .B1(G116), .B2(new_n221), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n359), .B(new_n695), .C1(new_n259), .C2(new_n225), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n255), .A2(G45), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n226), .B1(G20), .B2(new_n386), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n750), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n753), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n353), .A2(G179), .A3(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n218), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(G20), .A2(G179), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n768), .A2(G190), .A3(G200), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n767), .A2(G294), .B1(new_n769), .B2(G311), .ZN(new_n770));
  INV_X1    g0570(.A(G326), .ZN(new_n771));
  INV_X1    g0571(.A(new_n768), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n772), .A2(G190), .A3(G200), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n770), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT93), .Z(new_n775));
  NAND3_X1  g0575(.A1(new_n772), .A2(new_n353), .A3(G200), .ZN(new_n776));
  OR2_X1    g0576(.A1(KEYINPUT33), .A2(G317), .ZN(new_n777));
  NAND2_X1  g0577(.A1(KEYINPUT33), .A2(G317), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n768), .A2(new_n353), .A3(G200), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n359), .B(new_n779), .C1(G322), .C2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(KEYINPUT91), .B1(new_n353), .B2(G20), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n353), .A2(KEYINPUT91), .A3(G20), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G329), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n785), .A2(new_n285), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G283), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n333), .A2(G20), .A3(G190), .A4(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n791), .A2(KEYINPUT92), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(KEYINPUT92), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G303), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n781), .A2(new_n787), .A3(new_n789), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n773), .A2(new_n202), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n766), .A2(new_n232), .ZN(new_n798));
  INV_X1    g0598(.A(new_n776), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n797), .B(new_n798), .C1(G68), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n780), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n359), .B1(new_n801), .B2(new_n230), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G77), .B2(new_n769), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n788), .A2(G107), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n794), .A2(G87), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n800), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n786), .A2(G159), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT32), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n775), .A2(new_n796), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n764), .B1(new_n809), .B2(new_n761), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n751), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n747), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(G396));
  OR2_X1    g0613(.A1(new_n420), .A2(new_n676), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n421), .A2(new_n422), .B1(new_n409), .B2(new_n683), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n420), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n716), .B(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n752), .B1(new_n818), .B2(new_n740), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n740), .B2(new_n818), .ZN(new_n820));
  INV_X1    g0620(.A(new_n753), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n761), .A2(new_n748), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(new_n210), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n761), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G143), .A2(new_n780), .B1(new_n769), .B2(G159), .ZN(new_n825));
  INV_X1    g0625(.A(G137), .ZN(new_n826));
  INV_X1    g0626(.A(G150), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n826), .B2(new_n773), .C1(new_n827), .C2(new_n776), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT34), .Z(new_n829));
  INV_X1    g0629(.A(KEYINPUT94), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n794), .A2(G50), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n788), .A2(G68), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n786), .A2(G132), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n280), .B1(new_n767), .B2(G58), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n831), .A2(new_n832), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n829), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n835), .A2(new_n830), .ZN(new_n837));
  INV_X1    g0637(.A(new_n769), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n280), .B1(new_n838), .B2(new_n478), .C1(new_n609), .C2(new_n801), .ZN(new_n839));
  INV_X1    g0639(.A(new_n773), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n798), .B1(G303), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(G283), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n842), .B2(new_n776), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n839), .B(new_n843), .C1(G107), .C2(new_n794), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G87), .A2(new_n788), .B1(new_n786), .B2(G311), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n836), .A2(new_n837), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n823), .B1(new_n824), .B2(new_n846), .C1(new_n817), .C2(new_n749), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n820), .A2(new_n847), .ZN(G384));
  NAND2_X1  g0648(.A1(new_n814), .A2(new_n816), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n443), .A2(new_n676), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n468), .A2(new_n473), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(G169), .B1(new_n456), .B2(new_n460), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT14), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(new_n464), .A3(new_n461), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n443), .B(new_n676), .C1(new_n854), .C2(new_n472), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n849), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n736), .A2(new_n733), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n738), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT99), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n674), .B1(new_n378), .B2(new_n373), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n397), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n391), .A2(new_n394), .ZN(new_n863));
  INV_X1    g0663(.A(new_n674), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n367), .A2(new_n372), .A3(new_n289), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n864), .B1(new_n865), .B2(new_n382), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n355), .A2(new_n373), .A3(new_n378), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n863), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT37), .B1(new_n861), .B2(KEYINPUT96), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n868), .B(KEYINPUT37), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT38), .B1(new_n874), .B2(new_n862), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT40), .B1(new_n860), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n878), .A2(KEYINPUT99), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n856), .A2(new_n859), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n872), .A2(KEYINPUT97), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n397), .A2(new_n861), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n868), .B(new_n869), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n868), .A2(new_n869), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n868), .A2(new_n869), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT97), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT38), .A4(new_n862), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n881), .A2(new_n878), .A3(new_n885), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n880), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n877), .A2(new_n892), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n475), .A2(new_n859), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n680), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n893), .B2(new_n894), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT100), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n898), .B2(new_n897), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n881), .A2(KEYINPUT39), .A3(new_n885), .A4(new_n890), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n854), .A2(new_n443), .A3(new_n683), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n873), .B2(new_n875), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n901), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n851), .A2(new_n855), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n817), .B(new_n683), .C1(new_n662), .C2(new_n651), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(new_n908), .B2(new_n814), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n881), .A2(new_n885), .A3(new_n890), .ZN(new_n910));
  INV_X1    g0710(.A(new_n665), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n909), .A2(new_n910), .B1(new_n911), .B2(new_n674), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT98), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n906), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n908), .A2(new_n814), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n851), .A2(new_n855), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n910), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n911), .A2(new_n674), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n917), .A2(new_n913), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n475), .B(new_n713), .C1(new_n716), .C2(KEYINPUT29), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n669), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(new_n922), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n900), .A2(new_n923), .B1(new_n217), .B2(new_n744), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n923), .B2(new_n900), .ZN(new_n925));
  OR3_X1    g0725(.A1(new_n224), .A2(new_n210), .A3(new_n363), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n211), .A2(G68), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n217), .B(G13), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n577), .A2(KEYINPUT35), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n577), .A2(KEYINPUT35), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n929), .A2(new_n930), .A3(G116), .A4(new_n227), .ZN(new_n931));
  XOR2_X1   g0731(.A(KEYINPUT95), .B(KEYINPUT36), .Z(new_n932));
  XNOR2_X1  g0732(.A(new_n931), .B(new_n932), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n925), .A2(new_n928), .A3(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT101), .Z(G367));
  NOR2_X1   g0735(.A1(new_n695), .A2(new_n359), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n247), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n763), .B1(new_n695), .B2(new_n403), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n821), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT104), .Z(new_n940));
  INV_X1    g0740(.A(new_n750), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n525), .A2(new_n519), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n676), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n659), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n658), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT46), .ZN(new_n947));
  INV_X1    g0747(.A(new_n794), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n947), .B1(new_n948), .B2(new_n478), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n788), .A2(G97), .ZN(new_n950));
  XOR2_X1   g0750(.A(KEYINPUT105), .B(G317), .Z(new_n951));
  NAND2_X1  g0751(.A1(new_n786), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n794), .A2(KEYINPUT46), .A3(G116), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n949), .A2(new_n950), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n280), .B1(new_n801), .B2(new_n586), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G283), .B2(new_n769), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n767), .A2(G107), .B1(new_n840), .B2(G311), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n956), .B(new_n957), .C1(new_n609), .C2(new_n776), .ZN(new_n958));
  INV_X1    g0758(.A(G159), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n776), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n766), .A2(new_n357), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(G143), .C2(new_n840), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n359), .B1(new_n801), .B2(new_n827), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n206), .B2(new_n769), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n962), .B(new_n964), .C1(new_n230), .C2(new_n948), .ZN(new_n965));
  INV_X1    g0765(.A(new_n788), .ZN(new_n966));
  INV_X1    g0766(.A(new_n786), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n210), .A2(new_n966), .B1(new_n967), .B2(new_n826), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n954), .A2(new_n958), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT47), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n761), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n940), .B1(new_n941), .B2(new_n946), .C1(new_n971), .C2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n583), .B1(new_n580), .B2(new_n683), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n649), .B2(new_n683), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n691), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT42), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n975), .A2(new_n635), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n676), .B1(new_n979), .B2(new_n649), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT102), .ZN(new_n982));
  AND3_X1   g0782(.A1(new_n981), .A2(new_n982), .A3(new_n946), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n946), .B1(new_n981), .B2(new_n982), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(KEYINPUT43), .B1(new_n983), .B2(new_n984), .ZN(new_n988));
  AND4_X1   g0788(.A1(new_n687), .A2(new_n987), .A3(new_n976), .A4(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n987), .A2(new_n988), .B1(new_n687), .B2(new_n976), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n693), .A2(new_n976), .ZN(new_n992));
  XOR2_X1   g0792(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n693), .A2(new_n976), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT45), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n994), .A2(new_n996), .A3(new_n687), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n686), .B(new_n690), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(new_n681), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n741), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n687), .B1(new_n994), .B2(new_n996), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n997), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n741), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n696), .B(KEYINPUT41), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n746), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n974), .B1(new_n991), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT106), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(G387));
  NAND2_X1  g0809(.A1(new_n999), .A2(new_n746), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n951), .A2(new_n780), .B1(new_n769), .B2(G303), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n840), .A2(G322), .ZN(new_n1012));
  INV_X1    g0812(.A(G311), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1011), .B(new_n1012), .C1(new_n1013), .C2(new_n776), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT48), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n794), .A2(G294), .B1(G283), .B2(new_n767), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT49), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n280), .B1(new_n967), .B2(new_n771), .C1(new_n478), .C2(new_n966), .ZN(new_n1023));
  OR3_X1    g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n773), .A2(new_n959), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT108), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G77), .B2(new_n794), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n359), .B1(new_n838), .B2(new_n357), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n766), .A2(new_n402), .B1(new_n776), .B2(new_n300), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G50), .C2(new_n780), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n786), .A2(G150), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n1030), .A3(new_n950), .A4(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n824), .B1(new_n1024), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n400), .A2(new_n202), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT50), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n698), .B(new_n259), .C1(new_n357), .C2(new_n210), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n936), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1037), .A2(KEYINPUT107), .B1(G45), .B2(new_n244), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(KEYINPUT107), .B2(new_n1037), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n221), .A2(new_n359), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1039), .B1(G107), .B2(new_n221), .C1(new_n698), .C2(new_n1040), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n821), .B(new_n1033), .C1(new_n762), .C2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1042), .A2(KEYINPUT109), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(KEYINPUT109), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n686), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1044), .B1(new_n1045), .B2(new_n941), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1000), .A2(new_n696), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n741), .A2(new_n999), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1010), .B1(new_n1043), .B2(new_n1046), .C1(new_n1047), .C2(new_n1048), .ZN(G393));
  NAND2_X1  g0849(.A1(new_n1002), .A2(KEYINPUT110), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(new_n997), .Z(new_n1051));
  OAI211_X1 g0851(.A(new_n696), .B(new_n1003), .C1(new_n1051), .C2(new_n1001), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n976), .A2(new_n941), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n762), .B1(new_n232), .B2(new_n221), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n252), .B2(new_n936), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n821), .A2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT111), .Z(new_n1057));
  NOR2_X1   g0857(.A1(new_n766), .A2(new_n478), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n280), .B1(new_n776), .B2(new_n586), .C1(new_n838), .C2(new_n609), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(G283), .C2(new_n794), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n786), .A2(G322), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1060), .A2(new_n804), .A3(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n840), .A2(G317), .B1(G311), .B2(new_n780), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT52), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1065), .A2(KEYINPUT112), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(KEYINPUT112), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n766), .A2(new_n210), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n359), .B1(new_n838), .B2(new_n300), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n206), .C2(new_n799), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n801), .A2(new_n959), .B1(new_n773), .B2(new_n827), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT51), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G87), .A2(new_n788), .B1(new_n786), .B2(G143), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n794), .A2(G68), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1066), .A2(new_n1067), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1057), .B1(new_n1076), .B2(new_n761), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1051), .A2(new_n746), .B1(new_n1053), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1052), .A2(new_n1078), .ZN(G390));
  NAND3_X1  g0879(.A1(new_n712), .A2(new_n683), .A3(new_n816), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n814), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT113), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1080), .A2(KEYINPUT113), .A3(new_n814), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n916), .A3(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n876), .A2(new_n903), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n901), .A2(new_n905), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n909), .B2(new_n903), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n739), .A2(new_n817), .A3(new_n916), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n915), .A2(new_n916), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n902), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1088), .A2(new_n1093), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n856), .A2(G330), .A3(new_n859), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1091), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n475), .A2(G330), .A3(new_n859), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n921), .A2(new_n669), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n916), .B1(new_n739), .B2(new_n817), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n915), .B1(new_n1100), .B2(new_n1095), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n859), .A2(G330), .A3(new_n817), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n907), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1084), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT113), .B1(new_n1080), .B2(new_n814), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1090), .B(new_n1103), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1099), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1097), .A2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1091), .B(new_n1107), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n696), .A3(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1091), .B(new_n746), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT115), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n822), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n753), .B1(new_n400), .B2(new_n1114), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n280), .B1(new_n838), .B2(new_n232), .C1(new_n478), .C2(new_n801), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n794), .B2(G87), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n773), .A2(new_n842), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1118), .B(new_n1068), .C1(G107), .C2(new_n799), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n786), .A2(G294), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1117), .A2(new_n832), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n794), .A2(G150), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT53), .Z(new_n1123));
  OAI22_X1  g0923(.A1(new_n766), .A2(new_n959), .B1(new_n776), .B2(new_n826), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT54), .B(G143), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1126), .A2(new_n769), .B1(new_n780), .B2(G132), .ZN(new_n1127));
  INV_X1    g0927(.A(G128), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1127), .B1(new_n1128), .B2(new_n773), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1124), .B(new_n1129), .C1(G125), .C2(new_n786), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1123), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n280), .B1(new_n788), .B2(new_n206), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT114), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1121), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1115), .B1(new_n1134), .B2(new_n761), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1088), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1135), .B1(new_n1136), .B2(new_n749), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1112), .A2(new_n1113), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1113), .B1(new_n1112), .B2(new_n1137), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1111), .B1(new_n1138), .B2(new_n1139), .ZN(G378));
  NAND2_X1  g0940(.A1(new_n893), .A2(G330), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n320), .A2(new_n864), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n331), .A2(new_n335), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n331), .B2(new_n335), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1144), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n336), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n331), .A2(new_n335), .A3(new_n1144), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n1150), .A3(new_n1142), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1147), .A2(new_n1151), .A3(KEYINPUT118), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1141), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1152), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n893), .A2(G330), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n920), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n917), .A2(new_n918), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT98), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n912), .A2(new_n913), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1159), .A3(new_n906), .ZN(new_n1160));
  INV_X1    g0960(.A(G330), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1161), .B(new_n1152), .C1(new_n877), .C2(new_n892), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1154), .B1(new_n893), .B2(G330), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1160), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1099), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1156), .A2(new_n1164), .B1(new_n1110), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n696), .B1(new_n1166), .B2(KEYINPUT57), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1156), .A2(new_n1164), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1110), .A2(new_n1165), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1168), .A2(KEYINPUT57), .A3(new_n1169), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1147), .A2(new_n1151), .A3(new_n748), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n752), .B1(new_n206), .B2(new_n1114), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(G33), .A2(G41), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT116), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n202), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n258), .B2(new_n280), .ZN(new_n1177));
  AOI211_X1 g0977(.A(G41), .B(new_n359), .C1(G107), .C2(new_n780), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n402), .B2(new_n838), .C1(new_n948), .C2(new_n210), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n230), .A2(new_n966), .B1(new_n967), .B2(new_n842), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n961), .B1(G97), .B2(new_n799), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n478), .B2(new_n773), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1177), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n801), .A2(new_n1128), .B1(new_n838), .B2(new_n826), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G132), .B2(new_n799), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n767), .A2(G150), .B1(new_n840), .B2(G125), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(new_n948), .C2(new_n1125), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1175), .B1(new_n786), .B2(G124), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(new_n959), .C2(new_n966), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1185), .B1(new_n1190), .B2(new_n1193), .C1(new_n1184), .C2(new_n1183), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1173), .B1(new_n1194), .B2(new_n761), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1168), .A2(new_n746), .B1(new_n1172), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1171), .A2(new_n1196), .ZN(G375));
  NAND3_X1  g0997(.A1(new_n1101), .A2(new_n1106), .A3(new_n1099), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1108), .A2(new_n1005), .A3(new_n1198), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT119), .Z(new_n1200));
  NAND2_X1  g1000(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n745), .B(KEYINPUT120), .Z(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n753), .B1(G68), .B2(new_n1114), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n948), .A2(new_n232), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n280), .B1(new_n838), .B2(new_n413), .C1(new_n842), .C2(new_n801), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n767), .A2(new_n403), .B1(new_n799), .B2(G116), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(new_n609), .C2(new_n773), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n210), .A2(new_n966), .B1(new_n967), .B2(new_n586), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n794), .A2(G159), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n799), .A2(new_n1126), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n767), .A2(G50), .B1(new_n840), .B2(G132), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n359), .B1(new_n838), .B2(new_n827), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G137), .B2(new_n780), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1216), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n230), .A2(new_n966), .B1(new_n967), .B2(new_n1128), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n1210), .A2(new_n1211), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1205), .B1(new_n1219), .B2(new_n761), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n916), .B2(new_n749), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1204), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1200), .A2(new_n1223), .ZN(G381));
  NOR4_X1   g1024(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1008), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(G375), .ZN(new_n1227));
  INV_X1    g1027(.A(G381), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1111), .A2(new_n1112), .A3(new_n1137), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(G407));
  INV_X1    g1030(.A(new_n1229), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n675), .A2(G213), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT121), .Z(new_n1233));
  OR3_X1    g1033(.A1(G375), .A2(new_n1231), .A3(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(G407), .A2(G213), .A3(new_n1234), .ZN(G409));
  XNOR2_X1  g1035(.A(G393), .B(new_n812), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(KEYINPUT106), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(G390), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1236), .B1(new_n1052), .B2(new_n1078), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n974), .B1(new_n1006), .B2(new_n991), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1007), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1240), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT60), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1198), .B1(new_n1107), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT123), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n696), .B1(new_n1198), .B2(new_n1245), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1251), .A2(G384), .A3(new_n1223), .ZN(new_n1252));
  AOI21_X1  g1052(.A(G384), .B1(new_n1251), .B2(new_n1223), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(G2897), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1233), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n1252), .A2(new_n1253), .B1(new_n1255), .B2(new_n1233), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT125), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1259), .B(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1156), .A2(new_n1164), .A3(KEYINPUT122), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1203), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT122), .B1(new_n1156), .B2(new_n1164), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1168), .A2(new_n1005), .A3(new_n1169), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1172), .A2(new_n1195), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1229), .B1(new_n1265), .B2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G378), .B(new_n1196), .C1(new_n1167), .C2(new_n1170), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1233), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1244), .B1(new_n1261), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1233), .A3(new_n1254), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT63), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT124), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1271), .A2(new_n1254), .A3(KEYINPUT124), .A4(new_n1233), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1273), .B(new_n1276), .C1(KEYINPUT63), .C2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1272), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1243), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT126), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1278), .A2(new_n1285), .A3(new_n1286), .A4(new_n1279), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1275), .A2(KEYINPUT62), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT126), .B1(new_n1280), .B2(KEYINPUT62), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1284), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1240), .A2(new_n1242), .A3(KEYINPUT127), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT127), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1293));
  OR2_X1    g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1281), .B1(new_n1291), .B2(new_n1294), .ZN(G405));
  OAI21_X1  g1095(.A(new_n1270), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1254), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(new_n1296), .B(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1294), .B(new_n1298), .ZN(G402));
endmodule


