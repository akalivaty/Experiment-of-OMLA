//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n571, new_n572, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n634, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n468), .A2(KEYINPUT67), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(new_n467), .A3(G2104), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n475), .A2(new_n464), .A3(new_n466), .A4(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n474), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n472), .A2(new_n480), .ZN(G160));
  NAND4_X1  g056(.A1(new_n475), .A2(G2105), .A3(new_n466), .A4(new_n477), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n464), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI22_X1  g060(.A1(new_n482), .A2(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n478), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(G136), .B2(new_n487), .ZN(G162));
  INV_X1    g063(.A(new_n482), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n464), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OR3_X1    g068(.A1(new_n491), .A2(new_n492), .A3(new_n490), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n489), .A2(G126), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n464), .A2(G138), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n475), .A2(new_n466), .A3(new_n477), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n466), .A2(new_n468), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT69), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n469), .A2(new_n503), .A3(new_n499), .A4(new_n496), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n498), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  AND3_X1   g081(.A1(new_n495), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n506), .B1(new_n495), .B2(new_n505), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(G164));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G62), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n515), .A2(G651), .B1(G50), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n512), .A2(new_n511), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT71), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n517), .A2(new_n518), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT5), .B(G543), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT72), .B(G88), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n524), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n520), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  INV_X1    g107(.A(new_n512), .ZN(new_n533));
  NAND2_X1  g108(.A1(KEYINPUT5), .A2(G543), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n533), .A2(KEYINPUT73), .A3(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n536), .B1(new_n511), .B2(new_n512), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n535), .A2(new_n537), .A3(G63), .A4(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n541));
  AOI22_X1  g116(.A1(G51), .A2(new_n519), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n524), .A2(new_n528), .ZN(new_n543));
  INV_X1    g118(.A(G89), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n538), .B(new_n542), .C1(new_n543), .C2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND3_X1  g121(.A1(new_n535), .A2(new_n537), .A3(G64), .ZN(new_n547));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n519), .A2(G52), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n524), .A2(G90), .A3(new_n528), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND3_X1  g129(.A1(new_n524), .A2(G81), .A3(new_n528), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n519), .A2(G43), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G651), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n535), .A2(new_n537), .A3(G56), .ZN(new_n559));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT74), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n560), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n564), .A2(new_n565), .A3(new_n556), .A4(new_n555), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  AOI22_X1  g148(.A1(new_n526), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n558), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n524), .A2(G91), .A3(new_n528), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n524), .A2(KEYINPUT78), .A3(G91), .A4(new_n528), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT9), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(KEYINPUT75), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(KEYINPUT76), .B2(new_n581), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n583), .A2(new_n519), .A3(G53), .ZN(new_n584));
  OAI211_X1 g159(.A(G53), .B(G543), .C1(new_n521), .C2(new_n522), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n582), .B1(new_n585), .B2(KEYINPUT76), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT77), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n587), .B1(new_n584), .B2(new_n586), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n580), .A2(new_n590), .ZN(G299));
  INV_X1    g166(.A(new_n543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G87), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n535), .A2(new_n537), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n594), .B2(G74), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n519), .A2(G49), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(G288));
  NAND3_X1  g172(.A1(new_n524), .A2(G86), .A3(new_n528), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G73), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G61), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n513), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G48), .B2(new_n519), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(G305));
  NAND3_X1  g180(.A1(new_n535), .A2(new_n537), .A3(G60), .ZN(new_n606));
  NAND2_X1  g181(.A1(G72), .A2(G543), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G651), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n519), .A2(G47), .ZN(new_n611));
  INV_X1    g186(.A(G85), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n543), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT80), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n592), .A2(G85), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n615), .A2(new_n616), .A3(new_n609), .A4(new_n611), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n614), .A2(new_n617), .ZN(G290));
  NAND2_X1  g193(.A1(G301), .A2(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  INV_X1    g195(.A(G66), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n513), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G651), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n519), .A2(G54), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n524), .A2(G92), .A3(new_n528), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g203(.A1(new_n524), .A2(KEYINPUT10), .A3(G92), .A4(new_n528), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n619), .B1(G868), .B2(new_n630), .ZN(G284));
  XNOR2_X1  g206(.A(G284), .B(KEYINPUT81), .ZN(G321));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(G299), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(G168), .ZN(G297));
  OAI21_X1  g210(.A(new_n634), .B1(new_n633), .B2(G168), .ZN(G280));
  INV_X1    g211(.A(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n630), .B1(new_n637), .B2(G860), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT82), .Z(G148));
  NAND2_X1  g214(.A1(new_n630), .A2(new_n637), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G868), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n568), .B2(G868), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g219(.A1(new_n469), .A2(new_n473), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT12), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT13), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2100), .ZN(new_n648));
  INV_X1    g223(.A(G2096), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n651));
  INV_X1    g226(.A(G111), .ZN(new_n652));
  AOI22_X1  g227(.A1(new_n650), .A2(new_n651), .B1(new_n652), .B2(G2105), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n651), .B2(new_n650), .ZN(new_n654));
  INV_X1    g229(.A(G135), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n478), .B2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(G123), .ZN(new_n657));
  OR3_X1    g232(.A1(new_n482), .A2(KEYINPUT84), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(KEYINPUT84), .B1(new_n482), .B2(new_n657), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n648), .B1(new_n649), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n649), .B2(new_n660), .ZN(G156));
  XNOR2_X1  g237(.A(G2427), .B(G2438), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2430), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT15), .B(G2435), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(KEYINPUT14), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1341), .B(G1348), .Z(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2451), .B(G2454), .Z(new_n673));
  XNOR2_X1  g248(.A(G2443), .B(G2446), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n672), .A2(new_n675), .ZN(new_n677));
  AND3_X1   g252(.A1(new_n676), .A2(G14), .A3(new_n677), .ZN(G401));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT87), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT17), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2084), .B(G2090), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n680), .B2(new_n682), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n681), .B2(new_n682), .ZN(new_n686));
  INV_X1    g261(.A(new_n682), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n687), .A2(new_n683), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n680), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT18), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n684), .A2(new_n686), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G2100), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT88), .B(G2096), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G227));
  XOR2_X1   g269(.A(G1961), .B(G1966), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT89), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1956), .B(G2474), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1971), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT19), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT20), .Z(new_n703));
  OR2_X1    g278(.A1(new_n696), .A2(new_n698), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n704), .A2(new_n701), .A3(new_n699), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n703), .B(new_n705), .C1(new_n701), .C2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT90), .ZN(new_n707));
  XOR2_X1   g282(.A(G1981), .B(G1986), .Z(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n707), .B(new_n712), .ZN(G229));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G23), .ZN(new_n715));
  INV_X1    g290(.A(G288), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n714), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT92), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT33), .B(G1976), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n714), .A2(G22), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G166), .B2(new_n714), .ZN(new_n722));
  INV_X1    g297(.A(G1971), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n714), .A2(G6), .ZN(new_n725));
  INV_X1    g300(.A(G305), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n714), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT32), .B(G1981), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n728), .B2(new_n727), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n720), .A2(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(KEYINPUT34), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(KEYINPUT34), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G25), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n487), .A2(G131), .ZN(new_n736));
  INV_X1    g311(.A(G119), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n464), .A2(G107), .ZN(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n739));
  OAI22_X1  g314(.A1(new_n482), .A2(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(new_n734), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT35), .B(G1991), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT91), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n742), .B(new_n744), .Z(new_n745));
  AND2_X1   g320(.A1(new_n714), .A2(G24), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G290), .B2(G16), .ZN(new_n747));
  INV_X1    g322(.A(G1986), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n748), .B2(new_n747), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n732), .A2(new_n733), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT93), .B(KEYINPUT36), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n734), .A2(G32), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n489), .A2(G129), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT99), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT100), .B(KEYINPUT26), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G105), .B2(new_n473), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n487), .A2(G141), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT98), .Z(new_n764));
  AND2_X1   g339(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n754), .B1(new_n765), .B2(new_n734), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT27), .ZN(new_n767));
  INV_X1    g342(.A(G1996), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(G168), .A2(G16), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G16), .B2(G21), .ZN(new_n771));
  INV_X1    g346(.A(G1966), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  AOI211_X1 g349(.A(new_n773), .B(new_n774), .C1(G29), .C2(new_n660), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT24), .ZN(new_n776));
  INV_X1    g351(.A(G34), .ZN(new_n777));
  AOI21_X1  g352(.A(G29), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n776), .B2(new_n777), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G160), .B2(new_n734), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G2084), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT31), .B(G11), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT30), .B(G28), .Z(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G29), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n734), .A2(G33), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT25), .Z(new_n787));
  INV_X1    g362(.A(G139), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  OAI221_X1 g364(.A(new_n787), .B1(new_n788), .B2(new_n478), .C1(new_n789), .C2(new_n464), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n785), .B1(new_n790), .B2(G29), .ZN(new_n791));
  INV_X1    g366(.A(G2072), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n784), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AND3_X1   g368(.A1(new_n775), .A2(new_n781), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n734), .A2(G27), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT101), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G164), .B2(new_n734), .ZN(new_n797));
  INV_X1    g372(.A(G2078), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n714), .A2(G5), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G171), .B2(new_n714), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G1961), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G2084), .B2(new_n780), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n801), .A2(G1961), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n791), .A2(new_n792), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT97), .Z(new_n807));
  NAND4_X1  g382(.A1(new_n794), .A2(new_n799), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n769), .A2(new_n808), .A3(KEYINPUT102), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT102), .B1(new_n769), .B2(new_n808), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n734), .A2(G26), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(G104), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n815));
  INV_X1    g390(.A(G140), .ZN(new_n816));
  INV_X1    g391(.A(G128), .ZN(new_n817));
  OAI221_X1 g392(.A(new_n815), .B1(new_n478), .B2(new_n816), .C1(new_n817), .C2(new_n482), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(new_n734), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT96), .B(G2067), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(G4), .A2(G16), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n630), .B2(G16), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT94), .B(G1348), .Z(new_n825));
  AOI21_X1  g400(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT103), .B(KEYINPUT23), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n714), .A2(G20), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G299), .B2(G16), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G1956), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n826), .B(new_n831), .C1(new_n824), .C2(new_n825), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n734), .A2(G35), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G162), .B2(new_n734), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT29), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G2090), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n714), .A2(G19), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n568), .B2(new_n714), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G1341), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n832), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n809), .A2(new_n810), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n753), .A2(new_n841), .ZN(G311));
  INV_X1    g417(.A(G311), .ZN(G150));
  NAND3_X1  g418(.A1(new_n524), .A2(G93), .A3(new_n528), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n519), .A2(G55), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n535), .A2(new_n537), .A3(G67), .ZN(new_n847));
  NAND2_X1  g422(.A1(G80), .A2(G543), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n558), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(G860), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n847), .A2(new_n848), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n845), .B(new_n844), .C1(new_n854), .C2(new_n558), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n567), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n564), .A2(new_n556), .A3(new_n555), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n630), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT104), .Z(new_n866));
  OAI21_X1  g441(.A(new_n851), .B1(new_n863), .B2(new_n864), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n853), .B1(new_n866), .B2(new_n867), .ZN(G145));
  NAND2_X1  g443(.A1(new_n495), .A2(new_n505), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n819), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n765), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n762), .A2(new_n764), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n870), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n790), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n790), .A2(new_n875), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n872), .A2(new_n874), .A3(new_n878), .A4(new_n876), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(G106), .A2(G2105), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n883), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n884));
  INV_X1    g459(.A(G142), .ZN(new_n885));
  INV_X1    g460(.A(G130), .ZN(new_n886));
  OAI221_X1 g461(.A(new_n884), .B1(new_n478), .B2(new_n885), .C1(new_n886), .C2(new_n482), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT106), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n646), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n741), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n882), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n880), .A2(new_n890), .A3(new_n881), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(G162), .B(G160), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n895), .B(new_n660), .Z(new_n896));
  AOI21_X1  g471(.A(G37), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n896), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n892), .A2(new_n898), .A3(new_n893), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n897), .A2(KEYINPUT107), .A3(new_n899), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n902), .A2(KEYINPUT40), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT40), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(G395));
  NAND2_X1  g481(.A1(new_n855), .A2(new_n633), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n860), .B(new_n640), .ZN(new_n908));
  INV_X1    g483(.A(new_n630), .ZN(new_n909));
  NAND2_X1  g484(.A1(G299), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n580), .A2(new_n630), .A3(new_n590), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT108), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n580), .A2(new_n630), .A3(new_n590), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n628), .A2(new_n629), .ZN(new_n916));
  INV_X1    g491(.A(new_n625), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n580), .A2(new_n590), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n915), .A2(new_n918), .A3(KEYINPUT41), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n920), .B1(new_n910), .B2(new_n911), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n914), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n910), .A2(new_n920), .A3(new_n911), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT108), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n913), .B1(new_n925), .B2(new_n908), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT42), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n726), .A2(G288), .ZN(new_n928));
  NAND2_X1  g503(.A1(G305), .A2(new_n716), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(G303), .B(KEYINPUT109), .ZN(new_n931));
  NAND2_X1  g506(.A1(G290), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(G290), .A2(new_n931), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n934), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n936), .A2(new_n929), .A3(new_n928), .A4(new_n932), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n927), .B(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n907), .B1(new_n940), .B2(new_n633), .ZN(G295));
  OAI21_X1  g516(.A(new_n907), .B1(new_n940), .B2(new_n633), .ZN(G331));
  INV_X1    g517(.A(G37), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n552), .A2(new_n551), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n558), .B1(new_n547), .B2(new_n548), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n550), .A2(KEYINPUT110), .A3(new_n551), .A4(new_n552), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(G168), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n948), .A3(G286), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n856), .A2(new_n950), .A3(new_n859), .A4(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n947), .A2(new_n948), .A3(G286), .ZN(new_n953));
  AOI21_X1  g528(.A(G286), .B1(new_n947), .B2(new_n948), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n850), .B1(new_n562), .B2(new_n566), .ZN(new_n955));
  OAI22_X1  g530(.A1(new_n953), .A2(new_n954), .B1(new_n955), .B2(new_n858), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n912), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT41), .B1(new_n915), .B2(new_n918), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n923), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n952), .A2(new_n956), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n943), .B1(new_n961), .B2(new_n938), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT108), .B1(new_n958), .B2(new_n923), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n915), .A2(new_n918), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n914), .B1(new_n964), .B2(new_n920), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n960), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n957), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n938), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n966), .A2(KEYINPUT111), .A3(new_n938), .A4(new_n967), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n962), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n957), .B1(new_n925), .B2(new_n960), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n943), .B1(new_n975), .B2(new_n938), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n970), .B2(new_n971), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n974), .B1(new_n977), .B2(new_n973), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n962), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT111), .B1(new_n975), .B2(new_n938), .ZN(new_n982));
  INV_X1    g557(.A(new_n971), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n985), .A3(KEYINPUT43), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT112), .B1(new_n972), .B2(new_n973), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n979), .B1(new_n977), .B2(new_n973), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n989), .B1(new_n988), .B2(new_n990), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n980), .B1(new_n991), .B2(new_n992), .ZN(G397));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n869), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n996));
  XOR2_X1   g571(.A(KEYINPUT114), .B(G40), .Z(new_n997));
  NOR3_X1   g572(.A1(new_n472), .A2(new_n480), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n873), .A2(G1996), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  INV_X1    g579(.A(G2067), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n818), .B(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n873), .B2(G1996), .ZN(new_n1007));
  AOI211_X1 g582(.A(new_n1003), .B(new_n1004), .C1(new_n1000), .C2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n741), .B(new_n744), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n999), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(G290), .B(G1986), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1000), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(G288), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1384), .B1(new_n495), .B2(new_n505), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n998), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1017), .B(G8), .C1(G288), .C2(new_n1013), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(KEYINPUT52), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1981), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n604), .B2(new_n598), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(G305), .B2(G1981), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT116), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1017), .A2(G8), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1025), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1029), .B1(new_n1030), .B2(KEYINPUT49), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1021), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G303), .A2(G8), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT55), .ZN(new_n1034));
  INV_X1    g609(.A(new_n997), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G160), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n995), .B2(KEYINPUT50), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n994), .B1(new_n507), .B2(new_n508), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(new_n1038), .B2(KEYINPUT50), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(G2090), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n996), .ZN(new_n1041));
  AOI211_X1 g616(.A(new_n996), .B(G1384), .C1(new_n495), .C2(new_n505), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n998), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1040), .B1(new_n723), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G8), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1034), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n723), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1038), .A2(KEYINPUT50), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1036), .B1(new_n1050), .B2(new_n1016), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1048), .B1(G2090), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1034), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(G8), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1032), .A2(new_n1047), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT125), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n998), .B1(new_n1016), .B2(KEYINPUT45), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n869), .A2(KEYINPUT70), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n495), .A2(new_n505), .A3(new_n506), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1384), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1060), .B1(new_n1063), .B2(KEYINPUT45), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1059), .B1(new_n1064), .B2(G1966), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1038), .A2(new_n996), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT117), .B(new_n772), .C1(new_n1066), .C2(new_n1060), .ZN(new_n1067));
  INV_X1    g642(.A(G2084), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1049), .A2(new_n1068), .A3(new_n1051), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1065), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(G8), .B1(new_n1070), .B2(G286), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT51), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n1070), .B2(G286), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1072), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1032), .A2(new_n1047), .A3(new_n1055), .A4(KEYINPUT125), .ZN(new_n1076));
  XNOR2_X1  g651(.A(G301), .B(KEYINPUT54), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1044), .B2(G2078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT122), .B(G1961), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1052), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1064), .A2(KEYINPUT53), .A3(new_n798), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n995), .A2(new_n996), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n798), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n470), .A2(new_n471), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1086), .A2(KEYINPUT123), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n464), .B1(new_n1086), .B2(KEYINPUT123), .ZN(new_n1088));
  AOI211_X1 g663(.A(new_n480), .B(new_n1085), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1043), .A2(new_n1084), .A3(new_n1089), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1090), .A2(KEYINPUT124), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1077), .B1(new_n1090), .B2(KEYINPUT124), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1081), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1077), .A2(new_n1083), .B1(new_n1093), .B2(new_n1079), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1058), .A2(new_n1075), .A3(new_n1076), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n998), .A2(new_n768), .ZN(new_n1099));
  AOI211_X1 g674(.A(new_n1042), .B(new_n1099), .C1(new_n1038), .C2(new_n996), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT58), .B(G1341), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n1016), .B2(new_n998), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1102), .B(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1098), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1102), .B(KEYINPUT119), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1099), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1041), .A2(new_n1043), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(new_n1108), .A3(KEYINPUT120), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1097), .B1(new_n1110), .B2(new_n568), .ZN(new_n1111));
  AOI211_X1 g686(.A(KEYINPUT59), .B(new_n567), .C1(new_n1105), .C2(new_n1109), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1956), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1039), .A2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1041), .A2(new_n998), .A3(new_n1043), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n580), .B(KEYINPUT118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT57), .B1(new_n584), .B2(new_n586), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1119), .A2(new_n1120), .B1(KEYINPUT57), .B2(G299), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1121), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(KEYINPUT61), .A3(new_n1124), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1096), .B1(new_n1113), .B2(new_n1129), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1106), .A2(new_n1108), .A3(KEYINPUT120), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT120), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n568), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT59), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1110), .A2(new_n1097), .A3(new_n568), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1136), .A2(KEYINPUT121), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1017), .A2(G2067), .ZN(new_n1138));
  INV_X1    g713(.A(G1348), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1052), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT60), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(new_n630), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(KEYINPUT60), .B2(new_n1140), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1130), .A2(new_n1137), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1123), .B1(new_n909), .B2(new_n1140), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1124), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1095), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1148));
  NOR2_X1   g723(.A1(G288), .A2(G1976), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1148), .A2(new_n1149), .B1(new_n1022), .B2(new_n726), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1032), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1150), .A2(new_n1029), .B1(new_n1151), .B2(new_n1055), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT63), .ZN(new_n1153));
  NOR2_X1   g728(.A1(G286), .A2(new_n1046), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1070), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1056), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1070), .A2(KEYINPUT63), .A3(new_n1154), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1053), .A2(G8), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1157), .B1(new_n1034), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1159), .A2(new_n1055), .A3(new_n1032), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1152), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1075), .A2(KEYINPUT62), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1072), .B(new_n1163), .C1(new_n1071), .C2(new_n1074), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1058), .A2(G171), .A3(new_n1076), .A4(new_n1083), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1161), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1012), .B1(new_n1147), .B2(new_n1167), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n736), .A2(new_n744), .A3(new_n740), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1008), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n819), .A2(new_n1005), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n999), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT46), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n765), .B(new_n1006), .C1(new_n1176), .C2(G1996), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1176), .B1(new_n999), .B2(G1996), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1177), .A2(new_n1000), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1180), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT47), .ZN(new_n1182));
  NOR3_X1   g757(.A1(G290), .A2(new_n999), .A3(G1986), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT48), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1182), .B1(new_n1010), .B2(new_n1184), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1174), .A2(new_n1175), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1168), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  OR4_X1    g762(.A1(new_n462), .A2(G229), .A3(G401), .A4(G227), .ZN(new_n1189));
  AOI21_X1  g763(.A(new_n1189), .B1(new_n902), .B2(new_n903), .ZN(new_n1190));
  AND2_X1   g764(.A1(new_n1190), .A2(new_n978), .ZN(G308));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n978), .ZN(G225));
endmodule


