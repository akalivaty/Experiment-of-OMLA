//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182, new_n1183, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G101), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  NOR3_X1   g042(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(new_n466), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n470), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n475), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n479), .B1(new_n469), .B2(G125), .ZN(new_n480));
  NOR3_X1   g055(.A1(new_n480), .A2(KEYINPUT68), .A3(new_n471), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n478), .A2(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(new_n472), .A2(new_n473), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT69), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n469), .A2(new_n485), .A3(new_n461), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n471), .A2(G112), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n471), .A2(new_n483), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n490), .A2(new_n492), .B1(new_n493), .B2(G124), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  OAI21_X1  g074(.A(G2105), .B1(new_n499), .B2(G114), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT70), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(G126), .B(G2105), .C1(new_n472), .C2(new_n473), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(new_n461), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(G138), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT4), .B1(new_n509), .B2(new_n483), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n471), .A2(new_n469), .A3(new_n511), .A4(G138), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n505), .B1(new_n510), .B2(new_n512), .ZN(G164));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT72), .B1(new_n514), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n514), .A2(G543), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n519), .A2(G88), .A3(new_n520), .A4(new_n523), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n517), .B1(new_n521), .B2(new_n522), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n525), .A2(KEYINPUT71), .A3(G50), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT71), .B1(new_n525), .B2(G50), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n519), .A2(G62), .A3(new_n520), .ZN(new_n530));
  NAND2_X1  g105(.A1(G75), .A2(G543), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT73), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n529), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n528), .A2(new_n533), .ZN(G166));
  AND2_X1   g109(.A1(new_n519), .A2(new_n520), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n535), .A2(G63), .A3(G651), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n519), .A2(new_n520), .A3(new_n523), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G89), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n541));
  AOI22_X1  g116(.A1(G51), .A2(new_n525), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n536), .A2(new_n538), .A3(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  AOI22_X1  g119(.A1(new_n535), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n529), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n525), .A2(G52), .ZN(new_n547));
  INV_X1    g122(.A(new_n537), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n546), .A2(new_n550), .ZN(G171));
  AOI22_X1  g126(.A1(new_n535), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n554), .A2(G651), .A3(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n537), .A2(G81), .B1(G43), .B2(new_n525), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT75), .Z(G188));
  NAND4_X1  g140(.A1(new_n519), .A2(G91), .A3(new_n520), .A4(new_n523), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n525), .A2(new_n567), .A3(G53), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n567), .B1(new_n525), .B2(G53), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n519), .A2(G65), .A3(new_n520), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n529), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  INV_X1    g152(.A(G166), .ZN(G303));
  OAI21_X1  g153(.A(G651), .B1(new_n535), .B2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n537), .A2(G87), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n525), .A2(G49), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n525), .A2(new_n583), .A3(G48), .ZN(new_n584));
  AND2_X1   g159(.A1(KEYINPUT6), .A2(G651), .ZN(new_n585));
  NOR2_X1   g160(.A1(KEYINPUT6), .A2(G651), .ZN(new_n586));
  OAI211_X1 g161(.A(G48), .B(G543), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT76), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n537), .A2(G86), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n519), .A2(G61), .A3(new_n520), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n535), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n529), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n525), .A2(G47), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n548), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n525), .A2(G54), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n535), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n529), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT77), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n537), .A2(G92), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT10), .Z(new_n608));
  AND2_X1   g183(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n602), .B1(new_n609), .B2(G868), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(KEYINPUT78), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n612), .A2(KEYINPUT78), .ZN(new_n614));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(G299), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n613), .B1(new_n614), .B2(new_n616), .ZN(G297));
  AOI21_X1  g192(.A(new_n613), .B1(new_n614), .B2(new_n616), .ZN(G280));
  XOR2_X1   g193(.A(KEYINPUT79), .B(G559), .Z(new_n619));
  OAI21_X1  g194(.A(new_n609), .B1(G860), .B2(new_n619), .ZN(G148));
  NOR2_X1   g195(.A1(new_n558), .A2(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n609), .A2(new_n619), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(KEYINPUT80), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT80), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n609), .A2(new_n624), .A3(new_n619), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n621), .B1(new_n627), .B2(G868), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g204(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT13), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n493), .A2(G123), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT81), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n488), .A2(G135), .ZN(new_n636));
  OAI221_X1 g211(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n471), .C2(G111), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(G2096), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n639), .A3(new_n640), .ZN(G156));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT82), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT83), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(G14), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(G401));
  INV_X1    g234(.A(KEYINPUT18), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n660), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2100), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n663), .B2(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2096), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(new_n670), .ZN(G227));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n676), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n680), .A2(KEYINPUT20), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(KEYINPUT20), .ZN(new_n682));
  OAI221_X1 g257(.A(new_n677), .B1(new_n674), .B2(new_n678), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G229));
  MUX2_X1   g264(.A(G6), .B(G305), .S(G16), .Z(new_n690));
  XOR2_X1   g265(.A(KEYINPUT32), .B(G1981), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G23), .ZN(new_n694));
  INV_X1    g269(.A(G288), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(new_n693), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT33), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT86), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n696), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n693), .A2(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n693), .ZN(new_n701));
  INV_X1    g276(.A(G1971), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n692), .A2(new_n699), .A3(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT85), .B(KEYINPUT34), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G25), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n488), .A2(G131), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n471), .A2(G107), .ZN(new_n712));
  OAI21_X1  g287(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n712), .A2(new_n714), .B1(new_n493), .B2(G119), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n710), .B1(new_n717), .B2(new_n709), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G1986), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n600), .A2(new_n693), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n693), .B2(G24), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n720), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n721), .B2(new_n723), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n707), .A2(new_n708), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT87), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(KEYINPUT36), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n726), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G29), .A2(G32), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT98), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT26), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n493), .A2(G129), .ZN(new_n734));
  INV_X1    g309(.A(G105), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n462), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n488), .A2(G141), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(KEYINPUT97), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(KEYINPUT97), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n733), .B(new_n736), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT99), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n730), .B1(new_n743), .B2(G29), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT27), .B(G1996), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n693), .A2(G4), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n609), .B2(new_n693), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n744), .A2(new_n745), .B1(G1348), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G19), .ZN(new_n749));
  OR3_X1    g324(.A1(new_n749), .A2(KEYINPUT88), .A3(G16), .ZN(new_n750));
  OAI21_X1  g325(.A(KEYINPUT88), .B1(new_n749), .B2(G16), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n750), .B(new_n751), .C1(new_n559), .C2(new_n693), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(G1341), .Z(new_n753));
  OAI211_X1 g328(.A(new_n748), .B(new_n753), .C1(new_n745), .C2(new_n744), .ZN(new_n754));
  NOR2_X1   g329(.A1(G29), .A2(G33), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT91), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT92), .B(KEYINPUT25), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT93), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(new_n471), .ZN(new_n762));
  INV_X1    g337(.A(G139), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n760), .B(new_n762), .C1(new_n763), .C2(new_n487), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n756), .B1(new_n764), .B2(new_n709), .ZN(new_n765));
  INV_X1    g340(.A(G2072), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT94), .Z(new_n768));
  INV_X1    g343(.A(G34), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(KEYINPUT24), .ZN(new_n770));
  AOI21_X1  g345(.A(G29), .B1(new_n769), .B2(KEYINPUT24), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(KEYINPUT95), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(KEYINPUT95), .B2(new_n771), .ZN(new_n773));
  INV_X1    g348(.A(G160), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n709), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT96), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2084), .ZN(new_n777));
  NAND2_X1  g352(.A1(G171), .A2(G16), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G5), .B2(G16), .ZN(new_n779));
  INV_X1    g354(.A(G1961), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(G164), .A2(G29), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G27), .B2(G29), .ZN(new_n783));
  INV_X1    g358(.A(G2078), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n638), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G29), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT31), .B(G11), .Z(new_n788));
  XOR2_X1   g363(.A(KEYINPUT101), .B(G28), .Z(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(KEYINPUT30), .ZN(new_n790));
  AOI21_X1  g365(.A(G29), .B1(new_n789), .B2(KEYINPUT30), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n781), .A2(new_n785), .A3(new_n787), .A4(new_n792), .ZN(new_n793));
  OAI22_X1  g368(.A1(new_n765), .A2(new_n766), .B1(new_n779), .B2(new_n780), .ZN(new_n794));
  OR4_X1    g369(.A1(new_n768), .A2(new_n777), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(G168), .A2(G16), .ZN(new_n796));
  NOR2_X1   g371(.A1(G16), .A2(G21), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(KEYINPUT100), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(KEYINPUT100), .B2(new_n796), .ZN(new_n799));
  INV_X1    g374(.A(G1966), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n709), .A2(G26), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT28), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n493), .A2(G128), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT89), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n488), .A2(G140), .ZN(new_n806));
  NOR2_X1   g381(.A1(G104), .A2(G2105), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT90), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n808), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n805), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n803), .B1(new_n810), .B2(G29), .ZN(new_n811));
  INV_X1    g386(.A(G2067), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n801), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n709), .A2(G35), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT102), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G162), .B2(new_n709), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT103), .B(KEYINPUT29), .ZN(new_n818));
  INV_X1    g393(.A(G2090), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n817), .A2(new_n821), .B1(new_n783), .B2(new_n784), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n693), .A2(G20), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT23), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n575), .B2(new_n693), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1956), .ZN(new_n826));
  AOI211_X1 g401(.A(new_n822), .B(new_n826), .C1(new_n817), .C2(new_n821), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n814), .B(new_n827), .C1(G1348), .C2(new_n747), .ZN(new_n828));
  NOR4_X1   g403(.A1(new_n729), .A2(new_n754), .A3(new_n795), .A4(new_n828), .ZN(G311));
  INV_X1    g404(.A(G311), .ZN(G150));
  AOI22_X1  g405(.A1(new_n535), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(new_n529), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n525), .A2(G55), .ZN(new_n833));
  INV_X1    g408(.A(G93), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n548), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G860), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT105), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n609), .A2(G559), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT104), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n559), .A2(new_n836), .ZN(new_n846));
  INV_X1    g421(.A(new_n836), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n558), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n844), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n849), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n841), .B1(new_n855), .B2(KEYINPUT39), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n857));
  AOI211_X1 g432(.A(KEYINPUT105), .B(new_n857), .C1(new_n851), .C2(new_n854), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n837), .B1(new_n855), .B2(KEYINPUT39), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n840), .B1(new_n859), .B2(new_n860), .ZN(G145));
  NAND2_X1  g436(.A1(new_n488), .A2(G142), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT108), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n471), .A2(G118), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AOI22_X1  g441(.A1(new_n864), .A2(new_n866), .B1(new_n493), .B2(G130), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT109), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(new_n631), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n631), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n717), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n869), .B(new_n631), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n716), .ZN(new_n874));
  INV_X1    g449(.A(new_n764), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n742), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n740), .A2(new_n764), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n510), .A2(new_n512), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n503), .A2(new_n504), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT107), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT107), .B1(new_n879), .B2(new_n880), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n810), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n878), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n885), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n876), .A2(new_n887), .A3(new_n877), .ZN(new_n888));
  AND4_X1   g463(.A1(new_n872), .A2(new_n874), .A3(new_n886), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT111), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n495), .B(G160), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n786), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(KEYINPUT112), .Z(new_n893));
  NAND3_X1  g468(.A1(new_n874), .A2(KEYINPUT111), .A3(new_n872), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n886), .A2(new_n888), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(KEYINPUT110), .B(G37), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n872), .A2(new_n874), .B1(new_n886), .B2(new_n888), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n892), .B1(new_n889), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g477(.A1(new_n627), .A2(new_n850), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n850), .B1(new_n623), .B2(new_n625), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n606), .A2(new_n608), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n575), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT41), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n609), .A2(new_n575), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n906), .A2(G299), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n903), .A2(new_n905), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n626), .A2(new_n849), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(new_n904), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n914), .B1(new_n916), .B2(new_n907), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n600), .B(G288), .ZN(new_n919));
  XNOR2_X1  g494(.A(G166), .B(G305), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n919), .B(new_n920), .Z(new_n921));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n914), .B(new_n922), .C1(new_n907), .C2(new_n916), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n918), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n921), .B1(new_n918), .B2(new_n923), .ZN(new_n925));
  OAI21_X1  g500(.A(G868), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n847), .A2(new_n615), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(G295));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n927), .ZN(G331));
  NAND3_X1  g504(.A1(new_n846), .A2(G301), .A3(new_n848), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(G301), .B1(new_n846), .B2(new_n848), .ZN(new_n932));
  OAI21_X1  g507(.A(G286), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n932), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n934), .A2(G168), .A3(new_n930), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n913), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n907), .B1(new_n933), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n921), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n921), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n913), .A2(new_n933), .A3(new_n935), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n933), .A2(new_n935), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n939), .B(new_n940), .C1(new_n941), .C2(new_n907), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G37), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT43), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  INV_X1    g521(.A(new_n898), .ZN(new_n947));
  AOI211_X1 g522(.A(new_n946), .B(new_n947), .C1(new_n938), .C2(new_n942), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT44), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n946), .B1(new_n943), .B2(new_n944), .ZN(new_n950));
  AOI211_X1 g525(.A(KEYINPUT43), .B(new_n947), .C1(new_n938), .C2(new_n942), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n949), .B1(new_n952), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g528(.A(KEYINPUT113), .ZN(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n884), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n879), .A2(new_n880), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n959), .A2(new_n954), .A3(new_n955), .A4(new_n881), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT68), .B1(new_n480), .B2(new_n471), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n474), .A2(new_n475), .ZN(new_n964));
  INV_X1    g539(.A(new_n471), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n477), .A3(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n963), .A2(G40), .A3(new_n966), .A4(new_n470), .ZN(new_n967));
  OR3_X1    g542(.A1(new_n956), .A2(new_n962), .A3(new_n967), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n968), .A2(G1986), .A3(G290), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n969), .B(KEYINPUT48), .Z(new_n970));
  XNOR2_X1  g545(.A(new_n968), .B(KEYINPUT114), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n716), .B(new_n719), .Z(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n810), .B(new_n812), .ZN(new_n974));
  INV_X1    g549(.A(G1996), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(new_n975), .B2(new_n740), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n968), .A2(G1996), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n971), .A2(new_n976), .B1(new_n743), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n970), .A2(new_n973), .A3(new_n978), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n977), .B(KEYINPUT46), .Z(new_n980));
  NAND2_X1  g555(.A1(new_n974), .A2(new_n740), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n971), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n983), .A2(KEYINPUT47), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(KEYINPUT47), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n979), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n717), .A2(new_n719), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT126), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n978), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(G2067), .B2(new_n810), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n986), .B1(new_n971), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n957), .A2(new_n955), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n967), .B1(new_n993), .B2(new_n961), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n961), .A2(G1384), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n957), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(G1966), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G2084), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n999));
  INV_X1    g574(.A(G40), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n478), .A2(new_n481), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n957), .A2(new_n1002), .A3(new_n955), .ZN(new_n1003));
  AND4_X1   g578(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(G8), .B1(new_n997), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n992), .B1(new_n1005), .B2(KEYINPUT122), .ZN(new_n1006));
  OAI21_X1  g581(.A(G286), .B1(new_n997), .B2(new_n1004), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .A4(new_n998), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n961), .B1(G164), .B2(G1384), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1009), .A2(new_n1001), .A3(new_n996), .ZN(new_n1010));
  OAI211_X1 g585(.A(G168), .B(new_n1008), .C1(new_n1010), .C2(G1966), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1007), .A2(G8), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G8), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(new_n1001), .A3(new_n996), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n1015), .A2(new_n998), .B1(new_n1016), .B2(new_n800), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1014), .B1(new_n1017), .B2(G168), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT122), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1008), .B1(new_n1010), .B2(G1966), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n1020), .B2(G8), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1018), .B1(new_n1021), .B2(new_n992), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1013), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(G8), .B1(new_n993), .B2(new_n967), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT49), .ZN(new_n1025));
  INV_X1    g600(.A(G1981), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n589), .A2(new_n593), .A3(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n519), .A2(G86), .A3(new_n520), .A4(new_n523), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n583), .B1(new_n525), .B2(G48), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n587), .A2(KEYINPUT76), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n529), .B1(new_n590), .B2(new_n591), .ZN(new_n1032));
  OAI21_X1  g607(.A(G1981), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1027), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1024), .B1(new_n1025), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1027), .A2(new_n1033), .A3(KEYINPUT49), .ZN(new_n1036));
  NOR2_X1   g611(.A1(G164), .A2(G1384), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1001), .A2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n579), .A2(new_n580), .A3(G1976), .A4(new_n581), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(G8), .A3(new_n1039), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1035), .A2(new_n1036), .B1(KEYINPUT52), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(G166), .B2(new_n1014), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT55), .B(G8), .C1(new_n528), .C2(new_n533), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n959), .A2(new_n881), .A3(new_n995), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1971), .B1(new_n994), .B2(new_n1046), .ZN(new_n1047));
  AND4_X1   g622(.A1(new_n819), .A2(new_n999), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1048));
  OAI211_X1 g623(.A(G8), .B(new_n1045), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1024), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1039), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1041), .A2(new_n1049), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1045), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT116), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1056));
  INV_X1    g631(.A(new_n995), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n882), .A2(new_n883), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1009), .A2(new_n1001), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n702), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .A4(new_n819), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1056), .A2(new_n1063), .A3(G8), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1054), .B1(new_n1055), .B2(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1023), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT120), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .A4(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n780), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n994), .A2(new_n784), .A3(new_n1046), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1010), .A2(KEYINPUT53), .A3(new_n784), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1071), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G171), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n471), .B1(new_n964), .B2(KEYINPUT123), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(KEYINPUT123), .B2(new_n964), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n470), .A2(KEYINPUT53), .A3(G40), .A4(new_n784), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1046), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n956), .B2(new_n962), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1083), .A2(G301), .A3(new_n1074), .A4(new_n1071), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1077), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1071), .A2(new_n1074), .A3(G301), .A4(new_n1075), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1083), .A2(new_n1074), .A3(new_n1071), .ZN(new_n1089));
  OAI211_X1 g664(.A(KEYINPUT54), .B(new_n1088), .C1(new_n1089), .C2(G301), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1066), .A2(KEYINPUT124), .A3(new_n1087), .A4(new_n1090), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT118), .B(G1956), .Z(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1067), .A2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT56), .B(G2072), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1046), .A2(new_n1001), .A3(new_n1009), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n1097));
  INV_X1    g672(.A(new_n570), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1098), .A2(new_n568), .B1(new_n537), .B2(G91), .ZN(new_n1099));
  INV_X1    g674(.A(new_n574), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1097), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n571), .A2(KEYINPUT57), .A3(new_n574), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1094), .A2(new_n1096), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1094), .A2(new_n1096), .A3(KEYINPUT119), .A4(new_n1103), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1103), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1103), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT121), .B1(new_n1117), .B2(KEYINPUT61), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1111), .A2(KEYINPUT61), .A3(new_n1104), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n994), .A2(new_n975), .A3(new_n1046), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1038), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT58), .B(G1341), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n559), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n559), .A3(KEYINPUT59), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1119), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1348), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1068), .A2(new_n1129), .A3(new_n1070), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1121), .A2(new_n812), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n906), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n609), .A2(KEYINPUT60), .A3(new_n1131), .A4(new_n1130), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1115), .A2(new_n1118), .A3(new_n1128), .A4(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n906), .B1(new_n1131), .B2(new_n1130), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1108), .B1(new_n1139), .B2(new_n1116), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1087), .A2(new_n1090), .A3(new_n1023), .A4(new_n1065), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1091), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1034), .A2(new_n1025), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1146), .A2(new_n1050), .A3(new_n1036), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1147), .A2(new_n1051), .A3(new_n695), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1024), .B1(new_n1148), .B2(new_n1027), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1040), .A2(KEYINPUT52), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1147), .A2(new_n1150), .A3(new_n1053), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1151), .A2(new_n1049), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT115), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1005), .A2(G286), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT63), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1045), .B1(new_n1158), .B2(G8), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1157), .A2(new_n1159), .A3(new_n1054), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1064), .A2(new_n1055), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1041), .A2(new_n1049), .A3(new_n1053), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1161), .A2(new_n1162), .A3(new_n1156), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT63), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT117), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1160), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1163), .A2(KEYINPUT117), .A3(new_n1164), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1155), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1145), .A2(KEYINPUT125), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT125), .B1(new_n1145), .B2(new_n1169), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1023), .A2(KEYINPUT62), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1023), .A2(KEYINPUT62), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1065), .A2(G171), .A3(new_n1076), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1170), .A2(new_n1171), .A3(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n600), .B(G1986), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n978), .B(new_n973), .C1(new_n968), .C2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n991), .B1(new_n1176), .B2(new_n1178), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g754(.A1(new_n459), .A2(G227), .ZN(new_n1181));
  NOR3_X1   g755(.A1(G229), .A2(G401), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n1183));
  XNOR2_X1  g757(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  OAI211_X1 g758(.A(new_n1184), .B(new_n901), .C1(new_n950), .C2(new_n951), .ZN(G225));
  INV_X1    g759(.A(G225), .ZN(G308));
endmodule


