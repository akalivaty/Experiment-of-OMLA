

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595;

  XNOR2_X1 U327 ( .A(n402), .B(n401), .ZN(n543) );
  XNOR2_X1 U328 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n401) );
  XNOR2_X1 U329 ( .A(n314), .B(KEYINPUT41), .ZN(n315) );
  INV_X1 U330 ( .A(KEYINPUT73), .ZN(n304) );
  XNOR2_X1 U331 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U332 ( .A(n307), .B(n306), .ZN(n311) );
  XNOR2_X1 U333 ( .A(n388), .B(n315), .ZN(n392) );
  NOR2_X1 U334 ( .A1(n485), .A2(n465), .ZN(n574) );
  XOR2_X1 U335 ( .A(n332), .B(n403), .Z(n544) );
  XNOR2_X1 U336 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U337 ( .A(n472), .B(n471), .ZN(G1351GAT) );
  INV_X1 U338 ( .A(G92GAT), .ZN(n295) );
  NAND2_X1 U339 ( .A1(n295), .A2(G64GAT), .ZN(n298) );
  INV_X1 U340 ( .A(G64GAT), .ZN(n296) );
  NAND2_X1 U341 ( .A1(n296), .A2(G92GAT), .ZN(n297) );
  NAND2_X1 U342 ( .A1(n298), .A2(n297), .ZN(n300) );
  XNOR2_X1 U343 ( .A(G176GAT), .B(G204GAT), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n408) );
  XOR2_X1 U345 ( .A(G99GAT), .B(G85GAT), .Z(n380) );
  XOR2_X1 U346 ( .A(n408), .B(n380), .Z(n302) );
  NAND2_X1 U347 ( .A1(G230GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n307) );
  XNOR2_X1 U349 ( .A(G106GAT), .B(G78GAT), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n303), .B(G148GAT), .ZN(n456) );
  XNOR2_X1 U351 ( .A(n456), .B(KEYINPUT74), .ZN(n305) );
  XOR2_X1 U352 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n309) );
  XNOR2_X1 U353 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n308) );
  XOR2_X1 U354 ( .A(n309), .B(n308), .Z(n310) );
  XNOR2_X1 U355 ( .A(n311), .B(n310), .ZN(n313) );
  XOR2_X1 U356 ( .A(G120GAT), .B(G71GAT), .Z(n316) );
  XOR2_X1 U357 ( .A(G57GAT), .B(KEYINPUT13), .Z(n349) );
  XNOR2_X1 U358 ( .A(n316), .B(n349), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n313), .B(n312), .ZN(n388) );
  INV_X1 U360 ( .A(KEYINPUT65), .ZN(n314) );
  XNOR2_X1 U361 ( .A(KEYINPUT108), .B(n392), .ZN(n550) );
  XOR2_X1 U362 ( .A(G15GAT), .B(G127GAT), .Z(n350) );
  XOR2_X1 U363 ( .A(n316), .B(n350), .Z(n318) );
  NAND2_X1 U364 ( .A1(G227GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U366 ( .A(G134GAT), .B(KEYINPUT0), .Z(n439) );
  XOR2_X1 U367 ( .A(n319), .B(n439), .Z(n327) );
  XOR2_X1 U368 ( .A(KEYINPUT20), .B(G99GAT), .Z(n321) );
  XNOR2_X1 U369 ( .A(G43GAT), .B(G190GAT), .ZN(n320) );
  XNOR2_X1 U370 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U371 ( .A(G176GAT), .B(KEYINPUT84), .Z(n323) );
  XNOR2_X1 U372 ( .A(G169GAT), .B(G113GAT), .ZN(n322) );
  XNOR2_X1 U373 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n332) );
  XOR2_X1 U376 ( .A(G183GAT), .B(KEYINPUT85), .Z(n329) );
  XNOR2_X1 U377 ( .A(KEYINPUT18), .B(KEYINPUT86), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n331) );
  XOR2_X1 U379 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n330) );
  XNOR2_X1 U380 ( .A(n331), .B(n330), .ZN(n403) );
  INV_X1 U381 ( .A(n544), .ZN(n485) );
  XOR2_X1 U382 ( .A(KEYINPUT7), .B(KEYINPUT71), .Z(n334) );
  XNOR2_X1 U383 ( .A(G43GAT), .B(G29GAT), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U385 ( .A(KEYINPUT8), .B(n335), .Z(n386) );
  XOR2_X1 U386 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n337) );
  XNOR2_X1 U387 ( .A(G197GAT), .B(G15GAT), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U389 ( .A(G141GAT), .B(G22GAT), .Z(n453) );
  XNOR2_X1 U390 ( .A(n338), .B(n453), .ZN(n342) );
  XOR2_X1 U391 ( .A(G113GAT), .B(G1GAT), .Z(n440) );
  XOR2_X1 U392 ( .A(KEYINPUT29), .B(n440), .Z(n340) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U396 ( .A(G169GAT), .B(G8GAT), .Z(n413) );
  XOR2_X1 U397 ( .A(n343), .B(n413), .Z(n345) );
  XNOR2_X1 U398 ( .A(G50GAT), .B(G36GAT), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n386), .B(n346), .ZN(n581) );
  XOR2_X1 U401 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n348) );
  XNOR2_X1 U402 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n354) );
  XOR2_X1 U404 ( .A(n349), .B(G211GAT), .Z(n352) );
  XNOR2_X1 U405 ( .A(G22GAT), .B(n350), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U407 ( .A(n354), .B(n353), .Z(n356) );
  NAND2_X1 U408 ( .A1(G231GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U410 ( .A(G78GAT), .B(G155GAT), .Z(n358) );
  XNOR2_X1 U411 ( .A(G183GAT), .B(G71GAT), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U413 ( .A(n360), .B(n359), .Z(n368) );
  XOR2_X1 U414 ( .A(KEYINPUT82), .B(KEYINPUT12), .Z(n362) );
  XNOR2_X1 U415 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U417 ( .A(KEYINPUT77), .B(G64GAT), .Z(n364) );
  XNOR2_X1 U418 ( .A(G8GAT), .B(G1GAT), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U421 ( .A(n368), .B(n367), .ZN(n503) );
  XOR2_X1 U422 ( .A(G92GAT), .B(G106GAT), .Z(n370) );
  XNOR2_X1 U423 ( .A(G134GAT), .B(G218GAT), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U425 ( .A(KEYINPUT69), .B(KEYINPUT9), .Z(n372) );
  XNOR2_X1 U426 ( .A(KEYINPUT76), .B(KEYINPUT67), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U428 ( .A(n374), .B(n373), .Z(n379) );
  XOR2_X1 U429 ( .A(KEYINPUT11), .B(KEYINPUT68), .Z(n376) );
  NAND2_X1 U430 ( .A1(G232GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U432 ( .A(KEYINPUT10), .B(n377), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n381) );
  XOR2_X1 U434 ( .A(n381), .B(n380), .Z(n384) );
  XNOR2_X1 U435 ( .A(G50GAT), .B(KEYINPUT75), .ZN(n382) );
  XNOR2_X1 U436 ( .A(n382), .B(G162GAT), .ZN(n447) );
  XOR2_X1 U437 ( .A(G36GAT), .B(G190GAT), .Z(n409) );
  XNOR2_X1 U438 ( .A(n447), .B(n409), .ZN(n383) );
  XNOR2_X1 U439 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U440 ( .A(n386), .B(n385), .Z(n394) );
  XOR2_X1 U441 ( .A(KEYINPUT36), .B(n394), .Z(n592) );
  NOR2_X1 U442 ( .A1(n503), .A2(n592), .ZN(n387) );
  XNOR2_X1 U443 ( .A(KEYINPUT45), .B(n387), .ZN(n389) );
  NAND2_X1 U444 ( .A1(n389), .A2(n388), .ZN(n390) );
  NOR2_X1 U445 ( .A1(n581), .A2(n390), .ZN(n391) );
  XOR2_X1 U446 ( .A(KEYINPUT115), .B(n391), .Z(n400) );
  NAND2_X1 U447 ( .A1(n581), .A2(n392), .ZN(n393) );
  XNOR2_X1 U448 ( .A(KEYINPUT46), .B(n393), .ZN(n397) );
  INV_X1 U449 ( .A(n394), .ZN(n395) );
  INV_X1 U450 ( .A(n395), .ZN(n570) );
  INV_X1 U451 ( .A(n503), .ZN(n589) );
  NOR2_X1 U452 ( .A1(n570), .A2(n589), .ZN(n396) );
  AND2_X1 U453 ( .A1(n397), .A2(n396), .ZN(n398) );
  XOR2_X1 U454 ( .A(n398), .B(KEYINPUT47), .Z(n399) );
  NOR2_X1 U455 ( .A1(n400), .A2(n399), .ZN(n402) );
  INV_X1 U456 ( .A(n403), .ZN(n407) );
  XOR2_X1 U457 ( .A(KEYINPUT88), .B(G218GAT), .Z(n405) );
  XNOR2_X1 U458 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U460 ( .A(G197GAT), .B(n406), .Z(n459) );
  XNOR2_X1 U461 ( .A(n407), .B(n459), .ZN(n417) );
  XOR2_X1 U462 ( .A(n408), .B(n409), .Z(n411) );
  NAND2_X1 U463 ( .A1(G226GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U464 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U465 ( .A(n412), .B(KEYINPUT98), .Z(n415) );
  XNOR2_X1 U466 ( .A(n413), .B(KEYINPUT99), .ZN(n414) );
  XNOR2_X1 U467 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U468 ( .A(n417), .B(n416), .ZN(n531) );
  XNOR2_X1 U469 ( .A(n531), .B(KEYINPUT121), .ZN(n418) );
  NOR2_X1 U470 ( .A1(n543), .A2(n418), .ZN(n419) );
  XNOR2_X1 U471 ( .A(n419), .B(KEYINPUT54), .ZN(n445) );
  XOR2_X1 U472 ( .A(G57GAT), .B(G148GAT), .Z(n421) );
  XNOR2_X1 U473 ( .A(G120GAT), .B(G127GAT), .ZN(n420) );
  XNOR2_X1 U474 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U475 ( .A(G85GAT), .B(G162GAT), .Z(n423) );
  XNOR2_X1 U476 ( .A(G29GAT), .B(G141GAT), .ZN(n422) );
  XNOR2_X1 U477 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n444) );
  XOR2_X1 U479 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n427) );
  XNOR2_X1 U480 ( .A(KEYINPUT5), .B(KEYINPUT97), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U482 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n429) );
  XNOR2_X1 U483 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U485 ( .A(n431), .B(n430), .Z(n436) );
  XOR2_X1 U486 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n433) );
  NAND2_X1 U487 ( .A1(G225GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U489 ( .A(KEYINPUT92), .B(n434), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U491 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n437), .B(KEYINPUT2), .ZN(n458) );
  XOR2_X1 U493 ( .A(n438), .B(n458), .Z(n442) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n482) );
  NAND2_X1 U497 ( .A1(n445), .A2(n482), .ZN(n446) );
  XNOR2_X1 U498 ( .A(n446), .B(KEYINPUT66), .ZN(n580) );
  XOR2_X1 U499 ( .A(n447), .B(KEYINPUT22), .Z(n449) );
  NAND2_X1 U500 ( .A1(G228GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n463) );
  XOR2_X1 U502 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n451) );
  XNOR2_X1 U503 ( .A(G204GAT), .B(KEYINPUT87), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U505 ( .A(n452), .B(KEYINPUT89), .Z(n455) );
  XNOR2_X1 U506 ( .A(n453), .B(KEYINPUT23), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(n457) );
  XOR2_X1 U508 ( .A(n457), .B(n456), .Z(n461) );
  XNOR2_X1 U509 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U510 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U511 ( .A(n463), .B(n462), .ZN(n484) );
  NOR2_X1 U512 ( .A1(n580), .A2(n484), .ZN(n464) );
  XNOR2_X1 U513 ( .A(n464), .B(KEYINPUT55), .ZN(n465) );
  NAND2_X1 U514 ( .A1(n550), .A2(n574), .ZN(n468) );
  XOR2_X1 U515 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n466) );
  XNOR2_X1 U516 ( .A(n466), .B(G176GAT), .ZN(n467) );
  XNOR2_X1 U517 ( .A(n468), .B(n467), .ZN(G1349GAT) );
  NAND2_X1 U518 ( .A1(n574), .A2(n570), .ZN(n472) );
  XOR2_X1 U519 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n470) );
  INV_X1 U520 ( .A(G190GAT), .ZN(n469) );
  XOR2_X1 U521 ( .A(KEYINPUT103), .B(KEYINPUT34), .Z(n493) );
  NAND2_X1 U522 ( .A1(n388), .A2(n581), .ZN(n506) );
  XOR2_X1 U523 ( .A(KEYINPUT25), .B(KEYINPUT101), .Z(n473) );
  XNOR2_X1 U524 ( .A(KEYINPUT100), .B(n473), .ZN(n476) );
  AND2_X1 U525 ( .A1(n544), .A2(n531), .ZN(n474) );
  NOR2_X1 U526 ( .A1(n484), .A2(n474), .ZN(n475) );
  XNOR2_X1 U527 ( .A(n476), .B(n475), .ZN(n479) );
  NAND2_X1 U528 ( .A1(n484), .A2(n485), .ZN(n477) );
  XNOR2_X1 U529 ( .A(n477), .B(KEYINPUT26), .ZN(n579) );
  INV_X1 U530 ( .A(n579), .ZN(n559) );
  XNOR2_X1 U531 ( .A(n531), .B(KEYINPUT27), .ZN(n483) );
  NAND2_X1 U532 ( .A1(n559), .A2(n483), .ZN(n478) );
  NAND2_X1 U533 ( .A1(n479), .A2(n478), .ZN(n480) );
  NAND2_X1 U534 ( .A1(n482), .A2(n480), .ZN(n481) );
  XOR2_X1 U535 ( .A(KEYINPUT102), .B(n481), .Z(n488) );
  INV_X1 U536 ( .A(n482), .ZN(n529) );
  NAND2_X1 U537 ( .A1(n529), .A2(n483), .ZN(n542) );
  XOR2_X1 U538 ( .A(KEYINPUT28), .B(n484), .Z(n547) );
  NAND2_X1 U539 ( .A1(n485), .A2(n547), .ZN(n486) );
  NOR2_X1 U540 ( .A1(n542), .A2(n486), .ZN(n487) );
  NOR2_X1 U541 ( .A1(n488), .A2(n487), .ZN(n501) );
  XOR2_X1 U542 ( .A(KEYINPUT83), .B(KEYINPUT16), .Z(n490) );
  OR2_X1 U543 ( .A1(n503), .A2(n570), .ZN(n489) );
  XNOR2_X1 U544 ( .A(n490), .B(n489), .ZN(n491) );
  OR2_X1 U545 ( .A1(n501), .A2(n491), .ZN(n516) );
  NOR2_X1 U546 ( .A1(n506), .A2(n516), .ZN(n498) );
  NAND2_X1 U547 ( .A1(n498), .A2(n529), .ZN(n492) );
  XNOR2_X1 U548 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n494), .ZN(G1324GAT) );
  NAND2_X1 U550 ( .A1(n498), .A2(n531), .ZN(n495) );
  XNOR2_X1 U551 ( .A(n495), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .Z(n497) );
  NAND2_X1 U553 ( .A1(n498), .A2(n544), .ZN(n496) );
  XNOR2_X1 U554 ( .A(n497), .B(n496), .ZN(G1326GAT) );
  INV_X1 U555 ( .A(n547), .ZN(n537) );
  NAND2_X1 U556 ( .A1(n498), .A2(n537), .ZN(n499) );
  XNOR2_X1 U557 ( .A(n499), .B(KEYINPUT104), .ZN(n500) );
  XNOR2_X1 U558 ( .A(G22GAT), .B(n500), .ZN(G1327GAT) );
  XOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT39), .Z(n509) );
  NOR2_X1 U560 ( .A1(n592), .A2(n501), .ZN(n502) );
  NAND2_X1 U561 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U562 ( .A(KEYINPUT37), .B(n504), .ZN(n505) );
  XNOR2_X1 U563 ( .A(KEYINPUT105), .B(n505), .ZN(n526) );
  NOR2_X1 U564 ( .A1(n506), .A2(n526), .ZN(n507) );
  XNOR2_X1 U565 ( .A(n507), .B(KEYINPUT38), .ZN(n513) );
  NAND2_X1 U566 ( .A1(n513), .A2(n529), .ZN(n508) );
  XNOR2_X1 U567 ( .A(n509), .B(n508), .ZN(G1328GAT) );
  NAND2_X1 U568 ( .A1(n513), .A2(n531), .ZN(n510) );
  XNOR2_X1 U569 ( .A(n510), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U570 ( .A1(n513), .A2(n544), .ZN(n511) );
  XNOR2_X1 U571 ( .A(n511), .B(KEYINPUT40), .ZN(n512) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n512), .ZN(G1330GAT) );
  XNOR2_X1 U573 ( .A(G50GAT), .B(KEYINPUT106), .ZN(n515) );
  NAND2_X1 U574 ( .A1(n537), .A2(n513), .ZN(n514) );
  XNOR2_X1 U575 ( .A(n515), .B(n514), .ZN(G1331GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n518) );
  INV_X1 U577 ( .A(n581), .ZN(n561) );
  NAND2_X1 U578 ( .A1(n561), .A2(n550), .ZN(n527) );
  NOR2_X1 U579 ( .A1(n527), .A2(n516), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n523), .A2(n529), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U582 ( .A(G57GAT), .B(n519), .ZN(G1332GAT) );
  NAND2_X1 U583 ( .A1(n523), .A2(n531), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U585 ( .A(G71GAT), .B(KEYINPUT109), .Z(n522) );
  NAND2_X1 U586 ( .A1(n523), .A2(n544), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(G1334GAT) );
  XOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT43), .Z(n525) );
  NAND2_X1 U589 ( .A1(n523), .A2(n537), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(KEYINPUT110), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n536), .A2(n529), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U595 ( .A(G92GAT), .B(KEYINPUT111), .Z(n533) );
  NAND2_X1 U596 ( .A1(n531), .A2(n536), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(G1337GAT) );
  NAND2_X1 U598 ( .A1(n536), .A2(n544), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n534), .B(KEYINPUT112), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G99GAT), .B(n535), .ZN(G1338GAT) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n541) );
  XOR2_X1 U602 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n539) );
  NAND2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1339GAT) );
  NOR2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n560) );
  NAND2_X1 U607 ( .A1(n560), .A2(n544), .ZN(n545) );
  XOR2_X1 U608 ( .A(KEYINPUT116), .B(n545), .Z(n546) );
  NAND2_X1 U609 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U610 ( .A(n548), .B(KEYINPUT117), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n556), .A2(n581), .ZN(n549) );
  XNOR2_X1 U612 ( .A(G113GAT), .B(n549), .ZN(G1340GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n552) );
  NAND2_X1 U614 ( .A1(n556), .A2(n550), .ZN(n551) );
  XNOR2_X1 U615 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U616 ( .A(G120GAT), .B(n553), .ZN(G1341GAT) );
  NAND2_X1 U617 ( .A1(n589), .A2(n556), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n554), .B(KEYINPUT50), .ZN(n555) );
  XNOR2_X1 U619 ( .A(G127GAT), .B(n555), .ZN(G1342GAT) );
  XOR2_X1 U620 ( .A(G134GAT), .B(KEYINPUT51), .Z(n558) );
  NAND2_X1 U621 ( .A1(n556), .A2(n570), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n558), .B(n557), .ZN(G1343GAT) );
  NAND2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n564) );
  NOR2_X1 U624 ( .A1(n561), .A2(n564), .ZN(n563) );
  XNOR2_X1 U625 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n563), .B(n562), .ZN(G1344GAT) );
  INV_X1 U627 ( .A(n564), .ZN(n571) );
  NAND2_X1 U628 ( .A1(n392), .A2(n571), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(KEYINPUT120), .ZN(n566) );
  XOR2_X1 U630 ( .A(n566), .B(KEYINPUT52), .Z(n568) );
  XNOR2_X1 U631 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n589), .A2(n571), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U636 ( .A(n572), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U637 ( .A1(n574), .A2(n581), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G169GAT), .B(n573), .ZN(G1348GAT) );
  NAND2_X1 U639 ( .A1(n589), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U644 ( .A(KEYINPUT59), .B(n578), .Z(n583) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n588) );
  NAND2_X1 U646 ( .A1(n588), .A2(n581), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  INV_X1 U648 ( .A(n588), .ZN(n591) );
  NOR2_X1 U649 ( .A1(n591), .A2(n388), .ZN(n587) );
  XOR2_X1 U650 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n585) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n584) );
  XNOR2_X1 U652 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n590), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n594) );
  XNOR2_X1 U657 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n594), .B(n593), .ZN(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

