//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AND2_X1   g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT66), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT67), .B(G244), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G77), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G116), .A2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT68), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n212), .B1(new_n219), .B2(new_n220), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT70), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT69), .B(G50), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n245), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G1), .A2(G13), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  AND3_X1   g0054(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n206), .A2(G20), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G50), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT65), .B(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G33), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n259), .A2(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(G20), .B2(new_n203), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n254), .A2(new_n253), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI221_X1 g0067(.A(new_n257), .B1(G50), .B2(new_n252), .C1(new_n265), .C2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT9), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G222), .A2(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G223), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n253), .B1(G33), .B2(G41), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n278), .B(new_n279), .C1(G77), .C2(new_n274), .ZN(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n281), .B1(new_n217), .B2(new_n282), .ZN(new_n283));
  OR2_X1    g0083(.A1(KEYINPUT73), .A2(G41), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT73), .A2(G41), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n283), .B(new_n206), .C1(new_n286), .C2(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n217), .A2(new_n282), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G226), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n280), .A2(new_n287), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G200), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n269), .B(new_n293), .C1(new_n294), .C2(new_n292), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n295), .A2(KEYINPUT10), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(KEYINPUT10), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n292), .A2(G179), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT74), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT74), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n292), .B2(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n300), .B(new_n268), .C1(new_n299), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n255), .ZN(new_n306));
  INV_X1    g0106(.A(new_n260), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n256), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n306), .A2(new_n308), .B1(new_n252), .B2(new_n307), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT80), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT79), .B1(new_n270), .B2(KEYINPUT3), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT79), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(new_n272), .A3(G33), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n311), .A2(new_n313), .A3(new_n271), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT7), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n258), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(G68), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n311), .A2(new_n313), .A3(new_n271), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n315), .B1(new_n318), .B2(new_n207), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n310), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT7), .B1(new_n314), .B2(G20), .ZN(new_n321));
  INV_X1    g0121(.A(G68), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n213), .A2(new_n215), .A3(new_n315), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n318), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(KEYINPUT80), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G58), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n327), .A2(new_n322), .ZN(new_n328));
  OAI21_X1  g0128(.A(G20), .B1(new_n328), .B2(new_n202), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n262), .A2(G159), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT16), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n267), .B1(new_n326), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n271), .A2(new_n273), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n315), .B1(new_n335), .B2(new_n258), .ZN(new_n336));
  AOI211_X1 g0136(.A(KEYINPUT7), .B(G20), .C1(new_n271), .C2(new_n273), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n336), .A2(new_n337), .A3(new_n322), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n332), .B1(new_n338), .B2(new_n331), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n309), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G200), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G87), .ZN(new_n342));
  OR2_X1    g0142(.A1(G223), .A2(G1698), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(G226), .B2(new_n276), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n342), .B1(new_n318), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n345), .A2(new_n279), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n288), .A2(G232), .A3(new_n289), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n287), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT81), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n348), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n345), .A2(new_n279), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT81), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n341), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n346), .A2(new_n348), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n294), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n340), .A2(KEYINPUT17), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT17), .B1(new_n340), .B2(new_n357), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n302), .B1(new_n350), .B2(new_n353), .ZN(new_n361));
  INV_X1    g0161(.A(G179), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n340), .A2(new_n364), .A3(KEYINPUT18), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT18), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n317), .A2(new_n310), .A3(new_n319), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT80), .B1(new_n321), .B2(new_n324), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n333), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(new_n339), .A3(new_n266), .ZN(new_n370));
  INV_X1    g0170(.A(new_n309), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n349), .B1(new_n346), .B2(new_n348), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT81), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(new_n302), .B1(new_n362), .B2(new_n355), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n366), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n365), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n360), .A2(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n262), .A2(G50), .B1(G20), .B2(new_n322), .ZN(new_n380));
  INV_X1    g0180(.A(G77), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n380), .B1(new_n259), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n266), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT11), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n384), .A2(KEYINPUT78), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(KEYINPUT78), .ZN(new_n386));
  OR3_X1    g0186(.A1(new_n252), .A2(KEYINPUT12), .A3(G68), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT12), .B1(new_n252), .B2(G68), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n322), .B1(new_n206), .B2(G20), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n387), .A2(new_n388), .B1(new_n255), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n385), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(G226), .A2(G1698), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n233), .B2(G1698), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n274), .A2(new_n393), .B1(G33), .B2(G97), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT77), .ZN(new_n395));
  OR3_X1    g0195(.A1(new_n394), .A2(new_n395), .A3(new_n288), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n395), .B1(new_n394), .B2(new_n288), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n290), .A2(G238), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n399), .A2(new_n287), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT13), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT13), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n398), .A2(new_n403), .A3(new_n400), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT14), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(G169), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n362), .B2(new_n405), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n406), .B1(new_n405), .B2(G169), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n391), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n402), .A2(new_n404), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G190), .ZN(new_n412));
  INV_X1    g0212(.A(new_n391), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n405), .A2(G200), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n274), .A2(G238), .A3(G1698), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n274), .A2(G232), .A3(new_n276), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n335), .A2(G107), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n279), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n290), .A2(new_n221), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n422), .A2(new_n287), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G200), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n256), .A2(G77), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT75), .B1(new_n306), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT75), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n255), .A2(new_n428), .A3(G77), .A4(new_n256), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n216), .A2(G77), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT15), .B(G87), .ZN(new_n432));
  OAI221_X1 g0232(.A(new_n431), .B1(new_n263), .B2(new_n260), .C1(new_n259), .C2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n252), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n433), .A2(new_n266), .B1(new_n381), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n425), .A2(KEYINPUT76), .A3(new_n430), .A4(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT76), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n341), .B1(new_n421), .B2(new_n423), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n433), .A2(new_n266), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(new_n381), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(new_n430), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n437), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n421), .A2(G190), .A3(new_n423), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n436), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n424), .A2(new_n302), .B1(new_n435), .B2(new_n430), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n421), .A2(new_n423), .A3(new_n362), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NOR4_X1   g0248(.A1(new_n305), .A2(new_n379), .A3(new_n416), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G87), .ZN(new_n451));
  NOR4_X1   g0251(.A1(new_n216), .A2(new_n335), .A3(KEYINPUT22), .A4(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n258), .A2(new_n271), .A3(new_n311), .A4(new_n313), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT22), .B1(new_n453), .B2(new_n451), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT88), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(KEYINPUT88), .B(KEYINPUT22), .C1(new_n453), .C2(new_n451), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n452), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n258), .A2(KEYINPUT23), .A3(G107), .ZN(new_n459));
  NAND2_X1  g0259(.A1(KEYINPUT23), .A2(G107), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(G20), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n458), .A2(KEYINPUT24), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT24), .ZN(new_n466));
  INV_X1    g0266(.A(new_n452), .ZN(new_n467));
  INV_X1    g0267(.A(new_n457), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n270), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n272), .A2(G33), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n471), .A2(G87), .A3(new_n258), .A4(new_n311), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT88), .B1(new_n472), .B2(KEYINPUT22), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n467), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n466), .B1(new_n474), .B2(new_n463), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n266), .B1(new_n465), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G107), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT25), .B1(new_n434), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n434), .A2(KEYINPUT25), .A3(new_n477), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n206), .A2(G33), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n252), .A2(new_n481), .A3(new_n253), .A4(new_n254), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n479), .A2(new_n480), .B1(G107), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G294), .ZN(new_n485));
  INV_X1    g0285(.A(G250), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n276), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(G257), .B2(new_n276), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n485), .B1(new_n318), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n288), .B1(new_n489), .B2(KEYINPUT89), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT89), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n491), .B(new_n485), .C1(new_n318), .C2(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT5), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n206), .B(G45), .C1(new_n494), .C2(G41), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  AND2_X1   g0296(.A1(KEYINPUT73), .A2(G41), .ZN(new_n497));
  NOR2_X1   g0297(.A1(KEYINPUT73), .A2(G41), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n496), .A2(new_n499), .A3(new_n283), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n495), .B1(new_n286), .B2(new_n494), .ZN(new_n501));
  INV_X1    g0301(.A(G264), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n501), .A2(new_n502), .A3(new_n279), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n493), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n341), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(G190), .B2(new_n505), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n476), .A2(new_n484), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n505), .A2(G179), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n503), .B1(new_n490), .B2(new_n492), .ZN(new_n510));
  AOI21_X1  g0310(.A(G169), .B1(new_n510), .B2(new_n500), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT24), .B1(new_n458), .B2(new_n464), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n474), .A2(new_n466), .A3(new_n463), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n267), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n484), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n213), .A2(new_n215), .A3(G33), .A4(G97), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT19), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n453), .B2(new_n322), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT83), .ZN(new_n523));
  NAND3_X1  g0323(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n213), .A2(new_n215), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(G97), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n451), .A2(new_n526), .A3(new_n477), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n523), .B1(new_n258), .B2(new_n524), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n266), .B1(new_n522), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n432), .A2(new_n434), .ZN(new_n532));
  OR2_X1    g0332(.A1(new_n482), .A2(new_n432), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT84), .ZN(new_n535));
  INV_X1    g0335(.A(G244), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G1698), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(G238), .B2(G1698), .ZN(new_n538));
  INV_X1    g0338(.A(G116), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n318), .A2(new_n538), .B1(new_n270), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n279), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n206), .A2(new_n281), .A3(G45), .ZN(new_n542));
  INV_X1    g0342(.A(G45), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n486), .B1(new_n543), .B2(G1), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n288), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G169), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n541), .A2(G179), .A3(new_n545), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT84), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n531), .A2(new_n550), .A3(new_n532), .A4(new_n533), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n535), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n531), .A2(new_n532), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n541), .A2(G190), .A3(new_n545), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n483), .A2(G87), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n546), .A2(G200), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT85), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n279), .B1(new_n496), .B2(new_n499), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(G270), .B1(new_n501), .B2(new_n283), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n335), .A2(G303), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n502), .A2(G1698), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(G257), .B2(G1698), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n562), .B1(new_n318), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n279), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n567), .A2(new_n362), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n254), .A2(new_n253), .B1(G20), .B2(new_n539), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n270), .A2(G97), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G283), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n569), .B(KEYINPUT20), .C1(new_n216), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT87), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n569), .B1(new_n216), .B2(new_n572), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT20), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n258), .A2(new_n571), .A3(new_n570), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT87), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT20), .A4(new_n569), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n574), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n252), .A2(G116), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT86), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n255), .A2(new_n583), .A3(G116), .A4(new_n481), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT86), .B1(new_n482), .B2(new_n539), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n568), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n581), .A2(new_n586), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n567), .A2(G200), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n561), .A2(G190), .A3(new_n566), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n302), .B1(new_n561), .B2(new_n566), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT21), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n587), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n594), .B1(new_n587), .B2(new_n593), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n588), .B(new_n592), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n336), .A2(new_n337), .A3(new_n477), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n262), .A2(G77), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n599), .B(KEYINPUT82), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT6), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n601), .A2(new_n526), .A3(G107), .ZN(new_n602));
  XNOR2_X1  g0402(.A(G97), .B(G107), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n602), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n600), .B1(new_n258), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n266), .B1(new_n598), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n252), .A2(G97), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n483), .B2(G97), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT5), .B1(new_n284), .B2(new_n285), .ZN(new_n610));
  OAI211_X1 g0410(.A(G257), .B(new_n288), .C1(new_n610), .C2(new_n495), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n500), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n271), .A2(new_n273), .A3(G250), .A4(G1698), .ZN(new_n613));
  AND2_X1   g0413(.A1(KEYINPUT4), .A2(G244), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n271), .A2(new_n273), .A3(new_n614), .A4(new_n276), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n613), .A2(new_n615), .A3(new_n571), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT4), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n276), .A2(G244), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(new_n318), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n612), .B1(new_n620), .B2(new_n279), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n362), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n288), .B1(new_n616), .B2(new_n619), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n302), .B1(new_n623), .B2(new_n612), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n609), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n608), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n603), .A2(new_n601), .ZN(new_n627));
  INV_X1    g0427(.A(new_n602), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n258), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT82), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n599), .B(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT7), .B1(new_n274), .B2(new_n216), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n335), .A2(new_n315), .A3(new_n207), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G107), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n626), .B1(new_n636), .B2(new_n266), .ZN(new_n637));
  INV_X1    g0437(.A(new_n623), .ZN(new_n638));
  INV_X1    g0438(.A(new_n612), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(G190), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(G200), .B1(new_n623), .B2(new_n612), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n625), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n597), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT85), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n552), .A2(new_n645), .A3(new_n557), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n559), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n450), .A2(new_n518), .A3(new_n647), .ZN(G372));
  NAND2_X1  g0448(.A1(new_n549), .A2(new_n534), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n557), .A2(new_n625), .A3(new_n642), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n508), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n588), .B1(new_n595), .B2(new_n596), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n517), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n650), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n557), .A2(new_n649), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n658), .A2(KEYINPUT26), .A3(new_n625), .ZN(new_n659));
  INV_X1    g0459(.A(new_n625), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n559), .A2(new_n646), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n659), .B1(new_n661), .B2(KEYINPUT26), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n449), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g0464(.A(new_n664), .B(KEYINPUT90), .Z(new_n665));
  INV_X1    g0465(.A(new_n304), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n410), .A2(new_n447), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n360), .A2(new_n415), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n378), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n666), .B1(new_n669), .B2(new_n298), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n665), .A2(new_n670), .ZN(G369));
  NAND3_X1  g0471(.A1(new_n258), .A2(new_n206), .A3(G13), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n476), .B2(new_n484), .ZN(new_n679));
  OAI22_X1  g0479(.A1(new_n518), .A2(new_n679), .B1(new_n517), .B2(new_n678), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n678), .A2(new_n589), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n654), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n597), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n476), .A2(new_n484), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(new_n512), .A3(new_n678), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n508), .A2(new_n517), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n655), .A2(new_n677), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n686), .A2(new_n688), .A3(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n286), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n210), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n527), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n220), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(new_n545), .ZN(new_n699));
  AOI211_X1 g0499(.A(new_n362), .B(new_n699), .C1(new_n540), .C2(new_n279), .ZN(new_n700));
  NOR2_X1   g0500(.A1(G257), .A2(G1698), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n502), .B2(G1698), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n471), .A2(new_n311), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n288), .B1(new_n703), .B2(new_n562), .ZN(new_n704));
  OAI211_X1 g0504(.A(G270), .B(new_n288), .C1(new_n610), .C2(new_n495), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n500), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n510), .A2(new_n621), .A3(new_n700), .A4(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n567), .A2(new_n548), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(KEYINPUT30), .A3(new_n510), .A4(new_n621), .ZN(new_n712));
  INV_X1    g0512(.A(new_n621), .ZN(new_n713));
  AOI21_X1  g0513(.A(G179), .B1(new_n541), .B2(new_n545), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n505), .A2(new_n713), .A3(new_n567), .A4(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n710), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT31), .B1(new_n716), .B2(new_n677), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT91), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT91), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n716), .A2(new_n677), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(KEYINPUT31), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n647), .A2(new_n518), .A3(new_n677), .ZN(new_n724));
  OAI21_X1  g0524(.A(G330), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT92), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT92), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n727), .B(G330), .C1(new_n723), .C2(new_n724), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n677), .B1(new_n657), .B2(new_n662), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT26), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n658), .A2(new_n733), .A3(new_n625), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n661), .B2(new_n733), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n654), .B1(new_n687), .B2(new_n512), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n649), .B1(new_n736), .B2(new_n652), .ZN(new_n737));
  OAI211_X1 g0537(.A(KEYINPUT29), .B(new_n678), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n730), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n698), .B1(new_n741), .B2(G1), .ZN(G364));
  AND2_X1   g0542(.A1(new_n258), .A2(G13), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G45), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(new_n694), .A3(G1), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n210), .A2(new_n274), .ZN(new_n747));
  INV_X1    g0547(.A(G355), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n747), .A2(new_n748), .B1(G116), .B2(new_n210), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n245), .A2(G45), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n210), .A2(new_n318), .ZN(new_n751));
  INV_X1    g0551(.A(new_n220), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n751), .B1(new_n543), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n749), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n217), .B1(new_n207), .B2(G169), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n755), .A2(KEYINPUT93), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(KEYINPUT93), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G13), .A2(G33), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n746), .B1(new_n754), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n758), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n341), .A2(G179), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(G20), .A3(G190), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n274), .B1(new_n767), .B2(new_n451), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G190), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n216), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n526), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n258), .A2(G190), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n766), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n768), .B(new_n773), .C1(G107), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n362), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n216), .A2(G190), .A3(new_n778), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n779), .A2(new_n381), .B1(new_n327), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n362), .A2(new_n341), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n774), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G50), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n216), .A2(G190), .A3(new_n782), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n783), .A2(new_n322), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n774), .A2(new_n769), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n790));
  OR3_X1    g0590(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n790), .B1(new_n788), .B2(new_n789), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n777), .A2(new_n787), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n767), .B(KEYINPUT95), .Z(new_n794));
  AOI22_X1  g0594(.A1(new_n794), .A2(G303), .B1(new_n776), .B2(G283), .ZN(new_n795));
  INV_X1    g0595(.A(G294), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n335), .B1(new_n772), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n780), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(G322), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n779), .ZN(new_n800));
  INV_X1    g0600(.A(new_n788), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G311), .A2(new_n800), .B1(new_n801), .B2(G329), .ZN(new_n802));
  INV_X1    g0602(.A(new_n783), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT33), .B(G317), .ZN(new_n804));
  INV_X1    g0604(.A(new_n785), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n803), .A2(new_n804), .B1(G326), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n795), .A2(new_n799), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n765), .B1(new_n793), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n764), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n761), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n683), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n684), .A2(new_n745), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n683), .A2(G330), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(G396));
  NAND2_X1  g0614(.A1(new_n441), .A2(new_n677), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n444), .A2(new_n447), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n424), .A2(new_n302), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n817), .A2(new_n441), .A3(new_n446), .A4(new_n677), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT97), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n445), .A2(KEYINPUT97), .A3(new_n446), .A4(new_n677), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n816), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(KEYINPUT98), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT98), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n816), .A2(new_n825), .A3(new_n822), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n731), .B(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(KEYINPUT99), .B1(new_n829), .B2(new_n729), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n746), .B1(new_n829), .B2(new_n729), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n829), .A2(new_n729), .A3(KEYINPUT99), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n765), .A2(new_n760), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT96), .Z(new_n836));
  OAI21_X1  g0636(.A(new_n746), .B1(new_n836), .B2(G77), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n274), .B(new_n773), .C1(G283), .C2(new_n803), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G116), .A2(new_n800), .B1(new_n801), .B2(G311), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n794), .A2(G107), .B1(new_n776), .B2(G87), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G294), .A2(new_n798), .B1(new_n805), .B2(G303), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n314), .B1(new_n772), .B2(new_n327), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G132), .B2(new_n801), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n794), .A2(G50), .B1(new_n776), .B2(G68), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G137), .A2(new_n805), .B1(new_n798), .B2(G143), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n846), .B1(new_n261), .B2(new_n783), .C1(new_n789), .C2(new_n779), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT34), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n844), .B(new_n845), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n842), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n837), .B1(new_n851), .B2(new_n758), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n827), .B2(new_n760), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n834), .A2(new_n853), .ZN(G384));
  XOR2_X1   g0654(.A(new_n604), .B(KEYINPUT35), .Z(new_n855));
  NOR3_X1   g0655(.A1(new_n855), .A2(new_n539), .A3(new_n219), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT36), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n201), .A2(G68), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n752), .B(G77), .C1(new_n327), .C2(new_n322), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n206), .B(G13), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n675), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n378), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n369), .A2(new_n266), .ZN(new_n864));
  INV_X1    g0664(.A(new_n331), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT16), .B1(new_n326), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n371), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT100), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n331), .B1(new_n320), .B2(new_n325), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n369), .B(new_n266), .C1(new_n870), .C2(KEYINPUT16), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(KEYINPUT100), .A3(new_n371), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n869), .A2(new_n862), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n360), .B2(new_n378), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n364), .A2(new_n675), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n869), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n340), .A2(new_n357), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT101), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n372), .A2(new_n376), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n372), .A2(new_n862), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n883), .A3(new_n878), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n877), .B2(new_n878), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n889), .A2(new_n880), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n875), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(KEYINPUT38), .B(new_n875), .C1(new_n887), .C2(new_n890), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n447), .A2(new_n677), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n731), .B2(new_n827), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT14), .B1(new_n411), .B2(new_n302), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n898), .B(new_n407), .C1(new_n362), .C2(new_n405), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n391), .B(new_n677), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n391), .A2(new_n677), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n410), .A2(new_n415), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n897), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n863), .B1(new_n895), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n899), .A2(new_n391), .A3(new_n678), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n885), .B1(new_n889), .B2(new_n880), .ZN(new_n910));
  INV_X1    g0710(.A(new_n878), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n865), .B1(new_n367), .B2(new_n368), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n332), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n868), .B(new_n309), .C1(new_n913), .C2(new_n334), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT100), .B1(new_n871), .B2(new_n371), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n911), .B1(new_n916), .B2(new_n876), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT101), .B1(new_n917), .B2(new_n888), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n874), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n919), .A2(KEYINPUT38), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n892), .B(new_n874), .C1(new_n910), .C2(new_n918), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT39), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n379), .A2(new_n372), .A3(new_n862), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n884), .B(KEYINPUT37), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT38), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n919), .B2(KEYINPUT38), .ZN(new_n926));
  XOR2_X1   g0726(.A(KEYINPUT102), .B(KEYINPUT39), .Z(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n909), .B1(new_n922), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n908), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n449), .A2(new_n732), .A3(new_n738), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n670), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n930), .B(new_n932), .Z(new_n933));
  INV_X1    g0733(.A(KEYINPUT40), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n923), .A2(new_n924), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n892), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n894), .A2(new_n936), .ZN(new_n937));
  OR3_X1    g0737(.A1(new_n647), .A2(new_n518), .A3(new_n677), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n717), .A2(new_n718), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n904), .A2(new_n827), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n934), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n904), .A2(new_n940), .A3(new_n934), .A4(new_n827), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n893), .B2(new_n894), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n449), .A2(new_n940), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(G330), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n933), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n206), .B2(new_n743), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n933), .A2(new_n949), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n861), .B1(new_n951), .B2(new_n952), .ZN(G367));
  NAND2_X1  g0753(.A1(new_n744), .A2(G1), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n691), .A2(new_n688), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n660), .A2(new_n677), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n625), .B(new_n642), .C1(new_n637), .C2(new_n678), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT44), .Z(new_n962));
  NOR2_X1   g0762(.A1(new_n956), .A2(new_n960), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT45), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT104), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n686), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n680), .A2(new_n690), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n969), .A2(new_n691), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n685), .A2(KEYINPUT105), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n685), .A2(KEYINPUT105), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n972), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n740), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n686), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n965), .A2(new_n966), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n968), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT106), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT106), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n968), .A2(new_n981), .A3(new_n976), .A4(new_n978), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n740), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n694), .B(KEYINPUT41), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n955), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n678), .B1(new_n553), .B2(new_n555), .ZN(new_n986));
  MUX2_X1   g0786(.A(new_n658), .B(new_n649), .S(new_n986), .Z(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT103), .Z(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n689), .A2(new_n690), .A3(new_n959), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n990), .A2(KEYINPUT42), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n625), .B1(new_n517), .B2(new_n958), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n990), .A2(KEYINPUT42), .B1(new_n678), .B2(new_n992), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n989), .A2(KEYINPUT43), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n977), .A2(new_n959), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n985), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n762), .B1(new_n210), .B2(new_n432), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n239), .A2(new_n751), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n746), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n274), .B1(new_n767), .B2(new_n327), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n201), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G159), .A2(new_n803), .B1(new_n800), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n381), .B2(new_n775), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(KEYINPUT109), .B(G137), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1003), .B(new_n1006), .C1(new_n801), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT108), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n771), .A2(G68), .ZN(new_n1010));
  INV_X1    g0810(.A(G143), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1010), .B1(new_n780), .B2(new_n261), .C1(new_n1011), .C2(new_n785), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1008), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT110), .Z(new_n1015));
  INV_X1    g0815(.A(G317), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n318), .B1(new_n788), .B2(new_n1016), .C1(new_n526), .C2(new_n775), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1017), .A2(KEYINPUT107), .ZN(new_n1018));
  INV_X1    g0818(.A(G283), .ZN(new_n1019));
  INV_X1    g0819(.A(G303), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n779), .A2(new_n1019), .B1(new_n1020), .B2(new_n780), .ZN(new_n1021));
  AND3_X1   g0821(.A1(new_n794), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(G311), .C2(new_n805), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1017), .A2(KEYINPUT107), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n767), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT46), .B1(new_n1025), .B2(G116), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n772), .A2(new_n477), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(G294), .C2(new_n803), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1023), .A2(new_n1024), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1015), .B1(new_n1018), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(KEYINPUT47), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n765), .B1(new_n1031), .B2(KEYINPUT47), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1002), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n988), .A2(new_n761), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n999), .A2(new_n1036), .ZN(G387));
  INV_X1    g0837(.A(new_n975), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n680), .A2(new_n810), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n747), .A2(new_n695), .B1(G107), .B2(new_n210), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n236), .A2(new_n543), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n695), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n1042), .C1(G68), .C2(G77), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n260), .A2(G50), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT50), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n751), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1040), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n746), .B1(new_n1047), .B2(new_n763), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n772), .A2(new_n432), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n318), .B(new_n1049), .C1(G77), .C2(new_n1025), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G68), .A2(new_n800), .B1(new_n803), .B2(new_n307), .ZN(new_n1051));
  XOR2_X1   g0851(.A(KEYINPUT111), .B(G150), .Z(new_n1052));
  AOI22_X1  g0852(.A1(new_n801), .A2(new_n1052), .B1(G159), .B2(new_n805), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n776), .A2(G97), .B1(G50), .B2(new_n798), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n772), .A2(new_n1019), .B1(new_n796), .B2(new_n767), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(KEYINPUT112), .B(G322), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n800), .A2(G303), .B1(new_n805), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(G311), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1058), .B1(new_n1059), .B2(new_n783), .C1(new_n1016), .C2(new_n780), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1056), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n1061), .B2(new_n1060), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT49), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n314), .B1(new_n801), .B2(G326), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n539), .B2(new_n775), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT113), .Z(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1055), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1048), .B1(new_n1070), .B2(new_n758), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1038), .A2(new_n954), .B1(new_n1039), .B2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n741), .A2(new_n1038), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n694), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n740), .B2(new_n975), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1072), .B1(new_n1073), .B2(new_n1075), .ZN(G393));
  XNOR2_X1  g0876(.A(new_n965), .B(new_n686), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n954), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n250), .A2(new_n210), .A3(new_n318), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n762), .B1(new_n526), .B2(new_n210), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n314), .B1(new_n322), .B2(new_n767), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G87), .A2(new_n776), .B1(new_n800), .B2(new_n307), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n1011), .B2(new_n788), .C1(new_n201), .C2(new_n783), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1081), .B(new_n1083), .C1(G77), .C2(new_n771), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n261), .A2(new_n785), .B1(new_n780), .B2(new_n789), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT51), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1059), .A2(new_n780), .B1(new_n785), .B2(new_n1016), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT52), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n801), .A2(new_n1057), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1019), .B2(new_n767), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1090), .A2(KEYINPUT114), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1090), .A2(KEYINPUT114), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n335), .B1(new_n772), .B2(new_n539), .C1(new_n775), .C2(new_n477), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n796), .A2(new_n779), .B1(new_n783), .B2(new_n1020), .ZN(new_n1094));
  NOR4_X1   g0894(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1084), .A2(new_n1086), .B1(new_n1088), .B2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n746), .B1(new_n1079), .B2(new_n1080), .C1(new_n1096), .C2(new_n765), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT115), .Z(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n810), .B2(new_n959), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1078), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n980), .A2(new_n982), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1077), .A2(new_n976), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1102), .A2(new_n694), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1100), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(G390));
  INV_X1    g0905(.A(G330), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n938), .B2(new_n939), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n449), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n931), .A2(new_n670), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1107), .A2(new_n827), .A3(new_n904), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n828), .B1(new_n726), .B2(new_n728), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1110), .B1(new_n1111), .B2(new_n904), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n659), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n552), .A2(new_n645), .A3(new_n557), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n645), .B1(new_n552), .B2(new_n557), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n1114), .A2(new_n1115), .A3(new_n625), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1113), .B1(new_n1116), .B2(new_n733), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n827), .B(new_n678), .C1(new_n1117), .C2(new_n737), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n896), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1112), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n904), .B1(new_n1107), .B2(new_n827), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n827), .B(new_n678), .C1(new_n735), .C2(new_n737), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1119), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT116), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1123), .A2(KEYINPUT116), .A3(new_n1119), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1122), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n729), .A2(new_n827), .A3(new_n904), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1109), .B1(new_n1121), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1110), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT39), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n893), .B2(new_n894), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n894), .A2(new_n936), .A3(new_n927), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n909), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n1120), .B2(new_n904), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n909), .B1(new_n921), .B2(new_n925), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1123), .A2(KEYINPUT116), .A3(new_n1119), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT116), .B1(new_n1123), .B2(new_n1119), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1139), .B1(new_n1142), .B2(new_n904), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1132), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n909), .B1(new_n897), .B2(new_n905), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n922), .A2(new_n928), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1126), .A2(new_n904), .A3(new_n1127), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1136), .B1(new_n894), .B2(new_n936), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1146), .A2(new_n1149), .A3(new_n1129), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1131), .A2(new_n1144), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT117), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1131), .A2(new_n1144), .A3(KEYINPUT117), .A4(new_n1150), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1144), .A2(new_n1150), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1131), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n694), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1156), .A2(new_n955), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n794), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n1161), .A2(new_n451), .B1(new_n539), .B2(new_n780), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n526), .A2(new_n779), .B1(new_n788), .B2(new_n796), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n335), .B1(new_n772), .B2(new_n381), .C1(new_n775), .C2(new_n322), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n783), .A2(new_n477), .B1(new_n1019), .B2(new_n785), .ZN(new_n1165));
  NOR4_X1   g0965(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT120), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n805), .A2(G128), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1025), .A2(new_n1052), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT119), .ZN(new_n1170));
  XOR2_X1   g0970(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1171));
  XNOR2_X1  g0971(.A(new_n1170), .B(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1004), .A2(new_n776), .B1(new_n803), .B2(new_n1007), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n274), .B1(new_n772), .B2(new_n789), .ZN(new_n1174));
  INV_X1    g0974(.A(G125), .ZN(new_n1175));
  INV_X1    g0975(.A(G132), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n788), .A2(new_n1175), .B1(new_n1176), .B2(new_n780), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT54), .B(G143), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1174), .B(new_n1177), .C1(new_n800), .C2(new_n1179), .ZN(new_n1180));
  AND4_X1   g0980(.A1(new_n1168), .A2(new_n1172), .A3(new_n1173), .A4(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1167), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1182), .A2(new_n765), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n746), .B1(new_n836), .B2(new_n307), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1183), .B(new_n1184), .C1(new_n1185), .C2(new_n759), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1160), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1159), .A2(new_n1187), .ZN(G378));
  OAI21_X1  g0988(.A(new_n746), .B1(new_n835), .B2(new_n1004), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n772), .A2(new_n261), .B1(new_n767), .B2(new_n1178), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n800), .A2(G137), .B1(G128), .B2(new_n798), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n1175), .B2(new_n785), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(G132), .C2(new_n803), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n776), .A2(G159), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G33), .B(G41), .C1(new_n801), .C2(G124), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n776), .A2(G58), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT121), .Z(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n526), .A2(new_n783), .B1(new_n779), .B2(new_n432), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT122), .Z(new_n1204));
  OAI221_X1 g1004(.A(new_n1010), .B1(new_n381), .B2(new_n767), .C1(new_n539), .C2(new_n785), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n314), .A2(new_n286), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n477), .B2(new_n780), .C1(new_n788), .C2(new_n1019), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .A4(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1198), .A2(new_n1199), .B1(new_n1208), .B2(KEYINPUT58), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n784), .B1(G33), .B2(G41), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1209), .B1(KEYINPUT58), .B2(new_n1208), .C1(new_n1206), .C2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1189), .B1(new_n1211), .B2(new_n758), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n268), .A2(new_n862), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT123), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n305), .B(new_n1214), .ZN(new_n1215));
  XOR2_X1   g1015(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1216));
  XOR2_X1   g1016(.A(new_n1215), .B(new_n1216), .Z(new_n1217));
  OAI21_X1  g1017(.A(new_n1212), .B1(new_n1217), .B2(new_n760), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n904), .A2(new_n940), .A3(new_n827), .ZN(new_n1219));
  OAI21_X1  g1019(.A(KEYINPUT40), .B1(new_n926), .B2(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n934), .B(new_n941), .C1(new_n920), .C2(new_n921), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1106), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n908), .B2(new_n929), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1136), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1224), .B(new_n907), .C1(new_n945), .C2(new_n1106), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1217), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1223), .A2(new_n1225), .A3(new_n1217), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1218), .B1(new_n1230), .B2(new_n955), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1109), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1146), .A2(new_n1149), .A3(new_n1129), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1110), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT117), .B1(new_n1236), .B2(new_n1131), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1154), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1233), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1109), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1228), .A2(KEYINPUT57), .A3(new_n1229), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1074), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1232), .B1(new_n1241), .B2(new_n1244), .ZN(G375));
  NAND2_X1  g1045(.A1(new_n905), .A2(new_n759), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n746), .B1(new_n836), .B2(G68), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n1161), .A2(new_n526), .B1(new_n1020), .B2(new_n788), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n779), .A2(new_n477), .B1(new_n1019), .B2(new_n780), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n335), .B1(new_n772), .B2(new_n432), .C1(new_n775), .C2(new_n381), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n783), .A2(new_n539), .B1(new_n796), .B2(new_n785), .ZN(new_n1251));
  NOR4_X1   g1051(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n794), .A2(G159), .B1(new_n798), .B2(new_n1007), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1176), .B2(new_n785), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n314), .B1(new_n772), .B2(new_n784), .C1(new_n783), .C2(new_n1178), .ZN(new_n1255));
  INV_X1    g1055(.A(G128), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n1256), .A2(new_n788), .B1(new_n779), .B2(new_n261), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1252), .B1(new_n1258), .B2(new_n1201), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT124), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n765), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1247), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1246), .A2(new_n1263), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1112), .A2(new_n1120), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1264), .B1(new_n1265), .B2(new_n955), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1131), .A2(new_n984), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1109), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1267), .B1(new_n1268), .B2(new_n1270), .ZN(G381));
  OR2_X1    g1071(.A1(G393), .A2(G396), .ZN(new_n1272));
  OR4_X1    g1072(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1272), .ZN(new_n1273));
  OR4_X1    g1073(.A1(G387), .A2(new_n1273), .A3(G378), .A4(G375), .ZN(G407));
  AOI211_X1 g1074(.A(new_n1160), .B(new_n1186), .C1(new_n1155), .C2(new_n1158), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n676), .A2(G213), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G407), .B(G213), .C1(G375), .C2(new_n1278), .ZN(G409));
  NAND2_X1  g1079(.A1(new_n1277), .A2(G2897), .ZN(new_n1280));
  INV_X1    g1080(.A(G384), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1121), .A2(KEYINPUT60), .A3(new_n1109), .A4(new_n1130), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1074), .ZN(new_n1283));
  OAI21_X1  g1083(.A(KEYINPUT60), .B1(new_n1265), .B2(new_n1109), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1283), .B1(new_n1269), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1281), .B1(new_n1285), .B2(new_n1266), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1284), .A2(new_n1269), .ZN(new_n1287));
  OAI211_X1 g1087(.A(G384), .B(new_n1267), .C1(new_n1287), .C2(new_n1283), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1286), .A2(new_n1288), .A3(KEYINPUT125), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT125), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1280), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1288), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1286), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G2897), .B(new_n1277), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1291), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT126), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  OAI211_X1 g1097(.A(G378), .B(new_n1232), .C1(new_n1241), .C2(new_n1244), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1242), .A2(new_n984), .A3(new_n1230), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1275), .B1(new_n1299), .B2(new_n1231), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1277), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1291), .A2(KEYINPUT126), .A3(new_n1294), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1297), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  OR2_X1    g1104(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1301), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT127), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(new_n999), .B2(new_n1036), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1036), .ZN(new_n1312));
  AOI211_X1 g1112(.A(KEYINPUT127), .B(new_n1312), .C1(new_n985), .C2(new_n998), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(G393), .B(G396), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1104), .B(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1311), .A2(new_n1314), .A3(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1316), .B1(new_n1310), .B2(new_n1313), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT61), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1301), .A2(KEYINPUT63), .A3(new_n1305), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1304), .A2(new_n1308), .A3(new_n1320), .A4(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT62), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1301), .A2(new_n1323), .A3(new_n1305), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT61), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1325), .B1(new_n1301), .B2(new_n1295), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1323), .B1(new_n1301), .B2(new_n1305), .ZN(new_n1327));
  NOR3_X1   g1127(.A1(new_n1324), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1322), .B1(new_n1328), .B2(new_n1329), .ZN(G405));
  NAND2_X1  g1130(.A1(G375), .A2(new_n1275), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1298), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1305), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1331), .B(new_n1298), .C1(new_n1293), .C2(new_n1292), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1329), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1335), .B(new_n1336), .ZN(G402));
endmodule


