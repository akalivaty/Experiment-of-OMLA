//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1209, new_n1210, new_n1211, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1267, new_n1268;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT65), .Z(G353));
  OAI21_X1  g0010(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT66), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g0018(.A1(KEYINPUT66), .A2(G1), .A3(G13), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n206), .A2(new_n207), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(KEYINPUT67), .B(G238), .Z(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n203), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G107), .A2(G264), .ZN(new_n231));
  NAND4_X1  g0031(.A1(new_n228), .A2(new_n229), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n212), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n215), .B(new_n225), .C1(KEYINPUT1), .C2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G351));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G274), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n254), .A2(new_n257), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n258), .B1(G226), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n220), .A2(new_n253), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G222), .A2(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G223), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G77), .B2(new_n263), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n261), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G179), .ZN(new_n270));
  INV_X1    g0070(.A(G169), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(new_n269), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n208), .A2(G20), .ZN(new_n273));
  INV_X1    g0073(.A(G150), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n277), .B(KEYINPUT69), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n222), .A2(G33), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n273), .B1(new_n274), .B2(new_n276), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n218), .B(new_n219), .C1(new_n281), .C2(new_n212), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G13), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n284), .A2(new_n222), .A3(G1), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n222), .A2(G1), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n207), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n286), .A2(new_n288), .B1(new_n207), .B2(new_n285), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n272), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g0091(.A(KEYINPUT75), .B(KEYINPUT12), .Z(new_n292));
  NOR2_X1   g0092(.A1(new_n284), .A2(G1), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT70), .B1(new_n294), .B2(new_n222), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT70), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n285), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n292), .B1(new_n298), .B2(G68), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT76), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n203), .A2(G20), .ZN(new_n301));
  OR3_X1    g0101(.A1(new_n294), .A2(KEYINPUT12), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G77), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n301), .B1(new_n279), .B2(new_n304), .C1(new_n276), .C2(new_n207), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n282), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT11), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n282), .B1(new_n295), .B2(new_n297), .ZN(new_n308));
  INV_X1    g0108(.A(new_n287), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(G68), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n303), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G238), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n312), .A2(new_n259), .B1(new_n255), .B2(new_n257), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G97), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT73), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n314), .B(new_n315), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n265), .A2(G232), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(G226), .B2(G1698), .ZN(new_n318));
  INV_X1    g0118(.A(new_n263), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n262), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n313), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT13), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(new_n322), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G179), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n322), .B(new_n325), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT14), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(G169), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n329), .B1(new_n328), .B2(G169), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n311), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n326), .A2(G190), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n307), .A2(new_n310), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n328), .A2(G200), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n334), .A2(new_n303), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n263), .A2(G232), .A3(new_n265), .ZN(new_n339));
  INV_X1    g0139(.A(G107), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n263), .A2(G1698), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n339), .B1(new_n340), .B2(new_n263), .C1(new_n341), .C2(new_n226), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n321), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n258), .B1(G244), .B2(new_n260), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n271), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n277), .A2(new_n276), .B1(new_n222), .B2(new_n304), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT15), .B(G87), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(new_n279), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n282), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n308), .A2(G77), .A3(new_n309), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n350), .B(new_n351), .C1(G77), .C2(new_n298), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n343), .A2(new_n344), .ZN(new_n355));
  INV_X1    g0155(.A(G179), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT71), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n345), .A2(G179), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(KEYINPUT71), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n354), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n352), .B1(G200), .B2(new_n345), .ZN(new_n363));
  INV_X1    g0163(.A(G190), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(new_n364), .B2(new_n345), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n338), .B1(KEYINPUT72), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n269), .A2(new_n364), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(G200), .B2(new_n269), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n290), .A2(KEYINPUT9), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n290), .A2(KEYINPUT9), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT10), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n366), .A2(KEYINPUT72), .ZN(new_n374));
  AND4_X1   g0174(.A1(new_n291), .A2(new_n367), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n282), .ZN(new_n376));
  INV_X1    g0176(.A(G159), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n377), .A2(G20), .A3(G33), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G58), .A2(G68), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n204), .A2(new_n205), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n378), .B1(new_n380), .B2(G20), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT3), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(G33), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n222), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT79), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n383), .B2(G33), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n383), .A2(G33), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n281), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n382), .A2(G20), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n382), .A2(new_n386), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n381), .B1(new_n393), .B2(new_n203), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n376), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT78), .ZN(new_n397));
  AOI211_X1 g0197(.A(new_n395), .B(new_n378), .C1(new_n380), .C2(G20), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n383), .A2(KEYINPUT77), .A3(G33), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n263), .B2(KEYINPUT77), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n382), .B1(new_n400), .B2(new_n222), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(new_n389), .A3(KEYINPUT77), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT77), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(new_n281), .A3(KEYINPUT3), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n403), .A2(new_n382), .A3(new_n222), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G68), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n397), .B(new_n398), .C1(new_n401), .C2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n403), .A2(new_n222), .A3(new_n405), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT7), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n411), .A2(G68), .A3(new_n406), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n397), .B1(new_n412), .B2(new_n398), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n396), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT80), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT80), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n396), .B(new_n416), .C1(new_n409), .C2(new_n413), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n278), .A2(new_n287), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n286), .B1(new_n285), .B2(new_n278), .ZN(new_n420));
  INV_X1    g0220(.A(G200), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n403), .A2(new_n405), .ZN(new_n422));
  MUX2_X1   g0222(.A(G223), .B(G226), .S(G1698), .Z(new_n423));
  AOI22_X1  g0223(.A1(new_n422), .A2(new_n423), .B1(G33), .B2(G87), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n424), .A2(new_n262), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n258), .B1(G232), .B2(new_n260), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n421), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n425), .A2(new_n426), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n427), .B1(G190), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n418), .A2(new_n420), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT82), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n420), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n415), .B2(new_n417), .ZN(new_n435));
  NAND2_X1  g0235(.A1(KEYINPUT82), .A2(KEYINPUT17), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(new_n432), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n429), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n417), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n398), .B1(new_n401), .B2(new_n407), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT78), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n408), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n416), .B1(new_n443), .B2(new_n396), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n420), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n271), .B1(new_n425), .B2(new_n426), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(G179), .B2(new_n428), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT18), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n445), .A2(KEYINPUT18), .A3(new_n448), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n449), .B1(KEYINPUT81), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n447), .B1(new_n418), .B2(new_n420), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT81), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT18), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n439), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n375), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  OR2_X1    g0257(.A1(G257), .A2(G1698), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(G264), .B2(new_n265), .ZN(new_n459));
  INV_X1    g0259(.A(G303), .ZN(new_n460));
  OAI22_X1  g0260(.A1(new_n400), .A2(new_n459), .B1(new_n460), .B2(new_n263), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT87), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT87), .ZN(new_n463));
  OAI221_X1 g0263(.A(new_n463), .B1(new_n460), .B2(new_n263), .C1(new_n400), .C2(new_n459), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n464), .A3(new_n321), .ZN(new_n465));
  NOR2_X1   g0265(.A1(KEYINPUT84), .A2(G41), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT5), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(KEYINPUT84), .B2(G41), .ZN(new_n469));
  INV_X1    g0269(.A(G45), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G1), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n467), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n255), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT85), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n467), .A2(new_n469), .A3(new_n471), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT85), .B1(new_n476), .B2(new_n255), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n476), .A2(new_n254), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G270), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n465), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G200), .ZN(new_n483));
  INV_X1    g0283(.A(new_n298), .ZN(new_n484));
  INV_X1    g0284(.A(G116), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n281), .A2(G1), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(new_n485), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n484), .A2(new_n485), .B1(new_n308), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(G20), .B1(G33), .B2(G283), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n281), .A2(G97), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n489), .A2(new_n490), .B1(G20), .B2(new_n485), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n282), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT20), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n492), .B(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n465), .A2(new_n481), .A3(G190), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n483), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n478), .A2(G179), .A3(new_n480), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n465), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n271), .B1(new_n488), .B2(new_n494), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT21), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n501), .A2(new_n482), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n501), .B2(new_n482), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n498), .B(new_n500), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n263), .A2(KEYINPUT4), .A3(G244), .A4(new_n265), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  INV_X1    g0308(.A(G250), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n507), .B(new_n508), .C1(new_n509), .C2(new_n341), .ZN(new_n510));
  INV_X1    g0310(.A(G244), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(G1698), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT4), .B1(new_n422), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n321), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n475), .A2(new_n477), .B1(new_n479), .B2(G257), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT86), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT86), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n517), .A2(G190), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n516), .A2(G200), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n393), .A2(new_n340), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n275), .A2(G77), .ZN(new_n523));
  XNOR2_X1  g0323(.A(new_n523), .B(KEYINPUT83), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT6), .ZN(new_n525));
  INV_X1    g0325(.A(G97), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n525), .A2(new_n526), .A3(G107), .ZN(new_n527));
  XNOR2_X1  g0327(.A(G97), .B(G107), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n527), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n524), .B1(new_n222), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n282), .B1(new_n522), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n285), .A2(new_n526), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n282), .A2(new_n285), .A3(new_n486), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G97), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n521), .A2(new_n531), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(G169), .B1(new_n517), .B2(new_n519), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n514), .A2(new_n515), .A3(new_n356), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n520), .A2(new_n535), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n422), .A2(KEYINPUT22), .A3(new_n222), .A4(G87), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n263), .A2(new_n222), .A3(G87), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT22), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n281), .A2(new_n485), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n222), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT23), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n548), .A2(new_n222), .A3(G107), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n548), .B1(new_n222), .B2(G107), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n545), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT24), .B1(new_n542), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT24), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n550), .A2(new_n551), .B1(new_n222), .B2(new_n546), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n541), .A2(new_n555), .A3(new_n545), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n282), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n533), .A2(G107), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n222), .A2(G107), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n293), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT88), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT25), .ZN(new_n564));
  OR2_X1    g0364(.A1(new_n563), .A2(KEYINPUT25), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(KEYINPUT25), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n565), .A2(new_n293), .A3(new_n561), .A4(new_n566), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n560), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n509), .A2(new_n265), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(G257), .B2(new_n265), .ZN(new_n570));
  INV_X1    g0370(.A(G294), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n400), .A2(new_n570), .B1(new_n281), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n321), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n479), .A2(G264), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(G190), .A3(new_n478), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n573), .A2(new_n478), .A3(new_n574), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G200), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n559), .A2(new_n568), .A3(new_n576), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n511), .A2(G1698), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G238), .B2(G1698), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n400), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n321), .B1(new_n582), .B2(new_n546), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n471), .A2(new_n509), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n473), .A2(new_n471), .B1(new_n584), .B2(new_n254), .ZN(new_n585));
  AOI21_X1  g0385(.A(G169), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n583), .A2(new_n585), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n586), .B1(new_n356), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT19), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n222), .B1(new_n316), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(G87), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(new_n526), .A3(new_n340), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n422), .A2(new_n222), .A3(G68), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n589), .B1(new_n279), .B2(new_n526), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n596), .A2(new_n282), .B1(new_n484), .B2(new_n348), .ZN(new_n597));
  INV_X1    g0397(.A(new_n348), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n533), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n588), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n583), .A2(new_n585), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G200), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n533), .A2(G87), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n583), .A2(G190), .A3(new_n585), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n597), .A2(new_n603), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n579), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n540), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n577), .A2(new_n271), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n573), .A2(new_n356), .A3(new_n478), .A4(new_n574), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n376), .B1(new_n554), .B2(new_n557), .ZN(new_n611));
  INV_X1    g0411(.A(new_n568), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT89), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n613), .B(new_n614), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n457), .A2(new_n506), .A3(new_n608), .A4(new_n615), .ZN(G372));
  OAI211_X1 g0416(.A(new_n613), .B(new_n500), .C1(new_n503), .C2(new_n504), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n608), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT26), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n517), .A2(new_n519), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n271), .ZN(new_n621));
  INV_X1    g0421(.A(new_n539), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n601), .A2(new_n606), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n619), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n536), .A2(new_n539), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n626), .A2(KEYINPUT26), .A3(new_n601), .A4(new_n606), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n618), .A2(new_n628), .A3(new_n601), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n457), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n291), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT90), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n373), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n373), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n445), .A2(new_n448), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT18), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n450), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n333), .A2(new_n362), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n337), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n639), .B1(new_n641), .B2(new_n439), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n631), .B1(new_n635), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n630), .A2(new_n643), .ZN(G369));
  OR3_X1    g0444(.A1(new_n294), .A2(KEYINPUT27), .A3(G20), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT27), .B1(new_n294), .B2(G20), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G343), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n611), .B2(new_n612), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n615), .A2(new_n579), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n649), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n613), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n652), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT91), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n613), .A2(new_n649), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n495), .A2(new_n649), .ZN(new_n660));
  MUX2_X1   g0460(.A(new_n654), .B(new_n506), .S(new_n660), .Z(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n653), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n659), .A2(new_n664), .ZN(G399));
  INV_X1    g0465(.A(new_n213), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(G41), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n592), .A2(G116), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G1), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n224), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n668), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT28), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n613), .B(KEYINPUT89), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n608), .B1(new_n674), .B2(new_n654), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n627), .A2(KEYINPUT95), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n625), .A2(KEYINPUT95), .A3(new_n627), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n675), .A2(new_n676), .A3(new_n677), .A4(new_n601), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(KEYINPUT29), .A3(new_n652), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n629), .A2(new_n652), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(KEYINPUT29), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n587), .A2(new_n575), .A3(new_n499), .A4(new_n465), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT30), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n620), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AND4_X1   g0484(.A1(new_n356), .A2(new_n516), .A3(new_n577), .A4(new_n602), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n684), .B1(new_n482), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n465), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n583), .A2(new_n573), .A3(new_n574), .A4(new_n585), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n478), .A2(new_n480), .A3(G179), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(KEYINPUT93), .A3(new_n517), .A4(new_n519), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT93), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n620), .B2(new_n682), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n691), .A2(new_n693), .A3(new_n683), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n686), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g0495(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(new_n649), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n608), .A2(new_n506), .A3(new_n615), .A4(new_n652), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT94), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n694), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n691), .A2(new_n693), .A3(KEYINPUT94), .A4(new_n683), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(new_n702), .A3(new_n686), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT31), .B1(new_n703), .B2(new_n649), .ZN(new_n704));
  OAI21_X1  g0504(.A(G330), .B1(new_n699), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n681), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT96), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n673), .B1(new_n708), .B2(G1), .ZN(G364));
  NOR2_X1   g0509(.A1(new_n284), .A2(G20), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n256), .B1(new_n710), .B2(G45), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n667), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n663), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(G330), .B2(new_n661), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n319), .A2(new_n666), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G355), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(G116), .B2(new_n213), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n422), .A2(new_n666), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n470), .B2(new_n224), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n251), .A2(G45), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n221), .B1(G20), .B2(new_n271), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n713), .B1(new_n723), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n222), .A2(G179), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(G190), .A3(G200), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT101), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(KEYINPUT101), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n222), .A2(new_n356), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n737), .A2(KEYINPUT97), .ZN(new_n738));
  AOI21_X1  g0538(.A(G200), .B1(new_n737), .B2(KEYINPUT97), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(new_n364), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G311), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n460), .A2(new_n735), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n738), .A2(new_n739), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n364), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n742), .B1(G322), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n736), .A2(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n364), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G326), .ZN(new_n749));
  INV_X1    g0549(.A(G283), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n731), .A2(new_n364), .A3(G200), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n748), .A2(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n746), .A2(G190), .ZN(new_n753));
  XNOR2_X1  g0553(.A(KEYINPUT33), .B(G317), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(G20), .A3(new_n364), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT99), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G329), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n222), .B1(new_n756), .B2(G190), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n263), .B1(new_n765), .B2(G294), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n745), .A2(new_n755), .A3(new_n763), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n744), .B(KEYINPUT98), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n202), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n263), .B1(new_n748), .B2(new_n207), .ZN(new_n771));
  INV_X1    g0571(.A(new_n753), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n772), .A2(new_n203), .B1(new_n764), .B2(new_n526), .ZN(new_n773));
  INV_X1    g0573(.A(new_n751), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n771), .B(new_n773), .C1(G107), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n735), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G87), .ZN(new_n777));
  INV_X1    g0577(.A(new_n740), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G77), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n761), .A2(new_n377), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT100), .B(KEYINPUT32), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n775), .A2(new_n777), .A3(new_n779), .A4(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n767), .B1(new_n770), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n730), .B1(new_n784), .B2(new_n724), .ZN(new_n785));
  INV_X1    g0585(.A(new_n727), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n661), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n715), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(G396));
  NAND2_X1  g0589(.A1(new_n352), .A2(new_n649), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n362), .A2(new_n365), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n357), .A2(new_n358), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n360), .A2(KEYINPUT71), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n353), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n794), .A2(KEYINPUT104), .A3(new_n649), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(KEYINPUT104), .B1(new_n794), .B2(new_n649), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n791), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n680), .B(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n713), .B1(new_n799), .B2(new_n705), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n705), .B2(new_n799), .ZN(new_n801));
  INV_X1    g0601(.A(new_n713), .ZN(new_n802));
  INV_X1    g0602(.A(new_n724), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n726), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT102), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n802), .B1(new_n806), .B2(new_n304), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n744), .A2(G294), .B1(new_n776), .B2(G107), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n485), .B2(new_n740), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n751), .A2(new_n591), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n772), .A2(new_n750), .B1(new_n748), .B2(new_n460), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n319), .B1(new_n526), .B2(new_n764), .C1(new_n761), .C2(new_n741), .ZN(new_n812));
  NOR4_X1   g0612(.A1(new_n809), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G137), .A2(new_n747), .B1(new_n753), .B2(G150), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT103), .ZN(new_n815));
  INV_X1    g0615(.A(G143), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n815), .B1(new_n377), .B2(new_n740), .C1(new_n769), .C2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT34), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n422), .B1(new_n202), .B2(new_n764), .C1(new_n203), .C2(new_n751), .ZN(new_n819));
  INV_X1    g0619(.A(G132), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n761), .A2(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n819), .B(new_n821), .C1(G50), .C2(new_n776), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n813), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n807), .B1(new_n726), .B2(new_n798), .C1(new_n823), .C2(new_n803), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n801), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G384));
  NOR2_X1   g0626(.A1(new_n710), .A2(new_n256), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n412), .A2(new_n381), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n443), .B(new_n282), .C1(KEYINPUT16), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n420), .ZN(new_n830));
  INV_X1    g0630(.A(new_n647), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n453), .B1(new_n452), .B2(KEYINPUT18), .ZN(new_n834));
  NOR4_X1   g0634(.A1(new_n435), .A2(KEYINPUT81), .A3(new_n637), .A4(new_n447), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n834), .A2(new_n835), .A3(new_n449), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n833), .B1(new_n836), .B2(new_n439), .ZN(new_n837));
  INV_X1    g0637(.A(new_n430), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n829), .A2(new_n420), .B1(new_n447), .B2(new_n647), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT37), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n445), .A2(new_n831), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT37), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n636), .A2(new_n841), .A3(new_n842), .A4(new_n430), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT38), .B1(new_n837), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n450), .A2(KEYINPUT81), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n846), .A2(new_n454), .A3(new_n638), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n433), .A2(new_n438), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n832), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n844), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT39), .B1(new_n845), .B2(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n854));
  NAND3_X1  g0654(.A1(new_n636), .A2(new_n841), .A3(new_n430), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n843), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n841), .B1(new_n848), .B2(new_n639), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n854), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(KEYINPUT38), .B(new_n844), .C1(new_n455), .C2(new_n832), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT39), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n853), .A2(KEYINPUT105), .A3(new_n863), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n333), .A2(new_n649), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n851), .B1(new_n849), .B2(new_n850), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n861), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT105), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT39), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n864), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n311), .A2(new_n649), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n333), .B2(new_n337), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n333), .A2(new_n337), .A3(new_n872), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n680), .A2(new_n798), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n794), .A2(new_n652), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n638), .A2(new_n450), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n880), .A2(new_n868), .B1(new_n881), .B2(new_n647), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n871), .A2(new_n882), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n681), .A2(new_n456), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n643), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n883), .B(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(G330), .ZN(new_n887));
  INV_X1    g0687(.A(new_n875), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n798), .B1(new_n888), .B2(new_n873), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n698), .A2(new_n696), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n703), .A2(new_n649), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n893));
  AOI211_X1 g0693(.A(KEYINPUT40), .B(new_n889), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n868), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n797), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n795), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n874), .A2(new_n875), .B1(new_n897), .B2(new_n791), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n698), .A2(new_n696), .B1(new_n703), .B2(new_n649), .ZN(new_n899));
  INV_X1    g0699(.A(new_n893), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n861), .B2(new_n860), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n895), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n456), .B1(new_n892), .B2(new_n893), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n887), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n905), .B2(new_n904), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n827), .B1(new_n886), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n886), .B2(new_n907), .ZN(new_n909));
  INV_X1    g0709(.A(new_n529), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n910), .A2(KEYINPUT35), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(KEYINPUT35), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n911), .A2(G116), .A3(new_n223), .A4(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT36), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n224), .A2(G77), .A3(new_n379), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(G50), .B2(new_n203), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(G1), .A3(new_n284), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n909), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT107), .Z(G367));
  OAI22_X1  g0719(.A1(new_n202), .A2(new_n735), .B1(new_n740), .B2(new_n207), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(G150), .B2(new_n744), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n764), .A2(new_n203), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n751), .A2(new_n304), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n922), .B(new_n923), .C1(G159), .C2(new_n753), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n263), .B1(new_n748), .B2(new_n816), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(G137), .B2(new_n762), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n921), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT113), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n776), .B2(G116), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT46), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n769), .A2(new_n460), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n778), .A2(G283), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n748), .A2(new_n741), .B1(new_n764), .B2(new_n340), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(G294), .B2(new_n753), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n400), .B1(new_n526), .B2(new_n751), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n762), .B2(G317), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n932), .A2(new_n933), .A3(new_n935), .A4(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n927), .B1(new_n931), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT47), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n724), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n652), .B1(new_n597), .B2(new_n604), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n624), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(new_n600), .A3(new_n588), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(new_n727), .A3(new_n944), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n728), .B1(new_n213), .B2(new_n348), .C1(new_n242), .C2(new_n720), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n946), .A2(KEYINPUT112), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(KEYINPUT112), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n947), .A2(new_n948), .A3(new_n802), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n941), .A2(new_n945), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n667), .B(KEYINPUT41), .Z(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n537), .A2(new_n649), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n540), .A2(new_n954), .B1(new_n623), .B2(new_n652), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT109), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n659), .A2(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT45), .Z(new_n959));
  NOR2_X1   g0759(.A1(new_n659), .A2(new_n957), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT44), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n664), .A2(KEYINPUT111), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n662), .B(new_n653), .Z(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(new_n656), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(new_n707), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n953), .B1(new_n970), .B2(new_n707), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n711), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n657), .A2(new_n957), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT110), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT42), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n623), .B1(new_n956), .B2(new_n615), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n652), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n943), .A2(new_n944), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT43), .B1(new_n979), .B2(KEYINPUT108), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(KEYINPUT108), .B2(new_n979), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n978), .A2(new_n983), .A3(new_n981), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n664), .A2(new_n956), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n985), .B(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n951), .B1(new_n972), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(G387));
  NAND2_X1  g0789(.A1(new_n967), .A2(new_n707), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n969), .A2(new_n990), .A3(new_n667), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n776), .A2(G77), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n400), .B1(G97), .B2(new_n774), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n274), .C2(new_n761), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT114), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n747), .A2(G159), .B1(new_n598), .B2(new_n765), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n278), .B2(new_n772), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G68), .B2(new_n778), .ZN(new_n998));
  INV_X1    g0798(.A(new_n744), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n995), .B(new_n998), .C1(new_n207), .C2(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n776), .A2(G294), .B1(G283), .B2(new_n765), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G311), .A2(new_n753), .B1(new_n747), .B2(G322), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n460), .B2(new_n740), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n768), .B2(G317), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1001), .B1(new_n1004), .B2(KEYINPUT48), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(KEYINPUT48), .B2(new_n1004), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT49), .Z(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(KEYINPUT115), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n400), .B1(new_n485), .B2(new_n751), .C1(new_n761), .C2(new_n749), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT116), .Z(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1007), .A2(KEYINPUT115), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1000), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n724), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n669), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n716), .A2(new_n1015), .B1(new_n340), .B2(new_n666), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n239), .A2(new_n470), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n277), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n207), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT50), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n669), .B(new_n470), .C1(new_n203), .C2(new_n304), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n719), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1016), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n802), .B1(new_n1023), .B2(new_n728), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1014), .B(new_n1024), .C1(new_n653), .C2(new_n786), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n991), .B(new_n1025), .C1(new_n711), .C2(new_n967), .ZN(G393));
  NAND3_X1  g0826(.A1(new_n962), .A2(new_n663), .A3(new_n653), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n959), .A2(new_n664), .A3(new_n961), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1027), .A2(new_n712), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n246), .A2(new_n720), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n728), .B1(new_n526), .B2(new_n213), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n319), .B1(new_n751), .B2(new_n340), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n772), .A2(new_n460), .B1(new_n764), .B2(new_n485), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(G322), .C2(new_n762), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n750), .B2(new_n735), .C1(new_n571), .C2(new_n740), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n744), .A2(G311), .B1(G317), .B2(new_n747), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT52), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n772), .A2(new_n207), .B1(new_n764), .B2(new_n304), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n400), .B(new_n810), .C1(new_n762), .C2(G143), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n203), .B2(new_n735), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT117), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1039), .B(new_n1042), .C1(new_n1018), .C2(new_n778), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n744), .A2(G159), .B1(G150), .B2(new_n747), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT51), .Z(new_n1045));
  AOI21_X1  g0845(.A(new_n1038), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n713), .B1(new_n1030), .B2(new_n1031), .C1(new_n1046), .C2(new_n803), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n956), .B2(new_n727), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1029), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT118), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n968), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1052));
  OR3_X1    g0852(.A1(new_n970), .A2(new_n668), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(G390));
  AOI21_X1  g0854(.A(new_n887), .B1(new_n892), .B2(new_n893), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n898), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n880), .A2(new_n866), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n864), .B2(new_n870), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n678), .A2(new_n652), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n798), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n879), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n866), .B1(new_n1062), .B2(new_n876), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n860), .A2(new_n861), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1057), .B1(new_n1059), .B2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n898), .B(G330), .C1(new_n699), .C2(new_n704), .ZN(new_n1068));
  AOI211_X1 g0868(.A(KEYINPUT105), .B(new_n862), .C1(new_n867), .C2(new_n861), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n869), .B1(new_n868), .B2(KEYINPUT39), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1069), .B1(new_n863), .B2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1068), .B(new_n1065), .C1(new_n1071), .C2(new_n1058), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n457), .A2(new_n1055), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n884), .A2(new_n1074), .A3(new_n643), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1068), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1076), .A2(new_n1062), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n892), .A2(new_n893), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1078), .A2(G330), .A3(new_n798), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n877), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1077), .A2(new_n1080), .A3(KEYINPUT119), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT119), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1068), .B(new_n879), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n876), .B1(new_n1055), .B2(new_n798), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n877), .B1(new_n705), .B2(new_n1061), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n1056), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n878), .A2(new_n879), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1075), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1073), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1067), .A2(new_n1072), .A3(new_n1091), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n667), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1067), .A2(new_n1072), .A3(new_n712), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n802), .B1(new_n806), .B2(new_n278), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n777), .B1(new_n526), .B2(new_n740), .C1(new_n999), .C2(new_n485), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n753), .A2(G107), .B1(G77), .B2(new_n765), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n750), .B2(new_n748), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n319), .B1(new_n203), .B2(new_n751), .C1(new_n761), .C2(new_n571), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n753), .A2(G137), .B1(G159), .B2(new_n765), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n747), .A2(G128), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1103), .B(new_n1104), .C1(new_n740), .C2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n263), .B1(new_n751), .B2(new_n207), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n762), .B2(G125), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT120), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1106), .B(new_n1109), .C1(G132), .C2(new_n744), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n735), .A2(new_n274), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT53), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1102), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1097), .B1(new_n1113), .B2(new_n803), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT121), .Z(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n1071), .B2(new_n726), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1095), .A2(new_n1096), .A3(new_n1116), .ZN(G378));
  NAND2_X1  g0917(.A1(new_n635), .A2(new_n291), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n290), .A2(new_n831), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n635), .A2(new_n291), .A3(new_n1119), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1123), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1119), .B1(new_n635), .B2(new_n291), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n631), .B(new_n1120), .C1(new_n633), .C2(new_n634), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n904), .A2(G330), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n904), .B2(G330), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n883), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n854), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n841), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n881), .B2(new_n439), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1134), .B1(new_n1136), .B2(new_n857), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1078), .B(new_n898), .C1(new_n852), .C2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1138), .A2(KEYINPUT40), .B1(new_n868), .B2(new_n894), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1133), .B1(new_n1139), .B2(new_n887), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n904), .A2(G330), .A3(new_n1129), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1140), .A2(new_n871), .A3(new_n882), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1132), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n712), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n802), .B1(new_n806), .B2(new_n207), .ZN(new_n1145));
  INV_X1    g0945(.A(G137), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n735), .A2(new_n1105), .B1(new_n740), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n747), .A2(G125), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n753), .A2(G132), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n765), .A2(G150), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1147), .B(new_n1151), .C1(G128), .C2(new_n744), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n762), .A2(G124), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G33), .B(G41), .C1(new_n774), .C2(G159), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n992), .B1(new_n999), .B2(new_n340), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n772), .A2(new_n526), .B1(new_n202), .B2(new_n751), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n922), .B(new_n1160), .C1(G116), .C2(new_n747), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n422), .A2(G41), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1161), .B(new_n1162), .C1(new_n750), .C2(new_n761), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1159), .B(new_n1163), .C1(new_n598), .C2(new_n778), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(KEYINPUT58), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(KEYINPUT58), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1162), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1167), .B(new_n207), .C1(G33), .C2(G41), .ZN(new_n1168));
  AND4_X1   g0968(.A1(new_n1158), .A2(new_n1165), .A3(new_n1166), .A4(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1145), .B1(new_n803), .B2(new_n1169), .C1(new_n1129), .C2(new_n726), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1144), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1075), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1094), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n1143), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT57), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1132), .B2(new_n1142), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n668), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1171), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(G375));
  NAND3_X1  g0980(.A1(new_n1086), .A2(new_n1090), .A3(new_n1075), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1092), .A2(new_n953), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n711), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n877), .A2(new_n725), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n713), .B1(new_n805), .B2(G68), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n999), .A2(new_n750), .B1(new_n340), .B2(new_n740), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G97), .B2(new_n776), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n747), .A2(G294), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n753), .A2(G116), .B1(new_n598), .B2(new_n765), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n263), .B(new_n923), .C1(new_n762), .C2(G303), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n769), .A2(new_n1146), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G159), .A2(new_n776), .B1(new_n778), .B2(G150), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n748), .A2(new_n820), .B1(new_n764), .B2(new_n207), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1105), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n753), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n422), .B1(new_n202), .B2(new_n751), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n762), .B2(G128), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1193), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1191), .B1(new_n1192), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1185), .B1(new_n1200), .B2(new_n724), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1183), .B1(new_n1184), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1182), .A2(new_n1202), .ZN(G381));
  NOR3_X1   g1003(.A1(G387), .A2(G390), .A3(G381), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT122), .ZN(new_n1206));
  INV_X1    g1006(.A(G378), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1206), .A3(new_n1207), .A4(new_n1179), .ZN(G407));
  NAND2_X1  g1008(.A1(new_n648), .A2(G213), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1179), .A2(new_n1207), .A3(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(G407), .A2(G213), .A3(new_n1211), .ZN(G409));
  NOR2_X1   g1012(.A1(new_n988), .A2(G390), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT125), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n988), .A2(G390), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(G393), .B(new_n788), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1216), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1215), .B1(new_n988), .B2(G390), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1217), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n1219), .A2(new_n1213), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT61), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1218), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1174), .A2(new_n952), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1207), .B1(new_n1171), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT123), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1179), .B2(G378), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1173), .A2(new_n1177), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1094), .A2(new_n1172), .B1(new_n1142), .B2(new_n1132), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1229), .B(new_n667), .C1(KEYINPUT57), .C2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1171), .ZN(new_n1232));
  AND4_X1   g1032(.A1(new_n1227), .A2(new_n1231), .A3(G378), .A4(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1226), .B1(new_n1228), .B2(new_n1233), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1234), .A2(new_n1209), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1092), .A2(KEYINPUT60), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1236), .A2(new_n1181), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n667), .B1(new_n1236), .B2(new_n1181), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1202), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1239), .A2(new_n825), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n825), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT63), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1224), .B1(new_n1235), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1234), .A2(KEYINPUT124), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1242), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT124), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1226), .B(new_n1248), .C1(new_n1228), .C2(new_n1233), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1246), .A2(new_n1209), .A3(new_n1247), .A4(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1243), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1246), .A2(new_n1209), .A3(new_n1249), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1210), .A2(G2897), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1242), .B(new_n1253), .Z(new_n1254));
  OAI211_X1 g1054(.A(new_n1245), .B(new_n1251), .C1(new_n1252), .C2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1223), .B1(new_n1254), .B2(new_n1235), .ZN(new_n1256));
  AND4_X1   g1056(.A1(KEYINPUT62), .A2(new_n1234), .A3(new_n1209), .A4(new_n1247), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1250), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1257), .B1(new_n1259), .B2(KEYINPUT126), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT126), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1250), .A2(new_n1261), .A3(new_n1258), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1256), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1218), .A2(new_n1222), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(KEYINPUT127), .Z(new_n1265));
  OAI21_X1  g1065(.A(new_n1255), .B1(new_n1263), .B2(new_n1265), .ZN(G405));
  OAI22_X1  g1066(.A1(new_n1228), .A2(new_n1233), .B1(G378), .B2(new_n1179), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(new_n1247), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1268), .B(new_n1264), .ZN(G402));
endmodule


