//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  AOI211_X1 g0011(.A(new_n205), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n212), .A2(KEYINPUT0), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n218), .B1(KEYINPUT0), .B2(new_n212), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n202), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  INV_X1    g0025(.A(G97), .ZN(new_n226));
  INV_X1    g0026(.A(G107), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n225), .B1(new_n226), .B2(new_n210), .C1(new_n227), .C2(new_n211), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n207), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n219), .A2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  XNOR2_X1  g0047(.A(KEYINPUT65), .B(G41), .ZN(new_n248));
  INV_X1    g0048(.A(G45), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G274), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G1), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT66), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT66), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n250), .A2(new_n255), .A3(new_n252), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n254), .A2(new_n256), .B1(G244), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT67), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n257), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(KEYINPUT67), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G1698), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n275), .A2(G232), .B1(G107), .B2(new_n274), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n269), .A2(new_n273), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G1698), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT68), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n278), .B(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n276), .B1(new_n280), .B2(new_n222), .ZN(new_n281));
  INV_X1    g0081(.A(new_n259), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n265), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n283), .A2(G169), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G20), .A2(G77), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n214), .A2(G33), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT15), .B(G87), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n285), .B1(new_n286), .B2(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n213), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n202), .ZN(new_n297));
  INV_X1    g0097(.A(new_n293), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(G1), .B2(new_n214), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n297), .B1(new_n299), .B2(new_n202), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G179), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n283), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n284), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n254), .A2(new_n256), .ZN(new_n305));
  INV_X1    g0105(.A(G226), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(new_n262), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n278), .B(KEYINPUT68), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G223), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n275), .A2(G222), .B1(G77), .B2(new_n274), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n302), .B(new_n308), .C1(new_n312), .C2(new_n259), .ZN(new_n313));
  INV_X1    g0113(.A(new_n299), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G50), .ZN(new_n315));
  INV_X1    g0115(.A(G150), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n316), .A2(new_n288), .B1(new_n201), .B2(new_n214), .ZN(new_n317));
  XOR2_X1   g0117(.A(new_n286), .B(KEYINPUT69), .Z(new_n318));
  INV_X1    g0118(.A(KEYINPUT70), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n289), .B(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n317), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n315), .B1(G50), .B2(new_n295), .C1(new_n321), .C2(new_n298), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n259), .B1(new_n310), .B2(new_n311), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n307), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n313), .B(new_n322), .C1(G169), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n320), .A2(G77), .ZN(new_n326));
  INV_X1    g0126(.A(G50), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n326), .B1(new_n214), .B2(G68), .C1(new_n327), .C2(new_n288), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n293), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT11), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n296), .A2(new_n221), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT12), .B1(new_n332), .B2(KEYINPUT71), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(KEYINPUT71), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n332), .A2(KEYINPUT71), .A3(KEYINPUT12), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n335), .A2(new_n336), .B1(G68), .B2(new_n314), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n328), .A2(KEYINPUT11), .A3(new_n293), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n331), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n263), .A2(G238), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n305), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(G226), .A2(G1698), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n235), .B2(G1698), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n277), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n257), .A2(new_n226), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n259), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT13), .B1(new_n341), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n347), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n254), .A2(new_n256), .B1(G238), .B2(new_n263), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n339), .B1(G200), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G190), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n354), .B1(new_n355), .B2(new_n353), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n283), .A2(G190), .ZN(new_n357));
  INV_X1    g0157(.A(G200), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n357), .B(new_n301), .C1(new_n358), .C2(new_n283), .ZN(new_n359));
  AND4_X1   g0159(.A1(new_n304), .A2(new_n325), .A3(new_n356), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n324), .A2(G190), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n322), .B(KEYINPUT9), .ZN(new_n362));
  OAI21_X1  g0162(.A(G200), .B1(new_n323), .B2(new_n307), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT10), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT10), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n361), .A2(new_n366), .A3(new_n362), .A4(new_n363), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n348), .A2(new_n352), .A3(G179), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT72), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n348), .A2(new_n352), .A3(KEYINPUT72), .A4(G179), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n353), .A2(G169), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT14), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT14), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n353), .A2(new_n376), .A3(G169), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n373), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n339), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n360), .A2(new_n368), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n306), .A2(G1698), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(G223), .B2(G1698), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n267), .A2(new_n268), .ZN(new_n383));
  INV_X1    g0183(.A(G87), .ZN(new_n384));
  OAI22_X1  g0184(.A1(new_n382), .A2(new_n383), .B1(new_n257), .B2(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(new_n282), .B1(new_n263), .B2(G232), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n305), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(new_n355), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(G200), .B2(new_n387), .ZN(new_n389));
  INV_X1    g0189(.A(new_n318), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n296), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n390), .B2(new_n299), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G58), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(new_n221), .ZN(new_n395));
  NOR2_X1   g0195(.A1(G58), .A2(G68), .ZN(new_n396));
  OAI21_X1  g0196(.A(G20), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n287), .A2(G159), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n383), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n400));
  AOI21_X1  g0200(.A(G20), .B1(new_n269), .B2(new_n273), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(KEYINPUT7), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G68), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n399), .B1(new_n403), .B2(KEYINPUT74), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT74), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(new_n405), .A3(G68), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT16), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT73), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT7), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n271), .A2(new_n272), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(G20), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n221), .B1(new_n411), .B2(new_n400), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(new_n399), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n408), .B1(new_n413), .B2(KEYINPUT16), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT16), .ZN(new_n415));
  NOR4_X1   g0215(.A1(new_n412), .A2(KEYINPUT73), .A3(new_n399), .A4(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n293), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n389), .B(new_n393), .C1(new_n407), .C2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT17), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n418), .B(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n393), .B1(new_n407), .B2(new_n417), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n387), .A2(G169), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n302), .B2(new_n387), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT18), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n421), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n420), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n380), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT6), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n432), .A2(new_n226), .A3(G107), .ZN(new_n433));
  XNOR2_X1  g0233(.A(G97), .B(G107), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n433), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n435), .A2(new_n214), .B1(new_n202), .B2(new_n288), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n402), .A2(G107), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n436), .B1(new_n437), .B2(KEYINPUT75), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT75), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n402), .A2(new_n439), .A3(G107), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n298), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n295), .A2(G97), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n257), .A2(G1), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n296), .A2(new_n293), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n442), .B1(new_n444), .B2(G97), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT76), .B1(new_n441), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n249), .A2(G1), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n258), .A2(KEYINPUT5), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n448), .B(new_n449), .C1(new_n248), .C2(KEYINPUT5), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(G257), .A3(new_n259), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT80), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT80), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n450), .A2(new_n453), .A3(G257), .A4(new_n259), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT5), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT79), .B1(new_n456), .B2(G41), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT79), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(new_n258), .A3(KEYINPUT5), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(G274), .A3(new_n259), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n258), .A2(KEYINPUT65), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT65), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G41), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n456), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT78), .B1(new_n467), .B2(new_n448), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT5), .B1(new_n463), .B2(new_n465), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT78), .ZN(new_n470));
  INV_X1    g0270(.A(new_n448), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n462), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT4), .ZN(new_n474));
  INV_X1    g0274(.A(G1698), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(new_n475), .A3(G244), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n383), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n223), .A2(G1698), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n269), .A2(new_n273), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n477), .B1(new_n479), .B2(KEYINPUT4), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n269), .A2(new_n273), .A3(G250), .A4(G1698), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT77), .B1(G33), .B2(G283), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(KEYINPUT77), .A2(G33), .A3(G283), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n282), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n455), .A2(new_n473), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G200), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n455), .A2(new_n487), .A3(G190), .A4(new_n473), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT76), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n402), .A2(new_n439), .A3(G107), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n439), .B1(new_n402), .B2(G107), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n493), .A2(new_n494), .A3(new_n436), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n492), .B(new_n445), .C1(new_n495), .C2(new_n298), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n447), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n290), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n444), .A2(new_n498), .ZN(new_n499));
  XOR2_X1   g0299(.A(new_n499), .B(KEYINPUT81), .Z(new_n500));
  NAND3_X1  g0300(.A1(new_n410), .A2(new_n214), .A3(G68), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n384), .A2(new_n226), .A3(new_n227), .ZN(new_n502));
  OAI211_X1 g0302(.A(KEYINPUT19), .B(new_n502), .C1(new_n345), .C2(G20), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n289), .A2(new_n226), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n501), .B(new_n503), .C1(KEYINPUT19), .C2(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n505), .A2(new_n293), .B1(new_n296), .B2(new_n290), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n260), .A2(new_n251), .A3(G45), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n205), .B1(new_n249), .B2(G1), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n259), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n223), .A2(G1698), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(G238), .B2(G1698), .ZN(new_n512));
  INV_X1    g0312(.A(G116), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n512), .A2(new_n383), .B1(new_n257), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n510), .B1(new_n514), .B2(new_n282), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(G169), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n302), .B2(new_n515), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n515), .A2(new_n358), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n518), .B1(G190), .B2(new_n515), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n444), .A2(G87), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n506), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n507), .A2(new_n517), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n488), .A2(G169), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n302), .B2(new_n488), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n445), .B1(new_n495), .B2(new_n298), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n497), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n450), .A2(G264), .A3(new_n259), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n210), .A2(G1698), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(G250), .B2(G1698), .ZN(new_n530));
  INV_X1    g0330(.A(G294), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n530), .A2(new_n383), .B1(new_n257), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n282), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n473), .A2(new_n528), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(new_n355), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(G200), .B2(new_n534), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n410), .A2(KEYINPUT22), .A3(new_n214), .A4(G87), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n227), .A2(G20), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT23), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n214), .A2(G33), .A3(G116), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n537), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT22), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n214), .A2(G87), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n543), .B1(new_n274), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT24), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT24), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n542), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n298), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n444), .A2(G107), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n296), .A2(new_n227), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n552), .B(KEYINPUT84), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n553), .A2(KEYINPUT25), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(KEYINPUT25), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n536), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G169), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n534), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n473), .A2(new_n528), .A3(new_n533), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n302), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n560), .B(new_n562), .C1(new_n550), .C2(new_n556), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n450), .A2(G270), .A3(new_n259), .ZN(new_n565));
  INV_X1    g0365(.A(G303), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n269), .B2(new_n273), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n211), .A2(G1698), .ZN(new_n568));
  OAI221_X1 g0368(.A(new_n568), .B1(G257), .B2(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n282), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n473), .A2(new_n565), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT20), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n214), .B1(new_n226), .B2(G33), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n483), .B2(new_n484), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n513), .A2(G20), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n293), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n573), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(G20), .B1(new_n257), .B2(G97), .ZN(new_n579));
  INV_X1    g0379(.A(new_n484), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n579), .B1(new_n580), .B2(new_n482), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n581), .A2(KEYINPUT20), .A3(new_n293), .A4(new_n576), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n295), .A2(G116), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n444), .B2(G116), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n559), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n572), .A2(new_n586), .A3(KEYINPUT21), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT82), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n572), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n583), .A2(new_n585), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(G179), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n572), .A2(new_n586), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n589), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n572), .A2(new_n586), .A3(KEYINPUT82), .A4(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n590), .A2(G190), .ZN(new_n598));
  INV_X1    g0398(.A(new_n591), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n572), .A2(G200), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n596), .A2(KEYINPUT83), .A3(new_n597), .A4(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT83), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n589), .A2(new_n592), .A3(new_n595), .A4(new_n597), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  AND4_X1   g0407(.A1(new_n431), .A2(new_n527), .A3(new_n564), .A4(new_n607), .ZN(G372));
  INV_X1    g0408(.A(new_n325), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n365), .A2(new_n367), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n356), .A2(new_n284), .A3(new_n303), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n379), .ZN(new_n612));
  INV_X1    g0412(.A(new_n420), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n428), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT88), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n610), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n420), .B1(new_n611), .B2(new_n379), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT88), .B1(new_n617), .B2(new_n428), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n609), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n431), .ZN(new_n620));
  XOR2_X1   g0420(.A(new_n563), .B(KEYINPUT85), .Z(new_n621));
  OAI211_X1 g0421(.A(new_n527), .B(new_n558), .C1(new_n621), .C2(new_n604), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n467), .A2(KEYINPUT78), .A3(new_n448), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n470), .B1(new_n469), .B2(new_n471), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n461), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n479), .A2(KEYINPUT4), .ZN(new_n626));
  INV_X1    g0426(.A(new_n477), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n481), .A2(new_n485), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n625), .B1(new_n630), .B2(new_n282), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n559), .B1(new_n631), .B2(new_n455), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n488), .A2(new_n302), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT86), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT86), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n523), .B(new_n635), .C1(new_n302), .C2(new_n488), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n447), .A2(new_n496), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .A4(new_n522), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n507), .A2(new_n517), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n524), .A2(new_n522), .A3(new_n525), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n641), .B1(new_n642), .B2(KEYINPUT26), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT87), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n640), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n640), .B2(new_n643), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n622), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n619), .B1(new_n620), .B2(new_n648), .ZN(G369));
  INV_X1    g0449(.A(G330), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n260), .A2(new_n214), .A3(G13), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G343), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n604), .A2(new_n591), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g0457(.A(new_n657), .B(KEYINPUT89), .Z(new_n658));
  INV_X1    g0458(.A(new_n656), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n607), .B1(new_n599), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n650), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n564), .B1(new_n557), .B2(new_n659), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n563), .B2(new_n659), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT90), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n621), .A2(new_n659), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n604), .A2(new_n659), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n564), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n666), .A2(new_n671), .ZN(G399));
  NOR2_X1   g0472(.A1(new_n209), .A2(new_n466), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n502), .A2(G116), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n673), .A2(new_n260), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n217), .B2(new_n673), .ZN(new_n676));
  XOR2_X1   g0476(.A(new_n676), .B(KEYINPUT28), .Z(new_n677));
  NAND4_X1  g0477(.A1(new_n527), .A2(new_n607), .A3(new_n564), .A4(new_n659), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT30), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n515), .A2(new_n528), .A3(new_n533), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT91), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n515), .A2(KEYINPUT91), .A3(new_n533), .A4(new_n528), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n590), .A2(new_n682), .A3(G179), .A4(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n679), .B1(new_n684), .B2(new_n488), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n561), .A2(G179), .A3(new_n515), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n686), .A2(new_n488), .A3(new_n572), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n473), .A2(G179), .A3(new_n571), .A4(new_n565), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n681), .B2(new_n680), .ZN(new_n689));
  INV_X1    g0489(.A(new_n488), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(KEYINPUT30), .A3(new_n690), .A4(new_n683), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n685), .A2(new_n687), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n656), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT31), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(new_n695), .A3(new_n656), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n678), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  INV_X1    g0499(.A(new_n646), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n640), .A2(new_n643), .A3(new_n644), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n656), .B1(new_n702), .B2(new_n622), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(KEYINPUT29), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n637), .A2(new_n638), .A3(KEYINPUT26), .A4(new_n522), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT92), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n634), .A2(new_n636), .B1(new_n447), .B2(new_n496), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(KEYINPUT92), .A3(KEYINPUT26), .A4(new_n522), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n642), .A2(new_n639), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n592), .A2(new_n595), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n563), .A3(new_n597), .A4(new_n589), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n536), .A2(new_n557), .B1(new_n521), .B2(new_n519), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n497), .A2(new_n526), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n641), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n656), .B1(new_n711), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT29), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n699), .B1(new_n704), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n677), .B1(new_n723), .B2(G1), .ZN(G364));
  INV_X1    g0524(.A(new_n661), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n214), .A2(G13), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n260), .B1(new_n726), .B2(G45), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n673), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n658), .A2(new_n660), .A3(new_n650), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n725), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n658), .A2(new_n660), .A3(new_n735), .ZN(new_n736));
  OAI211_X1 g0536(.A(G1), .B(G13), .C1(new_n214), .C2(G169), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT94), .Z(new_n738));
  NOR2_X1   g0538(.A1(new_n214), .A2(G190), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G179), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G159), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n741), .A2(KEYINPUT32), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT32), .ZN(new_n744));
  INV_X1    g0544(.A(new_n741), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n744), .B1(new_n745), .B2(G159), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n214), .B1(new_n740), .B2(G190), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n743), .B(new_n746), .C1(G97), .C2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT95), .B1(new_n750), .B2(G190), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n750), .A2(KEYINPUT95), .A3(G190), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G68), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n214), .A2(new_n355), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n358), .A2(G179), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G87), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n739), .A2(new_n758), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(new_n227), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n302), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n757), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n739), .A2(new_n764), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n765), .A2(new_n394), .B1(new_n766), .B2(new_n202), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n750), .A2(new_n355), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n274), .B1(new_n769), .B2(G50), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n749), .A2(new_n756), .A3(new_n768), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT33), .B(G317), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n755), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G322), .ZN(new_n774));
  INV_X1    g0574(.A(G329), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n765), .A2(new_n774), .B1(new_n741), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n766), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n776), .B1(G311), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G283), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n759), .A2(new_n566), .B1(new_n762), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n277), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n748), .A2(G294), .B1(G326), .B2(new_n769), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n773), .A2(new_n778), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n738), .B1(new_n771), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n209), .A2(new_n410), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(G45), .B2(new_n216), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(G45), .B2(new_n243), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n209), .A2(new_n274), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(G355), .B(KEYINPUT93), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n790), .B1(G116), .B2(new_n208), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n738), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n735), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n730), .B(new_n784), .C1(new_n792), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n736), .A2(new_n795), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n732), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(G396));
  OAI21_X1  g0598(.A(new_n656), .B1(new_n294), .B2(new_n300), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n359), .A2(new_n799), .B1(new_n303), .B2(new_n284), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n284), .A2(new_n303), .A3(new_n659), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n703), .B(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n729), .B1(new_n804), .B2(new_n699), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n699), .B2(new_n804), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n738), .A2(new_n734), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT96), .Z(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT97), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n729), .B1(new_n809), .B2(G77), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n769), .A2(G137), .ZN(new_n811));
  INV_X1    g0611(.A(new_n765), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G143), .A2(new_n812), .B1(new_n777), .B2(G159), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n811), .B(new_n813), .C1(new_n754), .C2(new_n316), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT34), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n759), .A2(new_n327), .B1(new_n741), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n762), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(G68), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n410), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n817), .B(new_n820), .C1(G58), .C2(new_n748), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n755), .A2(G283), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n765), .A2(new_n531), .B1(new_n741), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G116), .B2(new_n777), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n759), .A2(new_n227), .B1(new_n762), .B2(new_n384), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n277), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n748), .A2(G97), .B1(G303), .B2(new_n769), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n823), .A2(new_n826), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n738), .B1(new_n822), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n810), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n803), .B2(new_n734), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n806), .A2(new_n833), .ZN(G384));
  INV_X1    g0634(.A(new_n435), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n835), .A2(KEYINPUT35), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(KEYINPUT35), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n836), .A2(G116), .A3(new_n215), .A4(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT36), .Z(new_n839));
  OAI211_X1 g0639(.A(new_n217), .B(G77), .C1(new_n394), .C2(new_n221), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n327), .A2(G68), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n260), .B(G13), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n647), .A2(new_n659), .A3(new_n803), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n801), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n379), .A2(KEYINPUT98), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT98), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n378), .A2(new_n847), .A3(new_n339), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n339), .A2(new_n656), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n356), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n846), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n378), .A2(new_n339), .A3(new_n656), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n845), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT99), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n404), .A2(new_n406), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n415), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n413), .A2(KEYINPUT16), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT73), .ZN(new_n860));
  INV_X1    g0660(.A(new_n416), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n298), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n392), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n413), .A2(KEYINPUT16), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n393), .B1(new_n417), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n422), .B(new_n654), .C1(new_n302), .C2(new_n387), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n863), .A2(new_n389), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n856), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n865), .A2(new_n866), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n418), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(KEYINPUT99), .A3(KEYINPUT37), .ZN(new_n872));
  INV_X1    g0672(.A(new_n654), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n421), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n424), .A2(new_n874), .A3(new_n868), .A4(new_n418), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n869), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n865), .A2(new_n873), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n420), .B2(new_n428), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n876), .A2(new_n878), .A3(KEYINPUT38), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT38), .B1(new_n876), .B2(new_n878), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n428), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n855), .A2(new_n882), .B1(new_n883), .B2(new_n873), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n846), .A2(new_n848), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n659), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n424), .A2(new_n874), .A3(new_n418), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(KEYINPUT100), .A3(new_n875), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n875), .A2(KEYINPUT100), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n889), .B(new_n890), .C1(new_n429), .C2(new_n874), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n879), .A2(KEYINPUT101), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT39), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT101), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n876), .A2(new_n878), .A3(new_n896), .A4(KEYINPUT38), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT39), .B1(new_n880), .B2(new_n881), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n886), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n884), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n720), .B(new_n431), .C1(new_n703), .C2(KEYINPUT29), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n619), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n901), .B(new_n903), .Z(new_n904));
  NAND3_X1  g0704(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n678), .A2(KEYINPUT102), .A3(new_n697), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT102), .B1(new_n678), .B2(new_n697), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n359), .A2(new_n799), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n304), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n801), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n851), .B2(new_n852), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n905), .A2(new_n909), .A3(KEYINPUT40), .A4(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT40), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n913), .B1(new_n906), .B2(new_n907), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n915), .B1(new_n916), .B2(new_n882), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n620), .B2(new_n908), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n914), .A2(new_n917), .A3(new_n431), .A4(new_n909), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(G330), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n904), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n260), .B2(new_n726), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n904), .A2(new_n921), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n843), .B1(new_n923), .B2(new_n924), .ZN(G367));
  AOI21_X1  g0725(.A(new_n716), .B1(new_n638), .B2(new_n656), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT103), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n708), .A2(new_n656), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n669), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT42), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n931), .B(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n929), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n526), .B1(new_n934), .B2(new_n563), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n659), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n522), .B1(new_n521), .B2(new_n659), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n521), .A2(new_n659), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n641), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT43), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n937), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n933), .A2(new_n943), .A3(new_n936), .A4(new_n942), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n666), .A2(new_n934), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n946), .A2(new_n947), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n666), .B2(new_n934), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n673), .B(KEYINPUT41), .Z(new_n952));
  INV_X1    g0752(.A(KEYINPUT44), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n934), .B2(new_n670), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n929), .A2(KEYINPUT44), .A3(new_n671), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT45), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n934), .B2(new_n670), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n929), .A2(KEYINPUT45), .A3(new_n671), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n665), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n669), .B1(new_n663), .B2(new_n668), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n725), .B2(KEYINPUT104), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT104), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n661), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n964), .B(new_n966), .Z(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(new_n722), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n956), .A2(new_n960), .A3(new_n666), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n962), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n952), .B1(new_n970), .B2(new_n723), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n949), .B(new_n951), .C1(new_n971), .C2(new_n728), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n274), .B1(G77), .B2(new_n818), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT106), .ZN(new_n974));
  AOI22_X1  g0774(.A1(G58), .A2(new_n760), .B1(new_n745), .B2(G137), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n975), .B1(new_n327), .B2(new_n766), .C1(new_n316), .C2(new_n765), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n754), .A2(new_n742), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n769), .A2(G143), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n221), .B2(new_n747), .ZN(new_n979));
  NOR4_X1   g0779(.A1(new_n974), .A2(new_n976), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT107), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n410), .B1(new_n745), .B2(G317), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n226), .B2(new_n762), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT105), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n765), .A2(new_n566), .B1(new_n766), .B2(new_n779), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n760), .A2(KEYINPUT46), .A3(G116), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT46), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n759), .B2(new_n513), .ZN(new_n988));
  INV_X1    g0788(.A(new_n769), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n986), .B(new_n988), .C1(new_n989), .C2(new_n824), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n985), .B(new_n990), .C1(G107), .C2(new_n748), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n531), .B2(new_n754), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n981), .B1(new_n984), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT47), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n738), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n994), .B2(new_n993), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n735), .B(new_n793), .C1(new_n209), .C2(new_n498), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n785), .A2(new_n239), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n730), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n735), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n996), .B(new_n999), .C1(new_n1000), .C2(new_n941), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n972), .A2(new_n1001), .ZN(G387));
  INV_X1    g0802(.A(new_n673), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n968), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n967), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(new_n723), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n785), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n236), .B2(G45), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n674), .B2(new_n788), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n286), .A2(G50), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT50), .Z(new_n1011));
  OAI21_X1  g0811(.A(new_n249), .B1(new_n221), .B2(new_n202), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n1011), .A2(new_n674), .A3(new_n1012), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1009), .A2(new_n1013), .B1(G107), .B2(new_n208), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n794), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n729), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n663), .A2(new_n1000), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n383), .B1(new_n818), .B2(G97), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(KEYINPUT108), .B(G150), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1018), .B1(new_n202), .B2(new_n759), .C1(new_n741), .C2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT109), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n747), .A2(new_n290), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n765), .A2(new_n327), .B1(new_n766), .B2(new_n221), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(G159), .C2(new_n769), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1021), .B(new_n1024), .C1(new_n390), .C2(new_n754), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n410), .B1(new_n745), .B2(G326), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n759), .A2(new_n531), .B1(new_n747), .B2(new_n779), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G317), .A2(new_n812), .B1(new_n777), .B2(G303), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n774), .B2(new_n989), .C1(new_n754), .C2(new_n824), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT48), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n1030), .B2(new_n1029), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1026), .B1(new_n513), .B2(new_n762), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1025), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1016), .B(new_n1017), .C1(new_n793), .C2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n1005), .B2(new_n728), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1006), .A2(new_n1038), .ZN(G393));
  NAND3_X1  g0839(.A1(new_n962), .A2(new_n728), .A3(new_n969), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n794), .B1(new_n226), .B2(new_n208), .C1(new_n1007), .C2(new_n246), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n729), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT110), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n410), .B1(new_n747), .B2(new_n202), .C1(new_n384), .C2(new_n762), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G68), .A2(new_n760), .B1(new_n745), .B2(G143), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n286), .B2(new_n766), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1044), .B(new_n1046), .C1(G50), .C2(new_n755), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n989), .A2(new_n316), .B1(new_n765), .B2(new_n742), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT51), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n754), .A2(new_n566), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n274), .B1(new_n513), .B2(new_n747), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n762), .A2(new_n227), .B1(new_n741), .B2(new_n774), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n759), .A2(new_n779), .B1(new_n766), .B2(new_n531), .ZN(new_n1053));
  NOR4_X1   g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n812), .A2(G311), .B1(G317), .B2(new_n769), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT52), .Z(new_n1056));
  AOI22_X1  g0856(.A1(new_n1047), .A2(new_n1049), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1043), .B1(new_n738), .B2(new_n1057), .C1(new_n929), .C2(new_n1000), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1040), .A2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n970), .A2(new_n673), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n962), .A2(new_n969), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n722), .B2(new_n967), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1059), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(G390));
  INV_X1    g0864(.A(KEYINPUT112), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n656), .B(new_n800), .C1(new_n711), .C2(new_n718), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n1066), .B2(new_n802), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n711), .A2(new_n718), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1068), .A2(new_n659), .A3(new_n911), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1069), .A2(KEYINPUT112), .A3(new_n801), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1067), .A2(new_n854), .A3(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n892), .A2(new_n891), .B1(new_n879), .B2(KEYINPUT101), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n886), .A2(KEYINPUT111), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT111), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n885), .A2(new_n1074), .A3(new_n659), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1072), .A2(new_n897), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n853), .B1(new_n844), .B2(new_n801), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n886), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n899), .B(new_n898), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n698), .A2(G330), .A3(new_n803), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n853), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1077), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n431), .B(G330), .C1(new_n907), .C2(new_n906), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n902), .A2(new_n619), .A3(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(G330), .B(new_n803), .C1(new_n906), .C2(new_n907), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n853), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1066), .A2(new_n1065), .A3(new_n802), .ZN(new_n1088));
  AOI21_X1  g0888(.A(KEYINPUT112), .B1(new_n1069), .B2(new_n801), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1087), .B(new_n1082), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n913), .B(G330), .C1(new_n907), .C2(new_n906), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n853), .A2(new_n1081), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n845), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1085), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n898), .A2(new_n899), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n855), .A2(new_n886), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1096), .A2(new_n1097), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1083), .B(new_n1095), .C1(new_n1098), .C2(new_n1091), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT113), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1091), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1104), .A2(KEYINPUT113), .A3(new_n1083), .A4(new_n1095), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1104), .A2(new_n1083), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1106), .B(new_n673), .C1(new_n1107), .C2(new_n1095), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n728), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1096), .A2(new_n733), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n729), .B1(new_n809), .B2(new_n318), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n748), .A2(G77), .B1(G283), .B2(new_n769), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1112), .A2(new_n274), .A3(new_n761), .A4(new_n819), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G97), .A2(new_n777), .B1(new_n745), .B2(G294), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n513), .B2(new_n765), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1113), .B(new_n1115), .C1(G107), .C2(new_n755), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT115), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G132), .A2(new_n812), .B1(new_n745), .B2(G125), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1118), .B1(new_n766), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(G128), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n989), .A2(new_n1121), .B1(new_n747), .B2(new_n742), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n759), .A2(new_n1019), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT53), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n274), .B1(G50), .B2(new_n818), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n1126), .A2(KEYINPUT114), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1126), .A2(KEYINPUT114), .B1(new_n755), .B2(G137), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1117), .A2(new_n1129), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1130), .A2(KEYINPUT116), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n738), .B1(new_n1130), .B2(KEYINPUT116), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1111), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1110), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1108), .A2(new_n1109), .A3(new_n1134), .ZN(G378));
  INV_X1    g0935(.A(KEYINPUT119), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n610), .A2(new_n609), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n322), .A2(new_n873), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1137), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n368), .B2(new_n325), .ZN(new_n1141));
  OR3_X1    g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1139), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n918), .B2(new_n650), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n914), .A2(new_n1144), .A3(new_n917), .A4(G330), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1146), .A2(new_n901), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n901), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1085), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n1106), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1136), .B1(new_n1152), .B2(KEYINPUT57), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1003), .B1(new_n1152), .B2(KEYINPUT57), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT57), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1085), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1156));
  OAI211_X1 g0956(.A(KEYINPUT119), .B(new_n1155), .C1(new_n1156), .C2(new_n1150), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1153), .A2(new_n1154), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1150), .A2(new_n727), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1145), .A2(new_n733), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1121), .A2(new_n765), .B1(new_n759), .B2(new_n1119), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G137), .B2(new_n777), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n748), .A2(G150), .B1(G125), .B2(new_n769), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n754), .C2(new_n816), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(G33), .A2(G41), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT117), .ZN(new_n1168));
  INV_X1    g0968(.A(G124), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n762), .A2(new_n742), .B1(new_n741), .B2(new_n1169), .ZN(new_n1170));
  NOR4_X1   g0970(.A1(new_n1165), .A2(new_n1166), .A3(new_n1168), .A4(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n747), .A2(new_n221), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n383), .B(new_n248), .C1(new_n759), .C2(new_n202), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(G116), .C2(new_n769), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n755), .A2(G97), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G58), .A2(new_n818), .B1(new_n745), .B2(G283), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n812), .A2(G107), .B1(new_n777), .B2(new_n498), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT58), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1168), .B(new_n327), .C1(new_n410), .C2(new_n466), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n793), .B1(new_n1171), .B2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT118), .Z(new_n1185));
  AOI211_X1 g0985(.A(new_n730), .B(new_n1185), .C1(new_n327), .C2(new_n808), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1159), .B1(new_n1160), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1158), .A2(new_n1187), .ZN(G375));
  INV_X1    g0988(.A(new_n1095), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n952), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1090), .A2(new_n1094), .A3(new_n1085), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n754), .A2(new_n513), .B1(new_n227), .B2(new_n766), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1193), .A2(KEYINPUT120), .B1(G294), .B2(new_n769), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(KEYINPUT120), .B2(new_n1193), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT121), .Z(new_n1196));
  AOI22_X1  g0996(.A1(G283), .A2(new_n812), .B1(new_n745), .B2(G303), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n202), .B2(new_n762), .C1(new_n226), .C2(new_n759), .ZN(new_n1198));
  NOR4_X1   g0998(.A1(new_n1196), .A2(new_n277), .A3(new_n1022), .A4(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n812), .A2(G137), .B1(G132), .B2(new_n769), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n754), .B2(new_n1119), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1202), .A2(KEYINPUT122), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n766), .A2(new_n316), .B1(new_n741), .B2(new_n1121), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n410), .B1(new_n747), .B2(new_n327), .C1(new_n394), .C2(new_n762), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(G159), .C2(new_n760), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1202), .A2(KEYINPUT122), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1203), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n793), .B1(new_n1199), .B2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1209), .B(new_n729), .C1(G68), .C2(new_n809), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n853), .B2(new_n733), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n728), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1192), .A2(new_n1213), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT123), .Z(G381));
  NOR2_X1   g1015(.A1(G375), .A2(G378), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n972), .A2(new_n1063), .A3(new_n1001), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1006), .A2(new_n797), .A3(new_n1038), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(new_n1217), .A2(G381), .A3(G384), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1216), .A2(new_n1219), .ZN(G407));
  NAND2_X1  g1020(.A1(new_n655), .A2(G213), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1216), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(G407), .A2(new_n1223), .A3(G213), .ZN(G409));
  NAND3_X1  g1024(.A1(new_n1158), .A2(G378), .A3(new_n1187), .ZN(new_n1225));
  INV_X1    g1025(.A(G378), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1187), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1156), .A2(new_n952), .A3(new_n1150), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1226), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1222), .B1(new_n1225), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1189), .A2(KEYINPUT60), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(KEYINPUT124), .A3(new_n1191), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT60), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1232), .B(new_n673), .C1(new_n1233), .C2(new_n1191), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT124), .B1(new_n1231), .B2(new_n1191), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1213), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT125), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G384), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n806), .A2(KEYINPUT125), .A3(new_n833), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1236), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1213), .B(new_n1239), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1230), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT63), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1218), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n797), .B1(new_n1006), .B2(new_n1038), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1217), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1063), .B1(new_n972), .B2(new_n1001), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1250), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G387), .A2(G390), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1250), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1217), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1253), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT126), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1258), .B(new_n1259), .ZN(new_n1260));
  AND4_X1   g1060(.A1(G2897), .A2(new_n1241), .A3(new_n1222), .A4(new_n1242), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1241), .A2(new_n1242), .B1(G2897), .B2(new_n1222), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1230), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1230), .A2(KEYINPUT63), .A3(new_n1244), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1247), .A2(new_n1260), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT62), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1230), .A2(new_n1267), .A3(new_n1244), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1257), .B1(new_n1230), .B2(new_n1263), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1267), .B1(new_n1230), .B2(new_n1244), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1253), .A2(new_n1256), .A3(KEYINPUT127), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT127), .B1(new_n1253), .B2(new_n1256), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1266), .B1(new_n1271), .B2(new_n1275), .ZN(G405));
  OAI21_X1  g1076(.A(new_n1244), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1274), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(new_n1272), .A3(new_n1243), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G375), .A2(new_n1226), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1225), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1280), .B(new_n1282), .ZN(G402));
endmodule


