//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n449, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n552, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1146, new_n1147, new_n1148;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT67), .Z(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT68), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT69), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  OR4_X1    g031(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n456), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XOR2_X1   g038(.A(KEYINPUT3), .B(G2104), .Z(new_n464));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT70), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n469), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  OR2_X1    g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND3_X1   g047(.A1(KEYINPUT71), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(KEYINPUT3), .B1(KEYINPUT71), .B2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n471), .A2(G2104), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n476), .A2(G137), .B1(G101), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(new_n471), .B2(G112), .ZN(new_n483));
  OAI22_X1  g058(.A1(new_n475), .A2(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n484), .B1(G124), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT72), .Z(G162));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G114), .C2(new_n471), .ZN(new_n490));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  XOR2_X1   g067(.A(new_n492), .B(KEYINPUT73), .Z(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n469), .A2(new_n494), .A3(G138), .A4(new_n471), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n475), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT74), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n509), .A2(new_n515), .ZN(G166));
  AND2_X1   g091(.A1(new_n510), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G51), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n506), .A2(new_n510), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT75), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n520), .A2(new_n522), .A3(new_n525), .ZN(G168));
  AOI22_X1  g101(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(new_n508), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n521), .A2(G90), .B1(new_n517), .B2(G52), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n527), .A2(new_n508), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n511), .A2(new_n533), .B1(new_n513), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g110(.A(KEYINPUT76), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n531), .A2(new_n536), .ZN(G171));
  AND2_X1   g112(.A1(G68), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(new_n506), .B2(G56), .ZN(new_n539));
  OR3_X1    g114(.A1(new_n539), .A2(KEYINPUT77), .A3(new_n508), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n521), .A2(G81), .B1(new_n517), .B2(G43), .ZN(new_n541));
  OAI21_X1  g116(.A(KEYINPUT77), .B1(new_n539), .B2(new_n508), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT78), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT78), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n540), .A2(new_n541), .A3(new_n545), .A4(new_n542), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(new_n548));
  XOR2_X1   g123(.A(new_n548), .B(KEYINPUT79), .Z(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT80), .ZN(G188));
  INV_X1    g130(.A(KEYINPUT81), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n504), .A2(KEYINPUT5), .A3(G543), .ZN(new_n557));
  AOI21_X1  g132(.A(KEYINPUT5), .B1(new_n504), .B2(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n503), .A2(KEYINPUT81), .A3(new_n505), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n559), .A2(G65), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT82), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT82), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n561), .A2(new_n565), .A3(new_n562), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(G651), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n517), .A2(new_n568), .A3(G53), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT9), .B1(new_n513), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n569), .A2(new_n571), .B1(G91), .B2(new_n521), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n567), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  NAND3_X1  g149(.A1(new_n520), .A2(new_n522), .A3(new_n525), .ZN(G286));
  INV_X1    g150(.A(G166), .ZN(G303));
  NAND2_X1  g151(.A1(new_n521), .A2(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n517), .A2(G49), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  AOI22_X1  g155(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n508), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n511), .A2(new_n583), .B1(new_n513), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n508), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n511), .A2(new_n590), .B1(new_n513), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G290));
  NAND3_X1  g169(.A1(new_n559), .A2(G66), .A3(new_n560), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G651), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n506), .A2(G92), .A3(new_n510), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n517), .A2(G54), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n604), .B2(G171), .ZN(G284));
  OAI21_X1  g181(.A(new_n605), .B1(new_n604), .B2(G171), .ZN(G321));
  NAND2_X1  g182(.A1(G299), .A2(new_n604), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n604), .B2(G168), .ZN(G297));
  XOR2_X1   g184(.A(G297), .B(KEYINPUT83), .Z(G280));
  XNOR2_X1  g185(.A(new_n599), .B(KEYINPUT10), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n508), .B1(new_n595), .B2(new_n596), .ZN(new_n612));
  INV_X1    g187(.A(new_n602), .ZN(new_n613));
  NOR3_X1   g188(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  OAI21_X1  g191(.A(G868), .B1(new_n603), .B2(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n547), .B2(G868), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n476), .A2(G135), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n620), .A2(KEYINPUT84), .B1(G123), .B2(new_n486), .ZN(new_n621));
  NOR2_X1   g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(new_n471), .B2(G111), .ZN(new_n623));
  OAI221_X1 g198(.A(new_n621), .B1(KEYINPUT84), .B2(new_n620), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT85), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n469), .A2(new_n477), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G2100), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(G2100), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n629), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT86), .Z(G156));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n640), .B(new_n641), .Z(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2435), .ZN(new_n644));
  XOR2_X1   g219(.A(G2427), .B(G2438), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n642), .B(new_n647), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n648), .A2(G14), .ZN(G401));
  XOR2_X1   g224(.A(G2067), .B(G2678), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n653), .B(KEYINPUT88), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT17), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n658), .A2(new_n652), .A3(new_n650), .ZN(new_n659));
  INV_X1    g234(.A(new_n652), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n658), .B2(new_n650), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n651), .A2(new_n653), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n656), .B(new_n659), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2096), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT89), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2100), .ZN(G227));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT20), .Z(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  INV_X1    g249(.A(new_n671), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n674), .B1(new_n668), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n668), .A2(KEYINPUT90), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n686), .A2(G27), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n499), .B2(G29), .ZN(new_n688));
  MUX2_X1   g263(.A(new_n687), .B(new_n688), .S(KEYINPUT102), .Z(new_n689));
  INV_X1    g264(.A(G2078), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT31), .B(G11), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT98), .B(G28), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(G29), .B1(new_n694), .B2(KEYINPUT30), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT99), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(KEYINPUT30), .B2(new_n694), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n692), .B(new_n697), .C1(new_n628), .C2(new_n686), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT100), .ZN(new_n699));
  MUX2_X1   g274(.A(G5), .B(G301), .S(G16), .Z(new_n700));
  MUX2_X1   g275(.A(G21), .B(G286), .S(G16), .Z(new_n701));
  AOI22_X1  g276(.A1(new_n700), .A2(G1961), .B1(G1966), .B2(new_n701), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n699), .B(new_n702), .C1(G1966), .C2(new_n701), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT101), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n486), .A2(G128), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n476), .A2(G140), .ZN(new_n706));
  NOR2_X1   g281(.A1(G104), .A2(G2105), .ZN(new_n707));
  OAI21_X1  g282(.A(G2104), .B1(new_n471), .B2(G116), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n705), .B(new_n706), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G29), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT95), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n686), .A2(G26), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G2067), .ZN(new_n715));
  OR2_X1    g290(.A1(KEYINPUT24), .A2(G34), .ZN(new_n716));
  NAND2_X1  g291(.A1(KEYINPUT24), .A2(G34), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n716), .A2(new_n686), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G160), .B2(new_n686), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n719), .A2(G2084), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n486), .A2(G129), .B1(G105), .B2(new_n477), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT26), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n476), .A2(G141), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT96), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G29), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G29), .B2(G32), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT27), .B(G1996), .ZN(new_n729));
  OAI22_X1  g304(.A1(new_n728), .A2(new_n729), .B1(new_n700), .B2(G1961), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n715), .A2(new_n720), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G4), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(G16), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n603), .B2(G16), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT94), .B(G1348), .Z(new_n735));
  XOR2_X1   g310(.A(new_n734), .B(new_n735), .Z(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT91), .B(G16), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(G19), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n547), .B2(new_n737), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(G1341), .Z(new_n740));
  NAND2_X1  g315(.A1(G299), .A2(G16), .ZN(new_n741));
  INV_X1    g316(.A(new_n737), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n742), .A2(KEYINPUT23), .A3(G20), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT23), .ZN(new_n744));
  INV_X1    g319(.A(G20), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n737), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n741), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G1956), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n731), .A2(new_n736), .A3(new_n740), .A4(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G29), .A2(G35), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G162), .B2(G29), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT29), .Z(new_n753));
  INV_X1    g328(.A(G2090), .ZN(new_n754));
  OAI22_X1  g329(.A1(new_n753), .A2(new_n754), .B1(new_n690), .B2(new_n689), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n754), .B2(new_n753), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n476), .A2(G139), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n477), .A2(G103), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT25), .Z(new_n759));
  AOI22_X1  g334(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n757), .B(new_n759), .C1(new_n760), .C2(new_n471), .ZN(new_n761));
  MUX2_X1   g336(.A(G33), .B(new_n761), .S(G29), .Z(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G2072), .Z(new_n763));
  AOI22_X1  g338(.A1(new_n728), .A2(new_n729), .B1(new_n719), .B2(G2084), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT97), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n756), .A2(new_n766), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n704), .A2(new_n750), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n593), .A2(new_n742), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G24), .B2(new_n742), .ZN(new_n770));
  INV_X1    g345(.A(G1986), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n486), .A2(G119), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n476), .A2(G131), .ZN(new_n774));
  NOR2_X1   g349(.A1(G95), .A2(G2105), .ZN(new_n775));
  OAI21_X1  g350(.A(G2104), .B1(new_n471), .B2(G107), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n773), .B(new_n774), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  MUX2_X1   g352(.A(G25), .B(new_n777), .S(G29), .Z(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT35), .B(G1991), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(G166), .A2(new_n737), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G22), .B2(new_n737), .ZN(new_n782));
  INV_X1    g357(.A(G1971), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G23), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(G16), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G288), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT92), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT33), .B(G1976), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G6), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(G16), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G305), .B2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT32), .B(G1981), .Z(new_n794));
  AND2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI22_X1  g370(.A1(new_n782), .A2(new_n783), .B1(new_n793), .B2(new_n794), .ZN(new_n796));
  OR4_X1    g371(.A1(new_n784), .A2(new_n790), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  AOI211_X1 g372(.A(new_n772), .B(new_n780), .C1(new_n797), .C2(KEYINPUT34), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n770), .A2(new_n771), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n797), .A2(KEYINPUT34), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT93), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(KEYINPUT93), .ZN(new_n803));
  AND3_X1   g378(.A1(new_n802), .A2(KEYINPUT36), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(KEYINPUT36), .B1(new_n802), .B2(new_n803), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n691), .B(new_n768), .C1(new_n804), .C2(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  AOI22_X1  g382(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(new_n508), .ZN(new_n809));
  INV_X1    g384(.A(G93), .ZN(new_n810));
  INV_X1    g385(.A(G55), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n511), .A2(new_n810), .B1(new_n513), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G860), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT37), .Z(new_n816));
  NAND2_X1  g391(.A1(new_n614), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n547), .A2(new_n814), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n543), .A2(new_n813), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n818), .B(new_n821), .Z(new_n822));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(G860), .B1(new_n824), .B2(KEYINPUT103), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(KEYINPUT103), .B2(new_n824), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n822), .A2(new_n823), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n816), .B1(new_n826), .B2(new_n827), .ZN(G145));
  INV_X1    g403(.A(new_n631), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n726), .A2(new_n709), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n726), .A2(new_n709), .ZN(new_n831));
  INV_X1    g406(.A(new_n492), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n498), .A2(new_n832), .ZN(new_n833));
  OR3_X1    g408(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n830), .B2(new_n831), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n829), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n834), .A2(new_n829), .A3(new_n835), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n628), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(new_n471), .B2(G118), .ZN(new_n841));
  INV_X1    g416(.A(G106), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n471), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n486), .A2(G130), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT104), .Z(new_n845));
  AOI211_X1 g420(.A(new_n843), .B(new_n845), .C1(G142), .C2(new_n476), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n761), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n777), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n837), .A2(new_n628), .A3(new_n838), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n840), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n848), .B1(new_n840), .B2(new_n849), .ZN(new_n851));
  XNOR2_X1  g426(.A(G160), .B(G162), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OR3_X1    g428(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(G37), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n853), .B1(new_n850), .B2(new_n851), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g433(.A(G166), .B(G288), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n859), .A2(new_n586), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n586), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G290), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n860), .A2(new_n593), .A3(new_n861), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT42), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(KEYINPUT107), .B2(new_n866), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n867), .A2(KEYINPUT108), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(KEYINPUT108), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n866), .A2(KEYINPUT107), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n870), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n614), .A2(new_n615), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n821), .B(new_n874), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n561), .A2(new_n565), .A3(new_n562), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n565), .B1(new_n561), .B2(new_n562), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n876), .A2(new_n877), .A3(new_n508), .ZN(new_n878));
  INV_X1    g453(.A(new_n572), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n614), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n567), .A2(new_n603), .A3(new_n572), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n875), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(KEYINPUT41), .A3(new_n881), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n885), .A2(KEYINPUT106), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT106), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n880), .A2(new_n887), .A3(new_n881), .A4(KEYINPUT41), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n882), .B2(new_n891), .ZN(new_n892));
  AOI211_X1 g467(.A(KEYINPUT105), .B(KEYINPUT41), .C1(new_n880), .C2(new_n881), .ZN(new_n893));
  OAI22_X1  g468(.A1(new_n886), .A2(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n884), .B1(new_n875), .B2(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n873), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n873), .A2(new_n895), .ZN(new_n897));
  OAI21_X1  g472(.A(G868), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(G868), .B2(new_n813), .ZN(G295));
  OAI21_X1  g474(.A(new_n898), .B1(G868), .B2(new_n813), .ZN(G331));
  INV_X1    g475(.A(KEYINPUT111), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n902));
  NAND3_X1  g477(.A1(G286), .A2(new_n531), .A3(new_n536), .ZN(new_n903));
  NAND2_X1  g478(.A1(G171), .A2(G168), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n819), .A2(new_n820), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n903), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n813), .B1(new_n544), .B2(new_n546), .ZN(new_n907));
  INV_X1    g482(.A(new_n820), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n567), .A2(new_n603), .A3(new_n572), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n603), .B1(new_n567), .B2(new_n572), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n891), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT105), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n882), .A2(new_n890), .A3(new_n891), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n885), .A2(KEYINPUT106), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n888), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n910), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n883), .B1(new_n905), .B2(new_n909), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n902), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n910), .A2(new_n882), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n914), .A2(new_n915), .B1(new_n917), .B2(new_n888), .ZN(new_n923));
  OAI211_X1 g498(.A(KEYINPUT109), .B(new_n922), .C1(new_n923), .C2(new_n910), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n921), .A2(new_n865), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n863), .A2(new_n864), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n926), .B(new_n922), .C1(new_n923), .C2(new_n910), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT110), .ZN(new_n928));
  INV_X1    g503(.A(new_n910), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n894), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT110), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n930), .A2(new_n931), .A3(new_n926), .A4(new_n922), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n932), .A3(new_n855), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n901), .B(KEYINPUT43), .C1(new_n925), .C2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n921), .A2(new_n865), .A3(new_n924), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n936), .A2(new_n855), .A3(new_n928), .A4(new_n932), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n901), .B1(new_n937), .B2(KEYINPUT43), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n933), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n910), .B1(new_n885), .B2(new_n913), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n865), .B1(new_n942), .B2(new_n920), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT44), .B1(new_n939), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n937), .A2(new_n941), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n940), .A2(KEYINPUT43), .A3(new_n943), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT112), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT111), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(new_n944), .A3(new_n934), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n946), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n955));
  INV_X1    g530(.A(new_n949), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n950), .A2(new_n957), .ZN(G397));
  INV_X1    g533(.A(KEYINPUT119), .ZN(new_n959));
  XNOR2_X1  g534(.A(G299), .B(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT57), .ZN(new_n961));
  AOI21_X1  g536(.A(G1384), .B1(new_n498), .B2(new_n832), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT45), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G1384), .B1(new_n493), .B2(new_n498), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(KEYINPUT45), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n472), .A2(G40), .A3(new_n478), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(KEYINPUT56), .B(G2072), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n472), .A2(G40), .A3(new_n478), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n971), .B(new_n972), .C1(new_n970), .C2(new_n962), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n968), .A2(new_n969), .B1(new_n748), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n961), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(KEYINPUT120), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT120), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n961), .B2(new_n974), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n833), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n967), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(G2067), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT121), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n962), .A2(new_n970), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n986), .B(new_n972), .C1(new_n970), .C2(new_n965), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n984), .A2(new_n985), .B1(new_n735), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT121), .B1(new_n983), .B2(G2067), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n603), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n961), .A2(new_n974), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n979), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT123), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n975), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n961), .A2(new_n974), .A3(KEYINPUT123), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(KEYINPUT61), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT61), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n976), .B2(new_n978), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT60), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n988), .A2(new_n999), .A3(new_n614), .A4(new_n989), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n988), .A2(new_n603), .A3(new_n989), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT60), .B1(new_n1001), .B2(new_n990), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n996), .A2(new_n998), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n499), .A2(new_n980), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1006), .A2(new_n972), .A3(new_n963), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT58), .B(G1341), .Z(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI22_X1  g584(.A1(new_n1007), .A2(G1996), .B1(new_n982), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT122), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n547), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT59), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n992), .B1(new_n1003), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n981), .A2(new_n1005), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n965), .A2(KEYINPUT45), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n972), .ZN(new_n1020));
  OAI22_X1  g595(.A1(new_n1020), .A2(G1966), .B1(new_n987), .B2(G2084), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(G8), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1022), .B(new_n1023), .C1(new_n1024), .C2(G168), .ZN(new_n1025));
  OAI211_X1 g600(.A(KEYINPUT51), .B(G8), .C1(new_n1021), .C2(G286), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1021), .A2(G8), .A3(G286), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G303), .A2(G8), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT55), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(KEYINPUT117), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1007), .A2(KEYINPUT116), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1006), .A2(new_n1034), .A3(new_n972), .A4(new_n963), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1971), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n987), .A2(G2090), .ZN(new_n1037));
  OAI211_X1 g612(.A(G8), .B(new_n1032), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n982), .A2(new_n1024), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1976), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G288), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT52), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n586), .B(G1981), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1044), .A2(KEYINPUT49), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(KEYINPUT49), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1039), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(G288), .B2(new_n1041), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1039), .B(new_n1048), .C1(new_n1041), .C2(G288), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1043), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1036), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n973), .A2(G2090), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1024), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1031), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1038), .B(new_n1050), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1029), .A2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT124), .B(G1961), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n987), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1033), .A2(new_n690), .A3(new_n1035), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT125), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1018), .A2(new_n972), .A3(KEYINPUT53), .A4(new_n690), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1019), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1061), .A2(new_n1062), .A3(G301), .A4(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1063), .A2(new_n964), .ZN(new_n1067));
  AOI211_X1 g642(.A(new_n1067), .B(new_n1058), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT125), .B1(new_n1068), .B2(G301), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  OAI211_X1 g646(.A(KEYINPUT54), .B(new_n1066), .C1(new_n1069), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(G171), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1068), .A2(G301), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1017), .A2(new_n1056), .A3(new_n1077), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1079), .A2(new_n1050), .A3(G8), .A4(new_n1032), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT118), .B1(new_n1079), .B2(G8), .ZN(new_n1081));
  OAI211_X1 g656(.A(KEYINPUT118), .B(G8), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1031), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1038), .A2(new_n1050), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1022), .A2(G286), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1084), .A2(KEYINPUT63), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1055), .A2(G286), .A3(new_n1022), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(KEYINPUT63), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G288), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1047), .A2(new_n1041), .A3(new_n1090), .ZN(new_n1091));
  OR2_X1    g666(.A1(G305), .A2(G1981), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1040), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1095), .A2(new_n1055), .A3(new_n1073), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1029), .A2(new_n1094), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1093), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1078), .A2(new_n1080), .A3(new_n1089), .A4(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT113), .B1(new_n1018), .B2(new_n967), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT113), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n972), .A2(new_n1101), .A3(new_n1005), .A4(new_n981), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1100), .A2(KEYINPUT114), .A3(new_n1102), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n726), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1103), .A2(G1996), .ZN(new_n1108));
  OAI22_X1  g683(.A1(new_n1107), .A2(new_n1108), .B1(G1996), .B2(new_n726), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n709), .B(G2067), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1110), .A2(KEYINPUT115), .A3(new_n1111), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1109), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n777), .A2(new_n779), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n777), .A2(new_n779), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1110), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1103), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n593), .B(new_n771), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1099), .A2(new_n1120), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1110), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1109), .A2(new_n1114), .A3(new_n1117), .A4(new_n1115), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n709), .A2(G2067), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT127), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1110), .A2(new_n1111), .B1(KEYINPUT46), .B2(new_n1108), .ZN(new_n1132));
  OAI221_X1 g707(.A(new_n1132), .B1(KEYINPUT46), .B2(new_n1108), .C1(new_n726), .C2(new_n1125), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT47), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1121), .A2(new_n771), .A3(new_n593), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT48), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1120), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1130), .A2(new_n1131), .A3(new_n1134), .A4(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1139));
  AOI211_X1 g714(.A(KEYINPUT126), .B(new_n1125), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1137), .B(new_n1134), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT127), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1124), .A2(new_n1143), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g719(.A1(G227), .A2(G401), .ZN(new_n1146));
  AND2_X1   g720(.A1(new_n857), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g721(.A1(G229), .A2(new_n462), .ZN(new_n1148));
  AND3_X1   g722(.A1(new_n1147), .A2(new_n953), .A3(new_n1148), .ZN(G308));
  NAND3_X1  g723(.A1(new_n1147), .A2(new_n953), .A3(new_n1148), .ZN(G225));
endmodule


