//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202));
  NAND2_X1  g001(.A1(G229gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(KEYINPUT13), .Z(new_n204));
  INV_X1    g003(.A(G1gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT16), .ZN(new_n206));
  INV_X1    g005(.A(G15gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G22gat), .ZN(new_n208));
  INV_X1    g007(.A(G22gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G15gat), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n206), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(G1gat), .B1(new_n208), .B2(new_n210), .ZN(new_n212));
  OAI21_X1  g011(.A(G8gat), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n206), .A2(new_n208), .A3(new_n210), .ZN(new_n214));
  INV_X1    g013(.A(G8gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n214), .B(new_n215), .C1(G1gat), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G29gat), .ZN(new_n219));
  INV_X1    g018(.A(G36gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT14), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT14), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(G29gat), .A2(G36gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  INV_X1    g025(.A(G43gat), .ZN(new_n227));
  INV_X1    g026(.A(G50gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G43gat), .A2(G50gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT94), .ZN(new_n233));
  INV_X1    g032(.A(new_n230), .ZN(new_n234));
  NOR2_X1   g033(.A1(G43gat), .A2(G50gat), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT15), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n229), .A2(new_n226), .A3(new_n230), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n232), .B(new_n233), .C1(new_n238), .C2(new_n225), .ZN(new_n239));
  INV_X1    g038(.A(new_n225), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n240), .A2(KEYINPUT94), .A3(new_n236), .A4(new_n237), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n218), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n218), .B1(new_n239), .B2(new_n241), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n204), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT92), .B(KEYINPUT11), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G169gat), .ZN(new_n249));
  INV_X1    g048(.A(G197gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G169gat), .A2(G197gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT93), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT93), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(new_n255), .A3(new_n252), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n245), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n248), .A2(new_n254), .A3(new_n256), .A4(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n248), .A2(new_n258), .B1(new_n254), .B2(new_n256), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n258), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n254), .A2(new_n256), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT12), .B1(new_n266), .B2(new_n259), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n239), .A2(new_n241), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT17), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n239), .A2(KEYINPUT17), .A3(new_n241), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n218), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n218), .A2(new_n239), .A3(new_n241), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(KEYINPUT18), .A3(new_n203), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n244), .B(new_n268), .C1(new_n273), .C2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n218), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n239), .A2(KEYINPUT17), .A3(new_n241), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT17), .B1(new_n239), .B2(new_n241), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n274), .A2(new_n203), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT18), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n202), .B1(new_n276), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT18), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(new_n273), .B2(new_n281), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n261), .B1(new_n260), .B2(new_n262), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n266), .A2(KEYINPUT12), .A3(new_n259), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n269), .A2(new_n277), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n274), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n289), .B1(new_n291), .B2(new_n204), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n280), .A2(KEYINPUT18), .A3(new_n282), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n286), .A2(new_n292), .A3(new_n293), .A4(KEYINPUT95), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n284), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n244), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n289), .B1(new_n296), .B2(new_n283), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G211gat), .B(G218gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT22), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT75), .B(G211gat), .ZN(new_n303));
  INV_X1    g102(.A(G218gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n308));
  XNOR2_X1  g107(.A(G197gat), .B(G204gat), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n308), .B1(new_n307), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n301), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n307), .A2(new_n309), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT77), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n315), .A3(new_n300), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G155gat), .B(G162gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G141gat), .B(G148gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n319), .B1(KEYINPUT2), .B2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(KEYINPUT83), .B(KEYINPUT3), .Z(new_n322));
  XOR2_X1   g121(.A(G141gat), .B(G148gat), .Z(new_n323));
  INV_X1    g122(.A(KEYINPUT80), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(KEYINPUT80), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n318), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT81), .B(G155gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n328), .B1(new_n329), .B2(G162gat), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n321), .B(new_n322), .C1(new_n327), .C2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(G228gat), .A3(G233gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n321), .B1(new_n327), .B2(new_n330), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT82), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT82), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n338), .B(new_n321), .C1(new_n327), .C2(new_n330), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n312), .A2(new_n316), .A3(new_n332), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OR2_X1    g142(.A1(new_n335), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G228gat), .A2(G233gat), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n345), .B(KEYINPUT86), .Z(new_n346));
  INV_X1    g145(.A(new_n336), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n347), .B1(new_n341), .B2(new_n322), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n317), .A2(new_n333), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n346), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT87), .B1(new_n344), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT31), .B(G50gat), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n352), .B(new_n353), .Z(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(G22gat), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT87), .ZN(new_n357));
  INV_X1    g156(.A(new_n350), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n335), .A2(new_n343), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(new_n209), .A3(new_n354), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n358), .A2(new_n357), .A3(new_n359), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n356), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(new_n356), .B2(new_n361), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(KEYINPUT67), .B(G190gat), .Z(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT27), .B(G183gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(KEYINPUT28), .ZN(new_n369));
  NOR2_X1   g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n370), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n371));
  OR2_X1    g170(.A1(new_n370), .A2(KEYINPUT26), .ZN(new_n372));
  INV_X1    g171(.A(G176gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n249), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n371), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  OR2_X1    g174(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G183gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n366), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT24), .ZN(new_n380));
  INV_X1    g179(.A(G190gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n380), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT66), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(G169gat), .B2(G176gat), .ZN(new_n385));
  OR2_X1    g184(.A1(new_n385), .A2(KEYINPUT23), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n374), .B1(KEYINPUT23), .B2(new_n385), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n383), .A2(KEYINPUT25), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n379), .A2(KEYINPUT65), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n382), .B(new_n389), .C1(G183gat), .C2(G190gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n379), .A2(KEYINPUT65), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n386), .B(new_n387), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G226gat), .A2(G233gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n332), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n388), .A2(new_n394), .A3(KEYINPUT68), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT68), .B1(new_n388), .B2(new_n394), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n376), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n398), .B1(new_n402), .B2(new_n397), .ZN(new_n403));
  INV_X1    g202(.A(new_n317), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT79), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT79), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n369), .A2(new_n375), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT68), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n413), .B2(new_n399), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n397), .B1(new_n414), .B2(KEYINPUT29), .ZN(new_n415));
  INV_X1    g214(.A(new_n397), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n410), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n402), .B2(new_n332), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(KEYINPUT78), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n317), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n409), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  OR3_X1    g225(.A1(new_n422), .A2(KEYINPUT30), .A3(new_n426), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n403), .A2(KEYINPUT79), .A3(new_n404), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT79), .B1(new_n403), .B2(new_n404), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n417), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT78), .B1(new_n419), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n410), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n404), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n426), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n409), .A2(new_n421), .A3(new_n425), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT30), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n427), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT4), .ZN(new_n439));
  XOR2_X1   g238(.A(G113gat), .B(G120gat), .Z(new_n440));
  INV_X1    g239(.A(KEYINPUT1), .ZN(new_n441));
  XNOR2_X1  g240(.A(G127gat), .B(G134gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n441), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT69), .B(G134gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G127gat), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(KEYINPUT70), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G134gat), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT70), .B1(new_n448), .B2(G127gat), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n445), .B2(G127gat), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n443), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT84), .B1(new_n451), .B2(new_n336), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n451), .A2(new_n336), .A3(KEYINPUT84), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n439), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(G225gat), .A2(G233gat), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n337), .A2(KEYINPUT3), .A3(new_n339), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n331), .A2(new_n451), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n451), .A2(KEYINPUT71), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT71), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n462), .B(new_n443), .C1(new_n447), .C2(new_n450), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n461), .A2(KEYINPUT4), .A3(new_n347), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n455), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT5), .ZN(new_n466));
  INV_X1    g265(.A(new_n451), .ZN(new_n467));
  OAI22_X1  g266(.A1(new_n453), .A2(new_n454), .B1(new_n340), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n466), .B1(new_n468), .B2(new_n457), .ZN(new_n469));
  OR3_X1    g268(.A1(new_n451), .A2(new_n336), .A3(KEYINPUT84), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(KEYINPUT4), .A3(new_n452), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n461), .A2(new_n463), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n439), .B1(new_n472), .B2(new_n336), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n460), .A2(new_n466), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n465), .A2(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  XOR2_X1   g275(.A(G1gat), .B(G29gat), .Z(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G57gat), .B(G85gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT6), .B1(new_n476), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n469), .A2(new_n465), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n474), .A2(new_n475), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n481), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(KEYINPUT6), .A3(new_n481), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n438), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n450), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n493), .B(new_n444), .C1(KEYINPUT70), .C2(new_n446), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n462), .B1(new_n494), .B2(new_n443), .ZN(new_n495));
  INV_X1    g294(.A(new_n463), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT72), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT72), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n461), .A2(new_n498), .A3(new_n463), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n402), .ZN(new_n501));
  NAND2_X1  g300(.A1(G227gat), .A2(G233gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT64), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n414), .A2(new_n497), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n501), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT34), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT74), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G43gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(G71gat), .B(G99gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n413), .A2(new_n399), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n513), .A2(new_n376), .B1(new_n497), .B2(new_n499), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n513), .A2(new_n497), .A3(new_n376), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n503), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT33), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n512), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n504), .B1(new_n501), .B2(new_n505), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT32), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT73), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT73), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n516), .A2(new_n522), .A3(KEYINPUT32), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n518), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n516), .B(KEYINPUT32), .C1(new_n517), .C2(new_n512), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n507), .A2(KEYINPUT74), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n527), .B1(new_n524), .B2(new_n525), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n509), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n524), .A2(new_n525), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n526), .ZN(new_n532));
  INV_X1    g331(.A(new_n509), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n524), .A2(new_n527), .A3(new_n525), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n365), .A2(new_n492), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT35), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT39), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n458), .A2(new_n459), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n471), .A2(new_n473), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(KEYINPUT88), .A3(new_n457), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT88), .B1(new_n541), .B2(new_n457), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n539), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n544), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n468), .A2(new_n457), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(new_n539), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(new_n542), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n545), .A2(new_n549), .A3(new_n482), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT40), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n550), .A2(new_n551), .B1(new_n481), .B2(new_n486), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(new_n427), .A3(new_n437), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n545), .A2(new_n549), .A3(KEYINPUT40), .A4(new_n482), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT89), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT90), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n427), .A2(new_n437), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT89), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n554), .B(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT90), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n557), .A2(new_n559), .A3(new_n560), .A4(new_n552), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n426), .A2(KEYINPUT37), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n435), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n404), .B1(new_n418), .B2(new_n420), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n403), .A2(new_n317), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(KEYINPUT37), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n564), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n488), .A2(new_n489), .A3(new_n436), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n435), .A2(new_n563), .B1(new_n422), .B2(KEYINPUT37), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n565), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n356), .A2(new_n361), .A3(new_n362), .ZN(new_n573));
  INV_X1    g372(.A(new_n364), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n562), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n530), .A2(new_n535), .A3(KEYINPUT36), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT36), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n536), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n574), .A2(new_n573), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n491), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n576), .A2(new_n577), .A3(new_n579), .A4(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n299), .B1(new_n538), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G71gat), .ZN(new_n586));
  INV_X1    g385(.A(G78gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT9), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n585), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n589), .B(new_n588), .C1(new_n584), .C2(new_n591), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n218), .B1(new_n596), .B2(KEYINPUT21), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT97), .ZN(new_n598));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT96), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n598), .A2(new_n602), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n595), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G127gat), .B(G155gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  XOR2_X1   g410(.A(new_n605), .B(new_n611), .Z(new_n612));
  NAND2_X1  g411(.A1(G85gat), .A2(G92gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT7), .ZN(new_n614));
  XNOR2_X1  g413(.A(G99gat), .B(G106gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(G99gat), .A2(G106gat), .ZN(new_n616));
  INV_X1    g415(.A(G85gat), .ZN(new_n617));
  INV_X1    g416(.A(G92gat), .ZN(new_n618));
  AOI22_X1  g417(.A1(KEYINPUT8), .A2(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n614), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n615), .B1(new_n614), .B2(new_n619), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n269), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n622), .B1(KEYINPUT41), .B2(new_n623), .ZN(new_n624));
  OAI22_X1  g423(.A1(new_n278), .A2(new_n279), .B1(new_n620), .B2(new_n621), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G190gat), .B(G218gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT98), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n632));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n629), .A2(new_n634), .A3(new_n630), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n612), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n614), .A2(new_n619), .ZN(new_n640));
  INV_X1    g439(.A(new_n615), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n614), .A2(new_n615), .A3(new_n619), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n642), .A2(new_n594), .A3(new_n593), .A4(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n595), .B1(new_n620), .B2(new_n621), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n596), .A2(KEYINPUT10), .A3(new_n643), .A4(new_n642), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n644), .A2(new_n645), .ZN(new_n652));
  INV_X1    g451(.A(new_n650), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  NAND3_X1  g456(.A1(new_n651), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT99), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n651), .A2(new_n654), .A3(new_n660), .A4(new_n657), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n651), .A2(new_n654), .ZN(new_n663));
  INV_X1    g462(.A(new_n657), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(KEYINPUT100), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT100), .B1(new_n663), .B2(new_n664), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n639), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n583), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n490), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(new_n205), .ZN(G1324gat));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n670), .A2(new_n438), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT16), .B(G8gat), .Z(new_n675));
  AOI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G8gat), .B1(new_n670), .B2(new_n438), .ZN(new_n677));
  NOR2_X1   g476(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n678));
  MUX2_X1   g477(.A(KEYINPUT101), .B(new_n678), .S(new_n675), .Z(new_n679));
  AOI22_X1  g478(.A1(new_n676), .A2(new_n677), .B1(new_n674), .B2(new_n679), .ZN(G1325gat));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n530), .A2(new_n535), .A3(KEYINPUT36), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT36), .B1(new_n530), .B2(new_n535), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n579), .A2(KEYINPUT102), .A3(new_n577), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G15gat), .B1(new_n670), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n536), .A2(new_n207), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n688), .B1(new_n670), .B2(new_n689), .ZN(G1326gat));
  NOR2_X1   g489(.A1(new_n670), .A2(new_n365), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  INV_X1    g492(.A(new_n612), .ZN(new_n694));
  INV_X1    g493(.A(new_n668), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n638), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n583), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n490), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n219), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT45), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n636), .A2(new_n637), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n702), .A2(KEYINPUT44), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT35), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n537), .B(new_n704), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n579), .B(new_n577), .C1(new_n365), .C2(new_n492), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n562), .B2(new_n575), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n703), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n298), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n295), .A2(KEYINPUT103), .A3(new_n297), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n365), .B2(new_n492), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n580), .A2(KEYINPUT104), .A3(new_n491), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n717), .A2(new_n576), .A3(new_n685), .A4(new_n684), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n638), .B1(new_n718), .B2(new_n538), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n708), .B(new_n713), .C1(new_n719), .C2(KEYINPUT44), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(KEYINPUT105), .A3(new_n490), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT105), .B1(new_n720), .B2(new_n490), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G29gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n701), .B1(new_n721), .B2(new_n723), .ZN(G1328gat));
  NAND3_X1  g523(.A1(new_n698), .A2(new_n220), .A3(new_n557), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT46), .Z(new_n726));
  OAI21_X1  g525(.A(G36gat), .B1(new_n720), .B2(new_n438), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1329gat));
  INV_X1    g527(.A(new_n536), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(G43gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n583), .A2(new_n697), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G43gat), .B1(new_n720), .B2(new_n687), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(KEYINPUT47), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n733), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n734), .A2(new_n735), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n734), .A2(new_n731), .A3(new_n736), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n737), .A2(new_n738), .B1(new_n739), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g539(.A(G50gat), .B1(new_n720), .B2(new_n365), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n365), .A2(G50gat), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n698), .A2(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n743), .A2(new_n744), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n746), .B(new_n748), .ZN(G1331gat));
  NAND2_X1  g548(.A1(new_n718), .A2(new_n538), .ZN(new_n750));
  INV_X1    g549(.A(new_n712), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n751), .A2(new_n639), .A3(new_n695), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n490), .B(KEYINPUT109), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT110), .B(G57gat), .Z(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1332gat));
  NOR2_X1   g557(.A1(new_n753), .A2(new_n438), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  AND2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n759), .B2(new_n760), .ZN(G1333gat));
  OAI21_X1  g562(.A(G71gat), .B1(new_n753), .B2(new_n687), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n536), .A2(new_n586), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n753), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g566(.A1(new_n753), .A2(new_n365), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(new_n587), .ZN(G1335gat));
  NOR2_X1   g568(.A1(new_n751), .A2(new_n612), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n719), .A2(KEYINPUT51), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT51), .B1(new_n719), .B2(new_n770), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n773), .A2(new_n617), .A3(new_n699), .A4(new_n668), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n770), .A2(new_n668), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n708), .B(new_n776), .C1(new_n719), .C2(KEYINPUT44), .ZN(new_n777));
  OAI21_X1  g576(.A(G85gat), .B1(new_n777), .B2(new_n490), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n774), .A2(new_n778), .ZN(G1336gat));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  OAI21_X1  g579(.A(G92gat), .B1(new_n777), .B2(new_n438), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n438), .A2(new_n695), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n618), .B(new_n784), .C1(new_n771), .C2(new_n772), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n781), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n785), .B(new_n781), .C1(new_n782), .C2(new_n780), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(G1337gat));
  NOR3_X1   g588(.A1(new_n729), .A2(G99gat), .A3(new_n695), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G99gat), .B1(new_n777), .B2(new_n687), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(G1338gat));
  NOR3_X1   g592(.A1(new_n365), .A2(G106gat), .A3(new_n695), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n771), .B2(new_n772), .ZN(new_n795));
  OAI21_X1  g594(.A(G106gat), .B1(new_n777), .B2(new_n365), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(KEYINPUT112), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n795), .B(new_n796), .C1(KEYINPUT112), .C2(KEYINPUT53), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(G1339gat));
  AND3_X1   g601(.A1(new_n295), .A2(KEYINPUT103), .A3(new_n297), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT103), .B1(new_n295), .B2(new_n297), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n647), .A2(new_n648), .A3(new_n653), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n651), .A2(KEYINPUT54), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n653), .B1(new_n647), .B2(new_n648), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n657), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n806), .A2(KEYINPUT55), .A3(new_n809), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n662), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n803), .A2(new_n804), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n203), .B1(new_n280), .B2(new_n274), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n291), .A2(new_n204), .ZN(new_n817));
  OAI22_X1  g616(.A1(new_n816), .A2(new_n817), .B1(new_n260), .B2(new_n262), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n295), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(new_n668), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n638), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n662), .A2(new_n812), .A3(new_n813), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n702), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n612), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n751), .A2(new_n639), .A3(new_n668), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT113), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n710), .A2(new_n822), .A3(new_n711), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n819), .A2(new_n668), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n702), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n819), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n638), .A2(new_n830), .A3(new_n814), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n694), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n669), .A2(new_n712), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AND4_X1   g634(.A1(new_n438), .A2(new_n826), .A3(new_n755), .A4(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n580), .A2(new_n729), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(G113gat), .B1(new_n838), .B2(new_n751), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n826), .A2(new_n835), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n580), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n557), .A2(new_n490), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n536), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT114), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n298), .A2(G113gat), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n839), .B1(new_n845), .B2(new_n846), .ZN(G1340gat));
  AOI21_X1  g646(.A(G120gat), .B1(new_n838), .B2(new_n668), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n668), .A2(G120gat), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n845), .B2(new_n849), .ZN(G1341gat));
  OAI21_X1  g649(.A(G127gat), .B1(new_n844), .B2(new_n694), .ZN(new_n851));
  INV_X1    g650(.A(G127gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n838), .A2(new_n852), .A3(new_n612), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(G1342gat));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n445), .A3(new_n702), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT56), .Z(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n844), .B2(new_n638), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n856), .A2(KEYINPUT115), .A3(new_n857), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1343gat));
  NOR2_X1   g661(.A1(new_n686), .A2(new_n365), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n836), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(G141gat), .A3(new_n299), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867));
  INV_X1    g666(.A(G141gat), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT57), .B1(new_n363), .B2(new_n364), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n299), .A2(new_n814), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n638), .B1(new_n820), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n823), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n825), .B1(new_n872), .B2(new_n694), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n826), .A2(new_n580), .A3(new_n835), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n684), .A2(new_n685), .A3(new_n842), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n877), .A2(new_n878), .A3(new_n299), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n866), .B(new_n867), .C1(new_n868), .C2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n875), .A2(new_n876), .ZN(new_n882));
  INV_X1    g681(.A(new_n874), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n684), .A2(new_n685), .A3(new_n842), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(KEYINPUT116), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n877), .B2(new_n878), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n886), .A2(new_n751), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(G141gat), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n865), .B1(new_n890), .B2(KEYINPUT117), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n889), .A2(new_n892), .A3(G141gat), .ZN(new_n893));
  AOI211_X1 g692(.A(new_n881), .B(new_n867), .C1(new_n891), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n890), .A2(KEYINPUT117), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n893), .A3(new_n866), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT118), .B1(new_n896), .B2(KEYINPUT58), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n880), .B1(new_n894), .B2(new_n897), .ZN(G1344gat));
  AND2_X1   g697(.A1(new_n886), .A2(new_n888), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n668), .ZN(new_n900));
  INV_X1    g699(.A(G148gat), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(KEYINPUT59), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n872), .A2(new_n694), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n669), .A2(new_n299), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT57), .B1(new_n905), .B2(new_n580), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n840), .A2(new_n869), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n885), .A2(new_n668), .ZN(new_n911));
  OAI21_X1  g710(.A(G148gat), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n900), .A2(new_n902), .B1(new_n912), .B2(KEYINPUT59), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n864), .A2(G148gat), .A3(new_n695), .ZN(new_n914));
  OR3_X1    g713(.A1(new_n913), .A2(KEYINPUT120), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT120), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1345gat));
  INV_X1    g716(.A(new_n329), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n918), .B1(new_n899), .B2(new_n612), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n864), .A2(new_n329), .A3(new_n694), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n919), .A2(new_n920), .ZN(G1346gat));
  NAND3_X1  g720(.A1(new_n899), .A2(G162gat), .A3(new_n702), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n864), .A2(new_n638), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(G162gat), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT121), .ZN(G1347gat));
  NOR3_X1   g724(.A1(new_n729), .A2(new_n438), .A3(new_n755), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n841), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n299), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT122), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n840), .A2(new_n699), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n837), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n931), .A2(new_n438), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n249), .A3(new_n751), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n929), .A2(new_n933), .ZN(G1348gat));
  OAI21_X1  g733(.A(G176gat), .B1(new_n927), .B2(new_n695), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n784), .A2(new_n373), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n931), .B2(new_n936), .ZN(G1349gat));
  NAND3_X1  g736(.A1(new_n932), .A2(new_n367), .A3(new_n612), .ZN(new_n938));
  OAI21_X1  g737(.A(G183gat), .B1(new_n927), .B2(new_n694), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n940));
  AOI22_X1  g739(.A1(new_n938), .A2(new_n939), .B1(KEYINPUT123), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n940), .A2(KEYINPUT123), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n941), .B(new_n942), .ZN(G1350gat));
  NAND3_X1  g742(.A1(new_n932), .A2(new_n366), .A3(new_n702), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT124), .ZN(new_n945));
  OAI21_X1  g744(.A(G190gat), .B1(new_n927), .B2(new_n638), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1351gat));
  AND2_X1   g747(.A1(new_n863), .A2(new_n930), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n949), .A2(new_n557), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n250), .A3(new_n751), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952));
  INV_X1    g751(.A(new_n910), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n686), .A2(new_n438), .A3(new_n755), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n952), .B1(new_n955), .B2(new_n299), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G197gat), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n955), .A2(new_n952), .A3(new_n299), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n951), .B1(new_n957), .B2(new_n958), .ZN(G1352gat));
  INV_X1    g758(.A(G204gat), .ZN(new_n960));
  INV_X1    g759(.A(new_n955), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(new_n668), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n949), .A2(new_n960), .A3(new_n784), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT126), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n963), .B(new_n967), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n968), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT127), .B1(new_n968), .B2(KEYINPUT62), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(G1353gat));
  NAND3_X1  g770(.A1(new_n950), .A2(new_n303), .A3(new_n612), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n961), .A2(new_n612), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(G1354gat));
  OAI21_X1  g775(.A(G218gat), .B1(new_n955), .B2(new_n638), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n950), .A2(new_n304), .A3(new_n702), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(G1355gat));
endmodule


