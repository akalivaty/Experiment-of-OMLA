//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n565, new_n567,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT66), .Z(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(KEYINPUT68), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(new_n463), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(G137), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT67), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n463), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n466), .A2(new_n474), .A3(G125), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n471), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n463), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n480), .B1(new_n461), .B2(new_n464), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n481), .A2(new_n471), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n484), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND3_X1  g066(.A1(new_n465), .A2(G126), .A3(new_n466), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n471), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n471), .A2(G102), .A3(G2104), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n466), .A2(new_n474), .A3(G138), .A4(new_n471), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT4), .A2(G138), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n465), .A2(new_n471), .A3(new_n466), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n494), .A2(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(G50), .A3(G543), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n510), .B(new_n512), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G88), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n510), .A2(new_n512), .A3(G62), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(KEYINPUT69), .B1(new_n520), .B2(G651), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n522));
  AOI211_X1 g097(.A(new_n522), .B(new_n504), .C1(new_n518), .C2(new_n519), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n508), .B(new_n517), .C1(new_n521), .C2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(new_n516), .A2(G89), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT74), .B(KEYINPUT7), .Z(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n530), .B1(new_n513), .B2(new_n514), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n505), .A2(KEYINPUT71), .A3(new_n506), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n531), .A2(new_n532), .A3(G543), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT72), .B(G51), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT5), .B(G543), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n536), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT70), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n536), .A2(new_n539), .A3(G63), .A4(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n535), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n542), .B1(new_n535), .B2(new_n541), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n526), .B(new_n529), .C1(new_n543), .C2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  AOI22_X1  g121(.A1(new_n536), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n504), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n533), .A2(G52), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n516), .A2(G90), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  AOI22_X1  g127(.A1(new_n533), .A2(G43), .B1(G81), .B2(new_n516), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n510), .A2(new_n512), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT75), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n557), .A2(new_n560), .A3(G651), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n553), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT76), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(G188));
  NAND3_X1  g145(.A1(new_n533), .A2(KEYINPUT9), .A3(G53), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n507), .A2(new_n536), .A3(G91), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n510), .A2(new_n512), .A3(G65), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n504), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n531), .A2(new_n532), .A3(G543), .ZN(new_n579));
  INV_X1    g154(.A(G53), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n571), .A2(new_n577), .A3(new_n581), .ZN(G299));
  NAND2_X1  g157(.A1(new_n533), .A2(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n536), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT77), .B1(new_n515), .B2(new_n585), .ZN(new_n586));
  OR3_X1    g161(.A1(new_n515), .A2(KEYINPUT77), .A3(new_n585), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n583), .A2(new_n584), .A3(new_n586), .A4(new_n587), .ZN(G288));
  AOI22_X1  g163(.A1(new_n536), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT78), .B1(new_n589), .B2(new_n504), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n555), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n593), .A2(new_n594), .A3(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n516), .A2(G86), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n507), .A2(G48), .A3(G543), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n590), .A2(new_n595), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(G305));
  INV_X1    g175(.A(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n579), .A2(new_n601), .B1(new_n602), .B2(new_n515), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n536), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(new_n504), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n579), .A2(KEYINPUT81), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n579), .A2(KEYINPUT81), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n610), .A2(G54), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n515), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT10), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n536), .A2(G66), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT82), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n616), .A2(new_n618), .A3(KEYINPUT83), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n621), .A2(G651), .A3(new_n622), .ZN(new_n623));
  AND3_X1   g198(.A1(new_n612), .A2(new_n615), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n609), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n609), .B1(new_n624), .B2(G868), .ZN(G321));
  NAND2_X1  g201(.A1(G286), .A2(G868), .ZN(new_n627));
  XOR2_X1   g202(.A(G299), .B(KEYINPUT84), .Z(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(G297));
  OAI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(new_n631), .B2(G860), .ZN(G148));
  NAND2_X1  g207(.A1(new_n624), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT85), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n483), .A2(G123), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n486), .A2(G135), .ZN(new_n639));
  NOR2_X1   g214(.A1(G99), .A2(G2105), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(new_n471), .B2(G111), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT12), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2100), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2435), .ZN(new_n650));
  XOR2_X1   g225(.A(G2427), .B(G2438), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT14), .ZN(new_n653));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT86), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n657), .B(new_n660), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(G14), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT88), .ZN(new_n665));
  XOR2_X1   g240(.A(G2067), .B(G2678), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2084), .B(G2090), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT87), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT18), .Z(new_n671));
  XOR2_X1   g246(.A(new_n665), .B(KEYINPUT17), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n672), .A2(new_n666), .A3(new_n669), .ZN(new_n673));
  INV_X1    g248(.A(new_n669), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n672), .B2(new_n666), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n665), .A2(new_n667), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n671), .B(new_n673), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2096), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2100), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G227));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT89), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n684), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(KEYINPUT91), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n685), .A2(new_n688), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT92), .B(G1981), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n695), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT93), .B(G1986), .Z(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n699), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G19), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n563), .B2(new_n705), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(G1341), .Z(new_n708));
  INV_X1    g283(.A(G35), .ZN(new_n709));
  OAI21_X1  g284(.A(KEYINPUT99), .B1(new_n709), .B2(G29), .ZN(new_n710));
  OR3_X1    g285(.A1(new_n709), .A2(KEYINPUT99), .A3(G29), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n710), .B(new_n711), .C1(G162), .C2(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT29), .Z(new_n714));
  INV_X1    g289(.A(G2090), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT100), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n708), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n705), .A2(KEYINPUT23), .A3(G20), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT23), .ZN(new_n720));
  INV_X1    g295(.A(G20), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G16), .ZN(new_n722));
  INV_X1    g297(.A(G299), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n719), .B(new_n722), .C1(new_n723), .C2(new_n705), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1956), .ZN(new_n725));
  OAI21_X1  g300(.A(KEYINPUT96), .B1(G29), .B2(G33), .ZN(new_n726));
  OR3_X1    g301(.A1(KEYINPUT96), .A2(G29), .A3(G33), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n466), .A2(new_n474), .A3(G127), .ZN(new_n728));
  INV_X1    g303(.A(G115), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n460), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G2105), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT25), .Z(new_n733));
  INV_X1    g308(.A(G139), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n731), .B(new_n733), .C1(new_n734), .C2(new_n485), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n726), .B(new_n727), .C1(new_n735), .C2(new_n712), .ZN(new_n736));
  INV_X1    g311(.A(G2072), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR3_X1   g313(.A1(new_n718), .A2(new_n725), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n716), .A2(new_n717), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n705), .A2(G5), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G171), .B2(new_n705), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1961), .ZN(new_n743));
  INV_X1    g318(.A(G2084), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT24), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(G34), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(G34), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n478), .B2(G29), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n743), .B1(new_n744), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n736), .A2(new_n737), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(G28), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(G28), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n753), .A2(new_n754), .A3(new_n712), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n755), .B1(new_n712), .B2(new_n642), .C1(new_n749), .C2(new_n744), .ZN(new_n756));
  INV_X1    g331(.A(G1348), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n624), .A2(G16), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G4), .B2(G16), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n751), .B(new_n756), .C1(new_n757), .C2(new_n759), .ZN(new_n760));
  AND3_X1   g335(.A1(new_n740), .A2(new_n750), .A3(new_n760), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n714), .A2(new_n715), .B1(new_n757), .B2(new_n759), .ZN(new_n762));
  NOR2_X1   g337(.A1(G16), .A2(G21), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G168), .B2(G16), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT98), .B(G1966), .Z(new_n765));
  XOR2_X1   g340(.A(new_n764), .B(new_n765), .Z(new_n766));
  NOR2_X1   g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n712), .A2(G27), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G164), .B2(new_n712), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(G2078), .Z(new_n770));
  NAND4_X1  g345(.A1(new_n739), .A2(new_n761), .A3(new_n767), .A4(new_n770), .ZN(new_n771));
  AOI22_X1  g346(.A1(G129), .A2(new_n483), .B1(new_n486), .B2(G141), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n471), .A2(G105), .A3(G2104), .ZN(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT97), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT26), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n772), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  MUX2_X1   g352(.A(G32), .B(new_n777), .S(G29), .Z(new_n778));
  XOR2_X1   g353(.A(KEYINPUT27), .B(G1996), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n771), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT31), .B(G11), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT36), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n705), .A2(G23), .ZN(new_n784));
  AND4_X1   g359(.A1(new_n583), .A2(new_n584), .A3(new_n586), .A4(new_n587), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n705), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(KEYINPUT33), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(KEYINPUT33), .ZN(new_n788));
  AND3_X1   g363(.A1(new_n787), .A2(G1976), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(G1976), .B1(new_n787), .B2(new_n788), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n705), .A2(G22), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G166), .B2(new_n705), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n792), .A2(G1971), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n792), .A2(G1971), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n789), .A2(new_n790), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(G6), .A2(G16), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G305), .B2(new_n705), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(KEYINPUT32), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT95), .B(G1981), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(KEYINPUT32), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n799), .B1(new_n798), .B2(new_n800), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n795), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n795), .B(KEYINPUT34), .C1(new_n801), .C2(new_n802), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n705), .A2(G24), .ZN(new_n808));
  INV_X1    g383(.A(G290), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n705), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(G1986), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(G1986), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n712), .A2(G25), .ZN(new_n813));
  OR2_X1    g388(.A1(G95), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n815));
  INV_X1    g390(.A(G119), .ZN(new_n816));
  INV_X1    g391(.A(G131), .ZN(new_n817));
  OAI221_X1 g392(.A(new_n815), .B1(new_n482), .B2(new_n816), .C1(new_n817), .C2(new_n485), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(new_n712), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT35), .B(G1991), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT94), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n811), .A2(new_n812), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n783), .B1(new_n807), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g401(.A(KEYINPUT36), .B(new_n824), .C1(new_n805), .C2(new_n806), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n781), .B(new_n782), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT28), .ZN(new_n829));
  INV_X1    g404(.A(G26), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(G29), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(G29), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n483), .A2(G128), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n486), .A2(G140), .ZN(new_n834));
  OR2_X1    g409(.A1(G104), .A2(G2105), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n835), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n832), .B1(new_n837), .B2(G29), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n831), .B1(new_n838), .B2(new_n829), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G2067), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n828), .A2(new_n840), .ZN(G311));
  AOI21_X1  g416(.A(new_n824), .B1(new_n805), .B2(new_n806), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n783), .ZN(new_n843));
  INV_X1    g418(.A(new_n840), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n843), .A2(new_n844), .A3(new_n782), .A4(new_n781), .ZN(G150));
  AOI22_X1  g420(.A1(new_n536), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(new_n504), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n533), .A2(G55), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n516), .A2(G93), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n563), .A2(new_n850), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n562), .A2(new_n848), .A3(new_n847), .A4(new_n849), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n612), .A2(new_n615), .A3(new_n623), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n858), .A2(new_n631), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n857), .B(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n852), .B1(new_n860), .B2(G860), .ZN(G145));
  NAND2_X1  g436(.A1(new_n819), .A2(new_n837), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n818), .A2(new_n833), .A3(new_n834), .A4(new_n836), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(G164), .A2(new_n735), .ZN(new_n865));
  NAND2_X1  g440(.A1(G164), .A2(new_n735), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n645), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n862), .A2(new_n863), .A3(new_n865), .A4(new_n866), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n869), .B1(new_n868), .B2(new_n870), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n483), .A2(G130), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n486), .A2(G142), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n471), .A2(G118), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT101), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n878), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n777), .A2(new_n875), .A3(new_n876), .A4(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n881), .A2(new_n773), .A3(new_n772), .A4(new_n776), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n874), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n880), .A2(new_n882), .A3(new_n874), .ZN(new_n884));
  OAI22_X1  g459(.A1(new_n872), .A2(new_n873), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n873), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n884), .A2(new_n883), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(new_n887), .A3(new_n871), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n642), .B(new_n478), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n490), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT103), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(G37), .B1(new_n889), .B2(new_n892), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n885), .A2(new_n888), .A3(new_n895), .A4(new_n891), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g473(.A1(new_n850), .A2(G868), .ZN(new_n899));
  NOR2_X1   g474(.A1(G305), .A2(G303), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(G305), .A2(G303), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n605), .A2(G288), .A3(new_n607), .ZN(new_n903));
  NAND2_X1  g478(.A1(G290), .A2(new_n785), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n901), .A2(new_n902), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n903), .ZN(new_n906));
  INV_X1    g481(.A(new_n902), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n906), .B1(new_n907), .B2(new_n900), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT104), .ZN(new_n911));
  XOR2_X1   g486(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n912));
  XNOR2_X1  g487(.A(new_n911), .B(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n853), .A2(new_n854), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n633), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n858), .B(new_n723), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n858), .B(G299), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(KEYINPUT41), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n917), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(KEYINPUT106), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n913), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n923), .B(KEYINPUT106), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n913), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n899), .B1(new_n927), .B2(G868), .ZN(G295));
  AOI21_X1  g503(.A(new_n899), .B1(new_n927), .B2(G868), .ZN(G331));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  AND2_X1   g505(.A1(G286), .A2(G171), .ZN(new_n931));
  NOR2_X1   g506(.A1(G286), .A2(G171), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n855), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(G168), .A2(G301), .ZN(new_n934));
  NAND2_X1  g509(.A1(G286), .A2(G171), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n914), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n936), .A3(new_n916), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT108), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n914), .B1(new_n934), .B2(new_n935), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n931), .A2(new_n932), .A3(new_n855), .ZN(new_n940));
  OAI22_X1  g515(.A1(new_n939), .A2(new_n940), .B1(new_n919), .B2(new_n921), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n933), .A2(new_n936), .A3(new_n942), .A4(new_n916), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n938), .A2(new_n909), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G37), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT109), .B1(new_n918), .B2(KEYINPUT41), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT110), .B1(new_n916), .B2(new_n920), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n918), .A2(new_n949), .A3(KEYINPUT41), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n916), .A2(new_n951), .A3(new_n920), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n947), .A2(new_n948), .A3(new_n950), .A4(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(new_n940), .B2(new_n939), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n909), .B1(new_n954), .B2(new_n937), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n930), .B1(new_n946), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n938), .A2(new_n943), .A3(new_n941), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n910), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n958), .A2(KEYINPUT43), .A3(new_n945), .A4(new_n944), .ZN(new_n959));
  XNOR2_X1  g534(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n956), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT43), .B1(new_n946), .B2(new_n955), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n958), .A2(new_n930), .A3(new_n945), .A4(new_n944), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(KEYINPUT44), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n961), .A2(new_n964), .ZN(G397));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n494), .B2(new_n501), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT111), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n481), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n477), .B(G40), .C1(new_n971), .C2(G2105), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT46), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n837), .B(G2067), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n973), .B1(new_n777), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n979), .B(KEYINPUT47), .Z(new_n980));
  INV_X1    g555(.A(new_n973), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n973), .A2(G1996), .A3(new_n777), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n777), .A2(G1996), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n973), .B1(new_n977), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(new_n983), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n818), .A2(new_n821), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n837), .A2(G2067), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n981), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n818), .A2(new_n821), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n973), .B1(new_n993), .B2(new_n989), .ZN(new_n994));
  OR2_X1    g569(.A1(G290), .A2(G1986), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n995), .A2(KEYINPUT112), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(KEYINPUT112), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n973), .A3(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT48), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n988), .A2(new_n994), .A3(new_n999), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n980), .A2(new_n992), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1971), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n967), .A2(new_n969), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n493), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n481), .B2(G126), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n500), .B(new_n498), .C1(new_n1006), .C2(new_n471), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1007), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n1008));
  INV_X1    g583(.A(G40), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n469), .A2(new_n1009), .A3(new_n476), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1002), .B1(new_n1004), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT115), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(new_n1007), .B2(new_n966), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1015), .B(new_n966), .C1(new_n494), .C2(new_n501), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1019), .A2(new_n1010), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1014), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1012), .B1(new_n1021), .B2(G2090), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n1023));
  NAND3_X1  g598(.A1(G303), .A2(new_n1023), .A3(G8), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1023), .B1(G303), .B2(G8), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT116), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1026), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n1024), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1022), .A2(new_n1031), .A3(G8), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1022), .A2(new_n1031), .A3(KEYINPUT117), .A4(G8), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1028), .A2(new_n1024), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1020), .A2(new_n715), .A3(new_n1013), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1012), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G8), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n967), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1040), .B1(new_n1042), .B2(new_n1010), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G288), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT52), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT49), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT118), .B(G86), .Z(new_n1049));
  NAND2_X1  g624(.A1(new_n516), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n590), .A2(new_n595), .A3(new_n597), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G1981), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n598), .A2(G1981), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1048), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n598), .A2(G1981), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(KEYINPUT49), .A3(new_n1052), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(new_n1057), .A3(new_n1043), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT52), .B1(G288), .B2(new_n1045), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1043), .B(new_n1059), .C1(new_n1045), .C2(G288), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1047), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1047), .A2(new_n1058), .A3(new_n1060), .A4(KEYINPUT119), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g640(.A(KEYINPUT115), .B(new_n1015), .C1(new_n1007), .C2(new_n966), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1017), .B1(new_n967), .B2(KEYINPUT50), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1019), .A2(new_n1010), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n744), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n765), .B1(new_n1004), .B2(new_n1011), .ZN(new_n1071));
  AOI211_X1 g646(.A(new_n1040), .B(G286), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1036), .A2(new_n1041), .A3(new_n1065), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT63), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1061), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1022), .A2(G8), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1074), .B1(new_n1077), .B2(new_n1037), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1036), .A2(new_n1076), .A3(new_n1072), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1036), .A2(new_n1061), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1058), .A2(new_n1045), .A3(new_n785), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1044), .B1(new_n1082), .B2(new_n1056), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1087), .B2(G286), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1070), .A2(new_n1071), .A3(G168), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G8), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1086), .B1(new_n1089), .B2(G8), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT62), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1092), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT62), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1094), .B(new_n1095), .C1(new_n1090), .C2(new_n1088), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1004), .A2(new_n1011), .A3(G2078), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1097), .A2(KEYINPUT53), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1069), .A2(G1961), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(KEYINPUT53), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1093), .A2(new_n1096), .A3(G171), .A4(new_n1101), .ZN(new_n1102));
  OR3_X1    g677(.A1(new_n967), .A2(new_n972), .A3(G2067), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1069), .B2(G1348), .ZN(new_n1104));
  INV_X1    g679(.A(G1956), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1068), .B2(new_n1016), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n573), .B2(new_n576), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n536), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n1109));
  OAI211_X1 g684(.A(KEYINPUT121), .B(new_n572), .C1(new_n1109), .C2(new_n504), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1108), .A2(new_n571), .A3(new_n1110), .A4(new_n581), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1113), .A2(KEYINPUT57), .A3(G299), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1003), .A2(new_n1010), .A3(new_n1008), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1111), .A2(KEYINPUT120), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1106), .A2(new_n1114), .A3(new_n1116), .A4(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1104), .A2(new_n624), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1106), .A2(new_n1116), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1114), .A2(new_n1119), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1124), .A2(KEYINPUT61), .A3(new_n1120), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT61), .B1(new_n1124), .B2(new_n1120), .ZN(new_n1127));
  OAI22_X1  g702(.A1(new_n1126), .A2(KEYINPUT125), .B1(new_n1127), .B2(KEYINPUT124), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1127), .A2(KEYINPUT124), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1124), .A2(KEYINPUT125), .A3(KEYINPUT61), .A4(new_n1120), .ZN(new_n1130));
  NOR2_X1   g705(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT58), .B(G1341), .Z(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n967), .B2(new_n972), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1003), .A2(new_n974), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1136));
  OAI211_X1 g711(.A(KEYINPUT122), .B(new_n1132), .C1(new_n967), .C2(new_n972), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n562), .B1(KEYINPUT123), .B2(KEYINPUT59), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1131), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1138), .A2(new_n1131), .A3(new_n1139), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1130), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1128), .A2(new_n1129), .A3(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(KEYINPUT60), .B(new_n1103), .C1(new_n1069), .C2(G1348), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1144), .A2(KEYINPUT126), .A3(new_n858), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n858), .B1(new_n1144), .B2(KEYINPUT126), .ZN(new_n1146));
  OAI22_X1  g721(.A1(new_n1145), .A2(new_n1146), .B1(KEYINPUT126), .B2(new_n1144), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1104), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1125), .B1(new_n1143), .B2(new_n1150), .ZN(new_n1151));
  XOR2_X1   g726(.A(G301), .B(KEYINPUT54), .Z(new_n1152));
  NOR2_X1   g727(.A1(new_n1011), .A2(G2078), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n970), .A2(KEYINPUT53), .A3(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1098), .A2(new_n1099), .A3(new_n1152), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1101), .ZN(new_n1156));
  OAI221_X1 g731(.A(new_n1155), .B1(new_n1152), .B2(new_n1156), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1102), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1036), .A2(new_n1041), .A3(new_n1065), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1085), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n973), .A2(G1986), .A3(G290), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n998), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT113), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1163), .A2(new_n994), .A3(new_n988), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1001), .B1(new_n1160), .B2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g740(.A1(new_n956), .A2(new_n458), .A3(new_n959), .ZN(new_n1167));
  AND3_X1   g741(.A1(new_n897), .A2(new_n662), .A3(new_n679), .ZN(new_n1168));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n1169));
  NAND4_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .A4(new_n703), .ZN(new_n1170));
  NAND4_X1  g744(.A1(new_n956), .A2(new_n959), .A3(new_n458), .A4(new_n703), .ZN(new_n1171));
  NAND3_X1  g745(.A1(new_n897), .A2(new_n662), .A3(new_n679), .ZN(new_n1172));
  OAI21_X1  g746(.A(KEYINPUT127), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1173), .ZN(G308));
  NAND3_X1  g748(.A1(new_n1167), .A2(new_n703), .A3(new_n1168), .ZN(G225));
endmodule


