

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(G651), .A2(n618), .ZN(n638) );
  XNOR2_X2 U551 ( .A(n676), .B(n675), .ZN(n763) );
  NOR2_X2 U552 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  XNOR2_X1 U553 ( .A(n679), .B(KEYINPUT30), .ZN(n680) );
  NAND2_X1 U554 ( .A1(n775), .A2(n773), .ZN(n730) );
  NOR2_X1 U555 ( .A1(n673), .A2(G1384), .ZN(n775) );
  NAND2_X1 U556 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U557 ( .A1(n568), .A2(n567), .ZN(n570) );
  AND2_X1 U558 ( .A1(n541), .A2(n540), .ZN(G160) );
  NOR2_X2 U559 ( .A1(G2104), .A2(n542), .ZN(n598) );
  AND2_X1 U560 ( .A1(n544), .A2(n543), .ZN(n517) );
  NOR2_X1 U561 ( .A1(n740), .A2(n677), .ZN(n518) );
  XOR2_X2 U562 ( .A(KEYINPUT17), .B(n533), .Z(n893) );
  INV_X1 U563 ( .A(G8), .ZN(n677) );
  INV_X1 U564 ( .A(KEYINPUT93), .ZN(n679) );
  XNOR2_X1 U565 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U566 ( .A1(G168), .A2(n682), .ZN(n683) );
  INV_X1 U567 ( .A(KEYINPUT29), .ZN(n722) );
  XNOR2_X1 U568 ( .A(n723), .B(n722), .ZN(n726) );
  INV_X1 U569 ( .A(KEYINPUT97), .ZN(n736) );
  XNOR2_X1 U570 ( .A(n737), .B(n736), .ZN(n738) );
  NAND2_X1 U571 ( .A1(G8), .A2(n730), .ZN(n676) );
  INV_X1 U572 ( .A(KEYINPUT12), .ZN(n561) );
  INV_X1 U573 ( .A(n1019), .ZN(n755) );
  XNOR2_X1 U574 ( .A(n561), .B(KEYINPUT69), .ZN(n562) );
  XNOR2_X1 U575 ( .A(n563), .B(n562), .ZN(n565) );
  NOR2_X1 U576 ( .A1(n758), .A2(n757), .ZN(n771) );
  XNOR2_X1 U577 ( .A(n523), .B(KEYINPUT64), .ZN(n640) );
  OR2_X1 U578 ( .A1(G2105), .A2(n534), .ZN(n535) );
  NAND2_X1 U579 ( .A1(n570), .A2(n569), .ZN(n1015) );
  INV_X1 U580 ( .A(G651), .ZN(n525) );
  NOR2_X1 U581 ( .A1(G543), .A2(n525), .ZN(n519) );
  XOR2_X2 U582 ( .A(KEYINPUT1), .B(n519), .Z(n639) );
  NAND2_X1 U583 ( .A1(G63), .A2(n639), .ZN(n521) );
  XOR2_X1 U584 ( .A(KEYINPUT0), .B(G543), .Z(n618) );
  NAND2_X1 U585 ( .A1(G51), .A2(n638), .ZN(n520) );
  NAND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U587 ( .A(KEYINPUT6), .B(n522), .ZN(n530) );
  NOR2_X1 U588 ( .A1(G543), .A2(G651), .ZN(n523) );
  NAND2_X1 U589 ( .A1(G89), .A2(n640), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(KEYINPUT4), .ZN(n527) );
  NOR2_X1 U591 ( .A1(n618), .A2(n525), .ZN(n643) );
  NAND2_X1 U592 ( .A1(G76), .A2(n643), .ZN(n526) );
  NAND2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U594 ( .A(n528), .B(KEYINPUT5), .Z(n529) );
  NOR2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U596 ( .A(KEYINPUT7), .B(n531), .Z(n532) );
  XOR2_X1 U597 ( .A(KEYINPUT71), .B(n532), .Z(G168) );
  XOR2_X1 U598 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U599 ( .A1(n893), .A2(G137), .ZN(n541) );
  NAND2_X1 U600 ( .A1(G2104), .A2(G101), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(KEYINPUT23), .ZN(n539) );
  AND2_X1 U602 ( .A1(G2104), .A2(G2105), .ZN(n890) );
  NAND2_X1 U603 ( .A1(G113), .A2(n890), .ZN(n537) );
  INV_X1 U604 ( .A(G2105), .ZN(n542) );
  NAND2_X1 U605 ( .A1(G125), .A2(n598), .ZN(n536) );
  NAND2_X1 U606 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n540) );
  AND2_X1 U608 ( .A1(G138), .A2(n893), .ZN(n547) );
  AND2_X1 U609 ( .A1(n542), .A2(G2104), .ZN(n895) );
  NAND2_X1 U610 ( .A1(G102), .A2(n895), .ZN(n545) );
  NAND2_X1 U611 ( .A1(G114), .A2(n890), .ZN(n544) );
  NAND2_X1 U612 ( .A1(G126), .A2(n598), .ZN(n543) );
  NAND2_X1 U613 ( .A1(n545), .A2(n517), .ZN(n546) );
  NOR2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n549) );
  INV_X1 U615 ( .A(KEYINPUT81), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n673) );
  BUF_X1 U617 ( .A(n673), .Z(G164) );
  NAND2_X1 U618 ( .A1(G64), .A2(n639), .ZN(n551) );
  NAND2_X1 U619 ( .A1(G52), .A2(n638), .ZN(n550) );
  NAND2_X1 U620 ( .A1(n551), .A2(n550), .ZN(n556) );
  NAND2_X1 U621 ( .A1(n643), .A2(G77), .ZN(n553) );
  NAND2_X1 U622 ( .A1(G90), .A2(n640), .ZN(n552) );
  NAND2_X1 U623 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U624 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U625 ( .A1(n556), .A2(n555), .ZN(G171) );
  AND2_X1 U626 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U627 ( .A(G57), .ZN(G237) );
  INV_X1 U628 ( .A(G82), .ZN(G220) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n557) );
  XNOR2_X1 U630 ( .A(n557), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U631 ( .A(KEYINPUT68), .B(KEYINPUT11), .Z(n559) );
  INV_X1 U632 ( .A(G223), .ZN(n825) );
  NAND2_X1 U633 ( .A1(G567), .A2(n825), .ZN(n558) );
  XNOR2_X1 U634 ( .A(n559), .B(n558), .ZN(G234) );
  NAND2_X1 U635 ( .A1(G56), .A2(n639), .ZN(n560) );
  XOR2_X1 U636 ( .A(KEYINPUT14), .B(n560), .Z(n568) );
  NAND2_X1 U637 ( .A1(n640), .A2(G81), .ZN(n563) );
  NAND2_X1 U638 ( .A1(G68), .A2(n643), .ZN(n564) );
  NAND2_X1 U639 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U640 ( .A(KEYINPUT13), .B(n566), .Z(n567) );
  NAND2_X1 U641 ( .A1(n638), .A2(G43), .ZN(n569) );
  INV_X1 U642 ( .A(G860), .ZN(n832) );
  OR2_X1 U643 ( .A1(n1015), .A2(n832), .ZN(G153) );
  INV_X1 U644 ( .A(G171), .ZN(G301) );
  NAND2_X1 U645 ( .A1(G66), .A2(n639), .ZN(n572) );
  NAND2_X1 U646 ( .A1(G92), .A2(n640), .ZN(n571) );
  NAND2_X1 U647 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U648 ( .A1(G79), .A2(n643), .ZN(n574) );
  NAND2_X1 U649 ( .A1(G54), .A2(n638), .ZN(n573) );
  NAND2_X1 U650 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U651 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U652 ( .A(KEYINPUT70), .B(KEYINPUT15), .ZN(n577) );
  XNOR2_X2 U653 ( .A(n578), .B(n577), .ZN(n1012) );
  NOR2_X1 U654 ( .A1(n1012), .A2(G868), .ZN(n580) );
  INV_X1 U655 ( .A(G868), .ZN(n655) );
  NOR2_X1 U656 ( .A1(n655), .A2(G301), .ZN(n579) );
  NOR2_X1 U657 ( .A1(n580), .A2(n579), .ZN(G284) );
  NAND2_X1 U658 ( .A1(G65), .A2(n639), .ZN(n582) );
  NAND2_X1 U659 ( .A1(G91), .A2(n640), .ZN(n581) );
  NAND2_X1 U660 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U661 ( .A1(n643), .A2(G78), .ZN(n583) );
  XOR2_X1 U662 ( .A(KEYINPUT66), .B(n583), .Z(n584) );
  NOR2_X1 U663 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U664 ( .A1(n638), .A2(G53), .ZN(n586) );
  NAND2_X1 U665 ( .A1(n587), .A2(n586), .ZN(G299) );
  NOR2_X1 U666 ( .A1(G286), .A2(n655), .ZN(n589) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n588) );
  NOR2_X1 U668 ( .A1(n589), .A2(n588), .ZN(G297) );
  NAND2_X1 U669 ( .A1(n832), .A2(G559), .ZN(n590) );
  INV_X1 U670 ( .A(n1012), .ZN(n635) );
  NAND2_X1 U671 ( .A1(n590), .A2(n635), .ZN(n591) );
  XNOR2_X1 U672 ( .A(n591), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n1015), .ZN(n594) );
  NAND2_X1 U674 ( .A1(n635), .A2(G868), .ZN(n592) );
  NOR2_X1 U675 ( .A1(G559), .A2(n592), .ZN(n593) );
  NOR2_X1 U676 ( .A1(n594), .A2(n593), .ZN(G282) );
  NAND2_X1 U677 ( .A1(G135), .A2(n893), .ZN(n595) );
  XNOR2_X1 U678 ( .A(n595), .B(KEYINPUT72), .ZN(n603) );
  NAND2_X1 U679 ( .A1(G99), .A2(n895), .ZN(n597) );
  NAND2_X1 U680 ( .A1(G111), .A2(n890), .ZN(n596) );
  NAND2_X1 U681 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U682 ( .A1(n598), .A2(G123), .ZN(n599) );
  XOR2_X1 U683 ( .A(KEYINPUT18), .B(n599), .Z(n600) );
  NOR2_X1 U684 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U685 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U686 ( .A(KEYINPUT73), .B(n604), .ZN(n976) );
  XNOR2_X1 U687 ( .A(n976), .B(G2096), .ZN(n606) );
  INV_X1 U688 ( .A(G2100), .ZN(n605) );
  NAND2_X1 U689 ( .A1(n606), .A2(n605), .ZN(G156) );
  NAND2_X1 U690 ( .A1(n643), .A2(G73), .ZN(n607) );
  XOR2_X1 U691 ( .A(KEYINPUT2), .B(n607), .Z(n612) );
  NAND2_X1 U692 ( .A1(G86), .A2(n640), .ZN(n609) );
  NAND2_X1 U693 ( .A1(n639), .A2(G61), .ZN(n608) );
  NAND2_X1 U694 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U695 ( .A(KEYINPUT76), .B(n610), .ZN(n611) );
  NOR2_X1 U696 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U697 ( .A1(n638), .A2(G48), .ZN(n613) );
  NAND2_X1 U698 ( .A1(n614), .A2(n613), .ZN(G305) );
  NAND2_X1 U699 ( .A1(G49), .A2(n638), .ZN(n616) );
  NAND2_X1 U700 ( .A1(G74), .A2(G651), .ZN(n615) );
  NAND2_X1 U701 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U702 ( .A1(n639), .A2(n617), .ZN(n620) );
  NAND2_X1 U703 ( .A1(n618), .A2(G87), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(G288) );
  NAND2_X1 U705 ( .A1(G62), .A2(n639), .ZN(n622) );
  NAND2_X1 U706 ( .A1(G88), .A2(n640), .ZN(n621) );
  NAND2_X1 U707 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U708 ( .A1(G75), .A2(n643), .ZN(n623) );
  XNOR2_X1 U709 ( .A(KEYINPUT77), .B(n623), .ZN(n624) );
  NOR2_X1 U710 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n638), .A2(G50), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n627), .A2(n626), .ZN(G303) );
  INV_X1 U713 ( .A(G303), .ZN(G166) );
  NAND2_X1 U714 ( .A1(n643), .A2(G72), .ZN(n629) );
  NAND2_X1 U715 ( .A1(G85), .A2(n640), .ZN(n628) );
  NAND2_X1 U716 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U717 ( .A(KEYINPUT65), .B(n630), .ZN(n634) );
  NAND2_X1 U718 ( .A1(G60), .A2(n639), .ZN(n632) );
  NAND2_X1 U719 ( .A1(G47), .A2(n638), .ZN(n631) );
  AND2_X1 U720 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U721 ( .A1(n634), .A2(n633), .ZN(G290) );
  NAND2_X1 U722 ( .A1(n635), .A2(G559), .ZN(n636) );
  XOR2_X1 U723 ( .A(n1015), .B(n636), .Z(n831) );
  XNOR2_X1 U724 ( .A(KEYINPUT19), .B(G305), .ZN(n637) );
  XNOR2_X1 U725 ( .A(n637), .B(G288), .ZN(n650) );
  NAND2_X1 U726 ( .A1(G55), .A2(n638), .ZN(n648) );
  NAND2_X1 U727 ( .A1(G67), .A2(n639), .ZN(n642) );
  NAND2_X1 U728 ( .A1(G93), .A2(n640), .ZN(n641) );
  NAND2_X1 U729 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U730 ( .A1(n643), .A2(G80), .ZN(n644) );
  XOR2_X1 U731 ( .A(KEYINPUT74), .B(n644), .Z(n645) );
  NOR2_X1 U732 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U733 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U734 ( .A(n649), .B(KEYINPUT75), .Z(n833) );
  XNOR2_X1 U735 ( .A(n650), .B(n833), .ZN(n652) );
  INV_X1 U736 ( .A(G299), .ZN(n698) );
  XNOR2_X1 U737 ( .A(n698), .B(G166), .ZN(n651) );
  XNOR2_X1 U738 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U739 ( .A(n653), .B(G290), .ZN(n908) );
  XNOR2_X1 U740 ( .A(n831), .B(n908), .ZN(n654) );
  NAND2_X1 U741 ( .A1(n654), .A2(G868), .ZN(n657) );
  NAND2_X1 U742 ( .A1(n655), .A2(n833), .ZN(n656) );
  NAND2_X1 U743 ( .A1(n657), .A2(n656), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2078), .A2(G2084), .ZN(n658) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n658), .Z(n659) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n659), .ZN(n660) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n660), .ZN(n661) );
  NAND2_X1 U748 ( .A1(n661), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(KEYINPUT67), .B(G132), .ZN(G219) );
  XNOR2_X1 U750 ( .A(KEYINPUT78), .B(G44), .ZN(n662) );
  XNOR2_X1 U751 ( .A(n662), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U752 ( .A1(G220), .A2(G219), .ZN(n663) );
  XNOR2_X1 U753 ( .A(KEYINPUT22), .B(n663), .ZN(n664) );
  NAND2_X1 U754 ( .A1(n664), .A2(G96), .ZN(n665) );
  NOR2_X1 U755 ( .A1(n665), .A2(G218), .ZN(n666) );
  XNOR2_X1 U756 ( .A(n666), .B(KEYINPUT79), .ZN(n829) );
  NAND2_X1 U757 ( .A1(n829), .A2(G2106), .ZN(n670) );
  NAND2_X1 U758 ( .A1(G69), .A2(G120), .ZN(n667) );
  NOR2_X1 U759 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U760 ( .A1(G108), .A2(n668), .ZN(n830) );
  NAND2_X1 U761 ( .A1(n830), .A2(G567), .ZN(n669) );
  NAND2_X1 U762 ( .A1(n670), .A2(n669), .ZN(n919) );
  NAND2_X1 U763 ( .A1(G483), .A2(G661), .ZN(n671) );
  NOR2_X1 U764 ( .A1(n919), .A2(n671), .ZN(n828) );
  NAND2_X1 U765 ( .A1(n828), .A2(G36), .ZN(n672) );
  XNOR2_X1 U766 ( .A(KEYINPUT80), .B(n672), .ZN(G176) );
  NAND2_X1 U767 ( .A1(G40), .A2(G160), .ZN(n674) );
  XNOR2_X1 U768 ( .A(n674), .B(KEYINPUT83), .ZN(n773) );
  INV_X1 U769 ( .A(KEYINPUT87), .ZN(n675) );
  NOR2_X1 U770 ( .A1(G1966), .A2(n763), .ZN(n743) );
  INV_X1 U771 ( .A(n743), .ZN(n678) );
  NOR2_X1 U772 ( .A1(G2084), .A2(n730), .ZN(n740) );
  NAND2_X1 U773 ( .A1(n678), .A2(n518), .ZN(n681) );
  XNOR2_X1 U774 ( .A(n683), .B(KEYINPUT94), .ZN(n689) );
  XOR2_X1 U775 ( .A(G2078), .B(KEYINPUT25), .Z(n929) );
  NOR2_X1 U776 ( .A1(n929), .A2(n730), .ZN(n684) );
  XNOR2_X1 U777 ( .A(n684), .B(KEYINPUT88), .ZN(n686) );
  INV_X1 U778 ( .A(n730), .ZN(n711) );
  NOR2_X1 U779 ( .A1(n711), .A2(G1961), .ZN(n685) );
  NOR2_X1 U780 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U781 ( .A(KEYINPUT89), .B(n687), .ZN(n724) );
  NOR2_X1 U782 ( .A1(n724), .A2(G171), .ZN(n688) );
  NOR2_X1 U783 ( .A1(n689), .A2(n688), .ZN(n691) );
  XNOR2_X1 U784 ( .A(KEYINPUT95), .B(KEYINPUT31), .ZN(n690) );
  XNOR2_X1 U785 ( .A(n691), .B(n690), .ZN(n728) );
  NAND2_X1 U786 ( .A1(G2072), .A2(n711), .ZN(n692) );
  XNOR2_X1 U787 ( .A(n692), .B(KEYINPUT27), .ZN(n693) );
  XNOR2_X1 U788 ( .A(n693), .B(KEYINPUT90), .ZN(n695) );
  INV_X1 U789 ( .A(G1956), .ZN(n951) );
  NOR2_X1 U790 ( .A1(n951), .A2(n711), .ZN(n694) );
  NOR2_X1 U791 ( .A1(n695), .A2(n694), .ZN(n699) );
  NOR2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n697) );
  XNOR2_X1 U793 ( .A(KEYINPUT91), .B(KEYINPUT28), .ZN(n696) );
  XNOR2_X1 U794 ( .A(n697), .B(n696), .ZN(n721) );
  NAND2_X1 U795 ( .A1(n699), .A2(n698), .ZN(n719) );
  NOR2_X1 U796 ( .A1(KEYINPUT26), .A2(G1996), .ZN(n700) );
  NOR2_X1 U797 ( .A1(n1015), .A2(n700), .ZN(n705) );
  NAND2_X1 U798 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n702) );
  NAND2_X1 U799 ( .A1(G2067), .A2(n1012), .ZN(n701) );
  NAND2_X1 U800 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U801 ( .A1(n711), .A2(n703), .ZN(n704) );
  NAND2_X1 U802 ( .A1(n705), .A2(n704), .ZN(n710) );
  NAND2_X1 U803 ( .A1(n1012), .A2(G1348), .ZN(n706) );
  NAND2_X1 U804 ( .A1(KEYINPUT26), .A2(n706), .ZN(n707) );
  NOR2_X1 U805 ( .A1(G1341), .A2(n707), .ZN(n708) );
  NOR2_X1 U806 ( .A1(n711), .A2(n708), .ZN(n709) );
  NOR2_X1 U807 ( .A1(n710), .A2(n709), .ZN(n716) );
  NAND2_X1 U808 ( .A1(G1348), .A2(n730), .ZN(n713) );
  NAND2_X1 U809 ( .A1(n711), .A2(G2067), .ZN(n712) );
  NAND2_X1 U810 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U811 ( .A1(n1012), .A2(n714), .ZN(n715) );
  NOR2_X1 U812 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U813 ( .A(KEYINPUT92), .B(n717), .ZN(n718) );
  NAND2_X1 U814 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U815 ( .A1(n721), .A2(n720), .ZN(n723) );
  NAND2_X1 U816 ( .A1(n724), .A2(G171), .ZN(n725) );
  NAND2_X1 U817 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U818 ( .A1(n728), .A2(n727), .ZN(n741) );
  NAND2_X1 U819 ( .A1(n741), .A2(G286), .ZN(n729) );
  XNOR2_X1 U820 ( .A(n729), .B(KEYINPUT96), .ZN(n735) );
  NOR2_X1 U821 ( .A1(G2090), .A2(n730), .ZN(n732) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n763), .ZN(n731) );
  NOR2_X1 U823 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U824 ( .A1(n733), .A2(G303), .ZN(n734) );
  NAND2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U826 ( .A1(n738), .A2(G8), .ZN(n739) );
  XNOR2_X1 U827 ( .A(n739), .B(KEYINPUT32), .ZN(n747) );
  NAND2_X1 U828 ( .A1(G8), .A2(n740), .ZN(n745) );
  INV_X1 U829 ( .A(n741), .ZN(n742) );
  NOR2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U831 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U832 ( .A1(n747), .A2(n746), .ZN(n761) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n1001) );
  NOR2_X1 U834 ( .A1(G1971), .A2(G303), .ZN(n748) );
  XNOR2_X1 U835 ( .A(KEYINPUT98), .B(n748), .ZN(n749) );
  NOR2_X1 U836 ( .A1(n1001), .A2(n749), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n761), .A2(n750), .ZN(n751) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n1002) );
  NAND2_X1 U839 ( .A1(n751), .A2(n1002), .ZN(n752) );
  NOR2_X1 U840 ( .A1(n752), .A2(n763), .ZN(n753) );
  NOR2_X1 U841 ( .A1(KEYINPUT33), .A2(n753), .ZN(n758) );
  AND2_X1 U842 ( .A1(n1001), .A2(KEYINPUT33), .ZN(n754) );
  INV_X1 U843 ( .A(n763), .ZN(n766) );
  NAND2_X1 U844 ( .A1(n754), .A2(n766), .ZN(n756) );
  XNOR2_X1 U845 ( .A(G1981), .B(G305), .ZN(n1019) );
  NOR2_X1 U846 ( .A1(G2090), .A2(G303), .ZN(n759) );
  NAND2_X1 U847 ( .A1(G8), .A2(n759), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n762) );
  AND2_X1 U849 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U850 ( .A(n764), .B(KEYINPUT99), .ZN(n769) );
  NOR2_X1 U851 ( .A1(G1981), .A2(G305), .ZN(n765) );
  XNOR2_X1 U852 ( .A(n765), .B(KEYINPUT24), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U854 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U855 ( .A1(n771), .A2(n770), .ZN(n806) );
  XNOR2_X1 U856 ( .A(KEYINPUT82), .B(G1986), .ZN(n772) );
  XNOR2_X1 U857 ( .A(n772), .B(G290), .ZN(n1007) );
  INV_X1 U858 ( .A(n773), .ZN(n774) );
  NOR2_X1 U859 ( .A1(n775), .A2(n774), .ZN(n819) );
  AND2_X1 U860 ( .A1(n1007), .A2(n819), .ZN(n804) );
  XNOR2_X1 U861 ( .A(G2067), .B(KEYINPUT37), .ZN(n817) );
  NAND2_X1 U862 ( .A1(G140), .A2(n893), .ZN(n777) );
  NAND2_X1 U863 ( .A1(G104), .A2(n895), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U865 ( .A(KEYINPUT34), .B(n778), .ZN(n783) );
  NAND2_X1 U866 ( .A1(G116), .A2(n890), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G128), .A2(n598), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U869 ( .A(KEYINPUT35), .B(n781), .Z(n782) );
  NOR2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U871 ( .A(KEYINPUT36), .B(n784), .ZN(n872) );
  NOR2_X1 U872 ( .A1(n817), .A2(n872), .ZN(n978) );
  NAND2_X1 U873 ( .A1(n819), .A2(n978), .ZN(n816) );
  NAND2_X1 U874 ( .A1(G131), .A2(n893), .ZN(n786) );
  NAND2_X1 U875 ( .A1(G95), .A2(n895), .ZN(n785) );
  NAND2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n598), .A2(G119), .ZN(n787) );
  XOR2_X1 U878 ( .A(KEYINPUT84), .B(n787), .Z(n788) );
  NOR2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n890), .A2(G107), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n885) );
  NAND2_X1 U882 ( .A1(G1991), .A2(n885), .ZN(n801) );
  NAND2_X1 U883 ( .A1(G105), .A2(n895), .ZN(n792) );
  XOR2_X1 U884 ( .A(KEYINPUT38), .B(n792), .Z(n797) );
  NAND2_X1 U885 ( .A1(G117), .A2(n890), .ZN(n794) );
  NAND2_X1 U886 ( .A1(G129), .A2(n598), .ZN(n793) );
  NAND2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U888 ( .A(KEYINPUT85), .B(n795), .Z(n796) );
  NOR2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n893), .A2(G141), .ZN(n798) );
  NAND2_X1 U891 ( .A1(n799), .A2(n798), .ZN(n880) );
  NAND2_X1 U892 ( .A1(G1996), .A2(n880), .ZN(n800) );
  NAND2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n983) );
  NAND2_X1 U894 ( .A1(n819), .A2(n983), .ZN(n809) );
  NAND2_X1 U895 ( .A1(n816), .A2(n809), .ZN(n802) );
  XNOR2_X1 U896 ( .A(n802), .B(KEYINPUT86), .ZN(n803) );
  OR2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n805) );
  OR2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n823) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n880), .ZN(n987) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n885), .ZN(n977) );
  NOR2_X1 U902 ( .A1(n807), .A2(n977), .ZN(n808) );
  XOR2_X1 U903 ( .A(KEYINPUT100), .B(n808), .Z(n810) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U905 ( .A(KEYINPUT101), .B(n811), .ZN(n812) );
  NOR2_X1 U906 ( .A1(n987), .A2(n812), .ZN(n814) );
  XNOR2_X1 U907 ( .A(KEYINPUT39), .B(KEYINPUT102), .ZN(n813) );
  XNOR2_X1 U908 ( .A(n814), .B(n813), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n818) );
  NAND2_X1 U910 ( .A1(n817), .A2(n872), .ZN(n984) );
  NAND2_X1 U911 ( .A1(n818), .A2(n984), .ZN(n820) );
  NAND2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U913 ( .A(KEYINPUT103), .B(n821), .Z(n822) );
  NAND2_X1 U914 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U915 ( .A(n824), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n825), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U918 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n828), .A2(n827), .ZN(G188) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(G69), .ZN(G235) );
  NOR2_X1 U925 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  NAND2_X1 U927 ( .A1(n832), .A2(n831), .ZN(n834) );
  XNOR2_X1 U928 ( .A(n834), .B(n833), .ZN(G145) );
  XNOR2_X1 U929 ( .A(G1341), .B(G2454), .ZN(n835) );
  XNOR2_X1 U930 ( .A(n835), .B(G2430), .ZN(n836) );
  XNOR2_X1 U931 ( .A(n836), .B(G1348), .ZN(n842) );
  XOR2_X1 U932 ( .A(G2443), .B(G2427), .Z(n838) );
  XNOR2_X1 U933 ( .A(G2438), .B(G2446), .ZN(n837) );
  XNOR2_X1 U934 ( .A(n838), .B(n837), .ZN(n840) );
  XOR2_X1 U935 ( .A(G2451), .B(G2435), .Z(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n842), .B(n841), .ZN(n843) );
  NAND2_X1 U938 ( .A1(n843), .A2(G14), .ZN(n844) );
  XOR2_X1 U939 ( .A(KEYINPUT104), .B(n844), .Z(G401) );
  XOR2_X1 U940 ( .A(KEYINPUT106), .B(G1991), .Z(n846) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1971), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U943 ( .A(n847), .B(KEYINPUT41), .Z(n849) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1961), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U946 ( .A(G1986), .B(G1956), .Z(n851) );
  XNOR2_X1 U947 ( .A(G1981), .B(G1976), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U949 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U950 ( .A(G2474), .B(KEYINPUT107), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n855), .B(n854), .ZN(G229) );
  XOR2_X1 U952 ( .A(KEYINPUT105), .B(G2090), .Z(n857) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2084), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U955 ( .A(n858), .B(G2100), .Z(n860) );
  XNOR2_X1 U956 ( .A(G2078), .B(G2072), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U958 ( .A(G2096), .B(KEYINPUT43), .Z(n862) );
  XNOR2_X1 U959 ( .A(KEYINPUT42), .B(G2678), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U961 ( .A(n864), .B(n863), .Z(G227) );
  NAND2_X1 U962 ( .A1(G124), .A2(n598), .ZN(n865) );
  XNOR2_X1 U963 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U964 ( .A1(n895), .A2(G100), .ZN(n866) );
  NAND2_X1 U965 ( .A1(n867), .A2(n866), .ZN(n871) );
  NAND2_X1 U966 ( .A1(G136), .A2(n893), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G112), .A2(n890), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U969 ( .A1(n871), .A2(n870), .ZN(G162) );
  XNOR2_X1 U970 ( .A(G160), .B(n872), .ZN(n883) );
  NAND2_X1 U971 ( .A1(G139), .A2(n893), .ZN(n874) );
  NAND2_X1 U972 ( .A1(G103), .A2(n895), .ZN(n873) );
  NAND2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n879) );
  NAND2_X1 U974 ( .A1(G115), .A2(n890), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G127), .A2(n598), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n877), .Z(n878) );
  NOR2_X1 U978 ( .A1(n879), .A2(n878), .ZN(n969) );
  XNOR2_X1 U979 ( .A(n969), .B(G162), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n906) );
  XOR2_X1 U982 ( .A(G164), .B(n976), .Z(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n889) );
  XOR2_X1 U984 ( .A(KEYINPUT48), .B(KEYINPUT110), .Z(n887) );
  XNOR2_X1 U985 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U987 ( .A(n889), .B(n888), .Z(n904) );
  NAND2_X1 U988 ( .A1(G118), .A2(n890), .ZN(n892) );
  NAND2_X1 U989 ( .A1(G130), .A2(n598), .ZN(n891) );
  NAND2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n901) );
  NAND2_X1 U991 ( .A1(n893), .A2(G142), .ZN(n894) );
  XNOR2_X1 U992 ( .A(KEYINPUT109), .B(n894), .ZN(n898) );
  NAND2_X1 U993 ( .A1(n895), .A2(G106), .ZN(n896) );
  XOR2_X1 U994 ( .A(KEYINPUT108), .B(n896), .Z(n897) );
  NOR2_X1 U995 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n899), .B(KEYINPUT45), .ZN(n900) );
  NOR2_X1 U997 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n902), .B(KEYINPUT111), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n907), .ZN(G395) );
  XOR2_X1 U1002 ( .A(n908), .B(G286), .Z(n910) );
  XNOR2_X1 U1003 ( .A(G171), .B(n1012), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1005 ( .A(n911), .B(n1015), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n912), .ZN(G397) );
  OR2_X1 U1007 ( .A1(n919), .A2(G401), .ZN(n916) );
  NOR2_X1 U1008 ( .A1(G229), .A2(G227), .ZN(n913) );
  XOR2_X1 U1009 ( .A(KEYINPUT113), .B(n913), .Z(n914) );
  XNOR2_X1 U1010 ( .A(n914), .B(KEYINPUT49), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(n919), .ZN(G319) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1017 ( .A(G2084), .B(G34), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(n920), .B(KEYINPUT54), .ZN(n937) );
  XNOR2_X1 U1019 ( .A(G2090), .B(G35), .ZN(n934) );
  XNOR2_X1 U1020 ( .A(G2072), .B(G33), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(G2067), .B(G26), .ZN(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n928) );
  XOR2_X1 U1023 ( .A(G1996), .B(G32), .Z(n923) );
  NAND2_X1 U1024 ( .A1(n923), .A2(G28), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(G25), .B(G1991), .ZN(n924) );
  XNOR2_X1 U1026 ( .A(KEYINPUT120), .B(n924), .ZN(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(G27), .B(n929), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(KEYINPUT53), .B(n932), .ZN(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1033 ( .A(n935), .B(KEYINPUT121), .ZN(n936) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1035 ( .A(KEYINPUT55), .B(n938), .Z(n939) );
  XNOR2_X1 U1036 ( .A(KEYINPUT122), .B(n939), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(G29), .A2(n940), .ZN(n968) );
  XNOR2_X1 U1038 ( .A(G1986), .B(G24), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(G1976), .B(G23), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(G22), .B(G1971), .ZN(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1042 ( .A(KEYINPUT127), .B(n943), .ZN(n944) );
  NOR2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(KEYINPUT58), .B(n946), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(G1966), .B(G21), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(G5), .B(G1961), .ZN(n947) );
  NOR2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n962) );
  XNOR2_X1 U1049 ( .A(G20), .B(n951), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G1981), .B(G6), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(G1341), .B(G19), .ZN(n952) );
  NOR2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1054 ( .A(KEYINPUT59), .B(G1348), .Z(n956) );
  XNOR2_X1 U1055 ( .A(G4), .B(n956), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1057 ( .A(KEYINPUT60), .B(n959), .Z(n960) );
  XNOR2_X1 U1058 ( .A(KEYINPUT126), .B(n960), .ZN(n961) );
  NOR2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1060 ( .A(n963), .B(KEYINPUT61), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(G16), .B(KEYINPUT125), .ZN(n964) );
  NAND2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n966), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n1000) );
  XOR2_X1 U1065 ( .A(G2072), .B(n969), .Z(n970) );
  XNOR2_X1 U1066 ( .A(KEYINPUT118), .B(n970), .ZN(n972) );
  XOR2_X1 U1067 ( .A(G164), .B(G2078), .Z(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1069 ( .A(KEYINPUT50), .B(n973), .Z(n994) );
  XOR2_X1 U1070 ( .A(G2084), .B(G160), .Z(n974) );
  XNOR2_X1 U1071 ( .A(KEYINPUT114), .B(n974), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1075 ( .A(KEYINPUT115), .B(n981), .Z(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n991) );
  XOR2_X1 U1078 ( .A(G2090), .B(G162), .Z(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1080 ( .A(KEYINPUT116), .B(n988), .Z(n989) );
  XOR2_X1 U1081 ( .A(KEYINPUT51), .B(n989), .Z(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(KEYINPUT117), .B(n992), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1085 ( .A(KEYINPUT52), .B(n995), .Z(n996) );
  NOR2_X1 U1086 ( .A1(KEYINPUT55), .A2(n996), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(KEYINPUT119), .B(n997), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n998), .A2(G29), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1028) );
  XOR2_X1 U1090 ( .A(KEYINPUT56), .B(G16), .Z(n1026) );
  INV_X1 U1091 ( .A(n1001), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G1956), .B(G299), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(G166), .B(G1971), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(n1006), .B(KEYINPUT123), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(KEYINPUT124), .B(n1011), .ZN(n1024) );
  XOR2_X1 U1100 ( .A(n1012), .B(G1348), .Z(n1014) );
  XNOR2_X1 U1101 ( .A(G171), .B(G1961), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(G1341), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1022) );
  XOR2_X1 U1105 ( .A(G1966), .B(G168), .Z(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1107 ( .A(KEYINPUT57), .B(n1020), .Z(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1112 ( .A(n1029), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

