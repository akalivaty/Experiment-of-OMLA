

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740;

  XNOR2_X1 U364 ( .A(n571), .B(n355), .ZN(n423) );
  NOR2_X1 U365 ( .A1(n581), .A2(n654), .ZN(n556) );
  NOR2_X1 U366 ( .A1(n543), .A2(n544), .ZN(n633) );
  XNOR2_X2 U367 ( .A(n370), .B(n347), .ZN(n567) );
  XNOR2_X2 U368 ( .A(n457), .B(n344), .ZN(n381) );
  XNOR2_X2 U369 ( .A(n583), .B(KEYINPUT41), .ZN(n685) );
  NOR2_X2 U370 ( .A1(n672), .A2(n671), .ZN(n583) );
  XNOR2_X2 U371 ( .A(KEYINPUT66), .B(G143), .ZN(n452) );
  INV_X2 U372 ( .A(G953), .ZN(n726) );
  AND2_X1 U373 ( .A1(n409), .A2(n406), .ZN(n389) );
  AND2_X1 U374 ( .A1(n411), .A2(n410), .ZN(n409) );
  XOR2_X1 U375 ( .A(n527), .B(KEYINPUT35), .Z(n537) );
  NAND2_X1 U376 ( .A1(n408), .A2(n407), .ZN(n406) );
  AND2_X1 U377 ( .A1(n570), .A2(n546), .ZN(n397) );
  NOR2_X1 U378 ( .A1(n528), .A2(n543), .ZN(n582) );
  XNOR2_X1 U379 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U380 ( .A(n398), .B(n455), .ZN(n693) );
  XNOR2_X1 U381 ( .A(n718), .B(n375), .ZN(n398) );
  XNOR2_X1 U382 ( .A(n374), .B(n510), .ZN(n718) );
  XNOR2_X1 U383 ( .A(n377), .B(n376), .ZN(n375) );
  XNOR2_X1 U384 ( .A(n496), .B(KEYINPUT16), .ZN(n374) );
  XNOR2_X1 U385 ( .A(n417), .B(n456), .ZN(n601) );
  XNOR2_X1 U386 ( .A(G110), .B(G107), .ZN(n453) );
  XNOR2_X1 U387 ( .A(n392), .B(KEYINPUT32), .ZN(n342) );
  INV_X1 U388 ( .A(n552), .ZN(n343) );
  XNOR2_X1 U389 ( .A(n392), .B(KEYINPUT32), .ZN(n737) );
  XNOR2_X1 U390 ( .A(n422), .B(n421), .ZN(n530) );
  NOR2_X2 U391 ( .A1(n587), .A2(n685), .ZN(n585) );
  XNOR2_X2 U392 ( .A(n465), .B(n464), .ZN(n401) );
  OR2_X1 U393 ( .A1(n710), .A2(G902), .ZN(n370) );
  XNOR2_X1 U394 ( .A(n556), .B(n557), .ZN(n561) );
  XNOR2_X1 U395 ( .A(n562), .B(n446), .ZN(n445) );
  INV_X1 U396 ( .A(KEYINPUT30), .ZN(n446) );
  XNOR2_X1 U397 ( .A(n512), .B(n371), .ZN(n724) );
  INV_X1 U398 ( .A(n475), .ZN(n371) );
  XNOR2_X1 U399 ( .A(n477), .B(n476), .ZN(n521) );
  INV_X1 U400 ( .A(KEYINPUT8), .ZN(n476) );
  NAND2_X1 U401 ( .A1(n726), .A2(G234), .ZN(n477) );
  NAND2_X1 U402 ( .A1(n530), .A2(n529), .ZN(n394) );
  AND2_X1 U403 ( .A1(n582), .A2(n433), .ZN(n529) );
  NOR2_X1 U404 ( .A1(n390), .A2(n405), .ZN(n361) );
  XNOR2_X1 U405 ( .A(n416), .B(KEYINPUT20), .ZN(n485) );
  NAND2_X1 U406 ( .A1(n601), .A2(G234), .ZN(n416) );
  XNOR2_X1 U407 ( .A(n386), .B(n385), .ZN(n566) );
  INV_X1 U408 ( .A(KEYINPUT78), .ZN(n385) );
  OR2_X1 U409 ( .A1(n387), .A2(n559), .ZN(n386) );
  XOR2_X1 U410 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n492) );
  XNOR2_X1 U411 ( .A(G137), .B(G101), .ZN(n491) );
  INV_X1 U412 ( .A(KEYINPUT44), .ZN(n430) );
  XNOR2_X1 U413 ( .A(G140), .B(G137), .ZN(n475) );
  INV_X1 U414 ( .A(KEYINPUT40), .ZN(n412) );
  XNOR2_X1 U415 ( .A(n366), .B(n384), .ZN(n365) );
  INV_X1 U416 ( .A(KEYINPUT28), .ZN(n384) );
  OR2_X1 U417 ( .A1(n607), .A2(G902), .ZN(n498) );
  OR2_X1 U418 ( .A1(n615), .A2(G902), .ZN(n414) );
  XNOR2_X1 U419 ( .A(G116), .B(G122), .ZN(n517) );
  XNOR2_X1 U420 ( .A(G134), .B(G107), .ZN(n516) );
  INV_X1 U421 ( .A(G128), .ZN(n451) );
  INV_X1 U422 ( .A(n381), .ZN(n420) );
  NAND2_X1 U423 ( .A1(n440), .A2(n441), .ZN(n598) );
  AND2_X1 U424 ( .A1(n437), .A2(n436), .ZN(n440) );
  NAND2_X1 U425 ( .A1(n381), .A2(n668), .ZN(n571) );
  XNOR2_X1 U426 ( .A(n593), .B(n400), .ZN(n572) );
  INV_X1 U427 ( .A(KEYINPUT111), .ZN(n400) );
  XNOR2_X1 U428 ( .A(n379), .B(G478), .ZN(n543) );
  NAND2_X1 U429 ( .A1(n705), .A2(n524), .ZN(n379) );
  INV_X1 U430 ( .A(G902), .ZN(n524) );
  INV_X1 U431 ( .A(n570), .ZN(n418) );
  XNOR2_X1 U432 ( .A(n372), .B(n724), .ZN(n710) );
  XNOR2_X1 U433 ( .A(n482), .B(n346), .ZN(n372) );
  BUF_X1 U434 ( .A(G953), .Z(n732) );
  XNOR2_X1 U435 ( .A(n569), .B(KEYINPUT68), .ZN(n580) );
  AND2_X1 U436 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U437 ( .A(n373), .B(G146), .ZN(n474) );
  INV_X1 U438 ( .A(G125), .ZN(n373) );
  INV_X1 U439 ( .A(KEYINPUT103), .ZN(n429) );
  XNOR2_X1 U440 ( .A(n474), .B(n425), .ZN(n377) );
  NAND2_X1 U441 ( .A1(n726), .A2(G224), .ZN(n425) );
  XNOR2_X1 U442 ( .A(n424), .B(KEYINPUT18), .ZN(n376) );
  XNOR2_X1 U443 ( .A(KEYINPUT88), .B(KEYINPUT17), .ZN(n424) );
  XNOR2_X1 U444 ( .A(n388), .B(n348), .ZN(n459) );
  XNOR2_X1 U445 ( .A(KEYINPUT89), .B(KEYINPUT14), .ZN(n388) );
  INV_X1 U446 ( .A(n561), .ZN(n393) );
  OR2_X1 U447 ( .A1(G902), .A2(G237), .ZN(n458) );
  NAND2_X1 U448 ( .A1(n434), .A2(n433), .ZN(n654) );
  INV_X1 U449 ( .A(n567), .ZN(n434) );
  XNOR2_X1 U450 ( .A(n367), .B(n497), .ZN(n607) );
  XNOR2_X1 U451 ( .A(G128), .B(G110), .ZN(n480) );
  XNOR2_X1 U452 ( .A(n474), .B(n447), .ZN(n512) );
  INV_X1 U453 ( .A(KEYINPUT10), .ZN(n447) );
  XNOR2_X1 U454 ( .A(G140), .B(KEYINPUT12), .ZN(n504) );
  XOR2_X1 U455 ( .A(KEYINPUT11), .B(KEYINPUT98), .Z(n505) );
  INV_X1 U456 ( .A(KEYINPUT15), .ZN(n456) );
  XNOR2_X1 U457 ( .A(G902), .B(KEYINPUT87), .ZN(n417) );
  XNOR2_X1 U458 ( .A(KEYINPUT91), .B(G104), .ZN(n466) );
  NOR2_X1 U459 ( .A1(n631), .A2(n412), .ZN(n407) );
  NAND2_X1 U460 ( .A1(n631), .A2(n412), .ZN(n410) );
  XNOR2_X1 U461 ( .A(n364), .B(n382), .ZN(n587) );
  INV_X1 U462 ( .A(KEYINPUT109), .ZN(n382) );
  INV_X1 U463 ( .A(n581), .ZN(n383) );
  XNOR2_X1 U464 ( .A(n395), .B(n515), .ZN(n544) );
  OR2_X1 U465 ( .A1(n700), .A2(G902), .ZN(n395) );
  INV_X1 U466 ( .A(KEYINPUT0), .ZN(n421) );
  XOR2_X1 U467 ( .A(n463), .B(KEYINPUT90), .Z(n449) );
  XNOR2_X1 U468 ( .A(n523), .B(n380), .ZN(n705) );
  NAND2_X1 U469 ( .A1(n597), .A2(n420), .ZN(n642) );
  NOR2_X1 U470 ( .A1(n575), .A2(n655), .ZN(n639) );
  NOR2_X1 U471 ( .A1(n655), .A2(n534), .ZN(n531) );
  NOR2_X1 U472 ( .A1(n443), .A2(n442), .ZN(n578) );
  NOR2_X1 U473 ( .A1(n403), .A2(n711), .ZN(n402) );
  NAND2_X1 U474 ( .A1(n709), .A2(G217), .ZN(n404) );
  XNOR2_X1 U475 ( .A(n389), .B(G131), .ZN(G33) );
  XNOR2_X1 U476 ( .A(n638), .B(G116), .ZN(G18) );
  AND2_X1 U477 ( .A1(G210), .A2(n458), .ZN(n344) );
  AND2_X1 U478 ( .A1(n642), .A2(n599), .ZN(n345) );
  XOR2_X1 U479 ( .A(n481), .B(n480), .Z(n346) );
  AND2_X1 U480 ( .A1(n600), .A2(n345), .ZN(n645) );
  INV_X1 U481 ( .A(n651), .ZN(n433) );
  XOR2_X1 U482 ( .A(n484), .B(n483), .Z(n347) );
  AND2_X1 U483 ( .A1(G237), .A2(G234), .ZN(n348) );
  AND2_X1 U484 ( .A1(n445), .A2(n439), .ZN(n349) );
  AND2_X1 U485 ( .A1(n633), .A2(n580), .ZN(n350) );
  NOR2_X1 U486 ( .A1(n532), .A2(n399), .ZN(n351) );
  AND2_X1 U487 ( .A1(n560), .A2(n579), .ZN(n352) );
  AND2_X1 U488 ( .A1(n345), .A2(KEYINPUT2), .ZN(n353) );
  XOR2_X1 U489 ( .A(KEYINPUT72), .B(KEYINPUT22), .Z(n354) );
  XNOR2_X1 U490 ( .A(KEYINPUT76), .B(KEYINPUT19), .ZN(n355) );
  XNOR2_X1 U491 ( .A(KEYINPUT74), .B(KEYINPUT38), .ZN(n356) );
  INV_X1 U492 ( .A(n579), .ZN(n444) );
  XNOR2_X1 U493 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n357) );
  XOR2_X1 U494 ( .A(n695), .B(n694), .Z(n358) );
  NAND2_X1 U495 ( .A1(n359), .A2(n589), .ZN(n415) );
  NAND2_X1 U496 ( .A1(n362), .A2(n360), .ZN(n359) );
  NAND2_X1 U497 ( .A1(n361), .A2(n369), .ZN(n360) );
  NAND2_X1 U498 ( .A1(n363), .A2(n413), .ZN(n362) );
  NAND2_X1 U499 ( .A1(n369), .A2(n389), .ZN(n363) );
  NAND2_X1 U500 ( .A1(n383), .A2(n365), .ZN(n364) );
  NAND2_X1 U501 ( .A1(n399), .A2(n580), .ZN(n366) );
  XNOR2_X1 U502 ( .A(n367), .B(n472), .ZN(n615) );
  XNOR2_X2 U503 ( .A(n401), .B(G146), .ZN(n367) );
  NAND2_X1 U504 ( .A1(n368), .A2(n423), .ZN(n630) );
  INV_X1 U505 ( .A(n587), .ZN(n368) );
  INV_X1 U506 ( .A(n735), .ZN(n369) );
  XNOR2_X2 U507 ( .A(n391), .B(G119), .ZN(n496) );
  XNOR2_X2 U508 ( .A(n378), .B(KEYINPUT4), .ZN(n465) );
  XNOR2_X1 U509 ( .A(n522), .B(n378), .ZN(n380) );
  XNOR2_X2 U510 ( .A(n452), .B(n451), .ZN(n378) );
  INV_X1 U511 ( .A(n633), .ZN(n631) );
  NAND2_X1 U512 ( .A1(n570), .A2(n350), .ZN(n593) );
  AND2_X1 U513 ( .A1(n563), .A2(n381), .ZN(n564) );
  NOR2_X1 U514 ( .A1(n566), .A2(n651), .ZN(n568) );
  NOR2_X1 U515 ( .A1(n558), .A2(G900), .ZN(n387) );
  XNOR2_X1 U516 ( .A(n585), .B(n584), .ZN(n735) );
  INV_X1 U517 ( .A(n409), .ZN(n390) );
  XNOR2_X2 U518 ( .A(G116), .B(KEYINPUT3), .ZN(n391) );
  XNOR2_X2 U519 ( .A(n420), .B(n356), .ZN(n667) );
  XNOR2_X1 U520 ( .A(n555), .B(n429), .ZN(n428) );
  NAND2_X2 U521 ( .A1(n540), .A2(n531), .ZN(n392) );
  NOR2_X1 U522 ( .A1(n711), .A2(n703), .ZN(n704) );
  NAND2_X1 U523 ( .A1(n598), .A2(n412), .ZN(n411) );
  NAND2_X1 U524 ( .A1(n393), .A2(n444), .ZN(n436) );
  NAND2_X1 U525 ( .A1(n532), .A2(n397), .ZN(n502) );
  XNOR2_X1 U526 ( .A(n404), .B(n710), .ZN(n403) );
  NAND2_X1 U527 ( .A1(n423), .A2(n449), .ZN(n422) );
  XNOR2_X2 U528 ( .A(n394), .B(n354), .ZN(n419) );
  XNOR2_X1 U529 ( .A(n510), .B(n448), .ZN(n511) );
  XNOR2_X1 U530 ( .A(n396), .B(n503), .ZN(n526) );
  NAND2_X1 U531 ( .A1(n676), .A2(n343), .ZN(n396) );
  XNOR2_X1 U532 ( .A(n432), .B(KEYINPUT82), .ZN(n431) );
  BUF_X2 U533 ( .A(n660), .Z(n399) );
  NAND2_X1 U534 ( .A1(n521), .A2(G221), .ZN(n479) );
  XNOR2_X1 U535 ( .A(n401), .B(n724), .ZN(n728) );
  XNOR2_X1 U536 ( .A(n402), .B(KEYINPUT124), .ZN(G66) );
  NAND2_X1 U537 ( .A1(n406), .A2(n586), .ZN(n405) );
  INV_X1 U538 ( .A(n598), .ZN(n408) );
  INV_X1 U539 ( .A(n586), .ZN(n413) );
  XNOR2_X2 U540 ( .A(n414), .B(n473), .ZN(n581) );
  NOR2_X2 U541 ( .A1(n590), .A2(n415), .ZN(n591) );
  NAND2_X1 U542 ( .A1(n419), .A2(n351), .ZN(n533) );
  AND2_X2 U543 ( .A1(n419), .A2(n418), .ZN(n540) );
  INV_X1 U544 ( .A(n530), .ZN(n552) );
  XNOR2_X2 U545 ( .A(n581), .B(KEYINPUT1), .ZN(n655) );
  OR2_X2 U546 ( .A1(n603), .A2(KEYINPUT2), .ZN(n604) );
  AND2_X4 U547 ( .A1(n605), .A2(n604), .ZN(n709) );
  NAND2_X1 U548 ( .A1(n426), .A2(n428), .ZN(n427) );
  XNOR2_X1 U549 ( .A(n539), .B(n430), .ZN(n426) );
  NAND2_X1 U550 ( .A1(n600), .A2(n353), .ZN(n432) );
  NOR2_X1 U551 ( .A1(n431), .A2(n644), .ZN(n643) );
  XNOR2_X2 U552 ( .A(n427), .B(n357), .ZN(n644) );
  NAND2_X1 U553 ( .A1(n445), .A2(n435), .ZN(n438) );
  AND2_X1 U554 ( .A1(n667), .A2(n560), .ZN(n435) );
  NAND2_X1 U555 ( .A1(n438), .A2(n444), .ZN(n437) );
  AND2_X1 U556 ( .A1(n667), .A2(n352), .ZN(n439) );
  NAND2_X1 U557 ( .A1(n349), .A2(n561), .ZN(n441) );
  INV_X1 U558 ( .A(n445), .ZN(n442) );
  NAND2_X1 U559 ( .A1(n561), .A2(n560), .ZN(n443) );
  NOR2_X1 U560 ( .A1(n711), .A2(n697), .ZN(n698) );
  NOR2_X1 U561 ( .A1(n572), .A2(n571), .ZN(n574) );
  XNOR2_X1 U562 ( .A(n696), .B(n358), .ZN(n697) );
  NAND2_X1 U563 ( .A1(n709), .A2(G210), .ZN(n696) );
  AND2_X1 U564 ( .A1(n509), .A2(G214), .ZN(n448) );
  INV_X1 U565 ( .A(n641), .ZN(n599) );
  INV_X1 U566 ( .A(n566), .ZN(n560) );
  INV_X1 U567 ( .A(KEYINPUT36), .ZN(n573) );
  BUF_X1 U568 ( .A(n645), .Z(n725) );
  XNOR2_X1 U569 ( .A(n702), .B(n701), .ZN(n703) );
  AND2_X1 U570 ( .A1(n610), .A2(n732), .ZN(n711) );
  XNOR2_X1 U571 ( .A(G104), .B(G113), .ZN(n450) );
  XNOR2_X1 U572 ( .A(n450), .B(G122), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n453), .B(G101), .ZN(n717) );
  INV_X1 U574 ( .A(KEYINPUT69), .ZN(n454) );
  XNOR2_X1 U575 ( .A(n717), .B(n454), .ZN(n471) );
  XOR2_X1 U576 ( .A(n465), .B(n471), .Z(n455) );
  NAND2_X1 U577 ( .A1(n693), .A2(n601), .ZN(n457) );
  NAND2_X1 U578 ( .A1(G214), .A2(n458), .ZN(n668) );
  XOR2_X1 U579 ( .A(KEYINPUT73), .B(n459), .Z(n460) );
  NAND2_X1 U580 ( .A1(G952), .A2(n460), .ZN(n683) );
  NOR2_X1 U581 ( .A1(n732), .A2(n683), .ZN(n559) );
  AND2_X1 U582 ( .A1(n732), .A2(n460), .ZN(n461) );
  NAND2_X1 U583 ( .A1(G902), .A2(n461), .ZN(n558) );
  NOR2_X1 U584 ( .A1(G898), .A2(n558), .ZN(n462) );
  NOR2_X1 U585 ( .A1(n559), .A2(n462), .ZN(n463) );
  XNOR2_X1 U586 ( .A(G134), .B(G131), .ZN(n464) );
  XNOR2_X1 U587 ( .A(n475), .B(n466), .ZN(n469) );
  NAND2_X1 U588 ( .A1(n726), .A2(G227), .ZN(n467) );
  XNOR2_X1 U589 ( .A(n467), .B(KEYINPUT77), .ZN(n468) );
  XNOR2_X1 U590 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U591 ( .A(n471), .B(n470), .ZN(n472) );
  INV_X1 U592 ( .A(G469), .ZN(n473) );
  INV_X1 U593 ( .A(n655), .ZN(n532) );
  XOR2_X1 U594 ( .A(KEYINPUT24), .B(G119), .Z(n478) );
  XNOR2_X1 U595 ( .A(n479), .B(n478), .ZN(n482) );
  XOR2_X1 U596 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n481) );
  NAND2_X1 U597 ( .A1(n485), .A2(G217), .ZN(n484) );
  INV_X1 U598 ( .A(KEYINPUT25), .ZN(n483) );
  XOR2_X1 U599 ( .A(KEYINPUT94), .B(KEYINPUT21), .Z(n487) );
  NAND2_X1 U600 ( .A1(n485), .A2(G221), .ZN(n486) );
  XNOR2_X1 U601 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U602 ( .A(n488), .B(KEYINPUT93), .ZN(n651) );
  INV_X1 U603 ( .A(n654), .ZN(n546) );
  XOR2_X1 U604 ( .A(G113), .B(KEYINPUT95), .Z(n490) );
  NOR2_X1 U605 ( .A1(n732), .A2(G237), .ZN(n509) );
  NAND2_X1 U606 ( .A1(G210), .A2(n509), .ZN(n489) );
  XNOR2_X1 U607 ( .A(n490), .B(n489), .ZN(n494) );
  XNOR2_X1 U608 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U609 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U610 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X2 U611 ( .A(n498), .B(G472), .ZN(n660) );
  INV_X1 U612 ( .A(KEYINPUT102), .ZN(n499) );
  XNOR2_X1 U613 ( .A(n499), .B(KEYINPUT6), .ZN(n500) );
  XNOR2_X1 U614 ( .A(n660), .B(n500), .ZN(n570) );
  XNOR2_X1 U615 ( .A(KEYINPUT104), .B(KEYINPUT33), .ZN(n501) );
  XNOR2_X1 U616 ( .A(n502), .B(n501), .ZN(n676) );
  XNOR2_X1 U617 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n503) );
  XNOR2_X1 U618 ( .A(KEYINPUT13), .B(G475), .ZN(n515) );
  XNOR2_X1 U619 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U620 ( .A(n506), .B(KEYINPUT99), .Z(n508) );
  XNOR2_X1 U621 ( .A(G143), .B(G131), .ZN(n507) );
  XNOR2_X1 U622 ( .A(n508), .B(n507), .ZN(n514) );
  XNOR2_X1 U623 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U624 ( .A(n514), .B(n513), .Z(n700) );
  INV_X1 U625 ( .A(n544), .ZN(n528) );
  XNOR2_X1 U626 ( .A(n516), .B(KEYINPUT100), .ZN(n520) );
  XOR2_X1 U627 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n518) );
  XNOR2_X1 U628 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U629 ( .A(n520), .B(n519), .Z(n523) );
  NAND2_X1 U630 ( .A1(G217), .A2(n521), .ZN(n522) );
  NAND2_X1 U631 ( .A1(n528), .A2(n543), .ZN(n525) );
  XNOR2_X1 U632 ( .A(n525), .B(KEYINPUT105), .ZN(n563) );
  NAND2_X1 U633 ( .A1(n526), .A2(n563), .ZN(n527) );
  XNOR2_X1 U634 ( .A(n537), .B(G122), .ZN(G24) );
  INV_X1 U635 ( .A(n567), .ZN(n534) );
  XNOR2_X1 U636 ( .A(n533), .B(KEYINPUT67), .ZN(n535) );
  INV_X1 U637 ( .A(n534), .ZN(n650) );
  NAND2_X1 U638 ( .A1(n535), .A2(n650), .ZN(n625) );
  NAND2_X1 U639 ( .A1(n737), .A2(n625), .ZN(n536) );
  XNOR2_X1 U640 ( .A(n536), .B(KEYINPUT85), .ZN(n538) );
  NAND2_X1 U641 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U642 ( .A1(n540), .A2(n655), .ZN(n541) );
  XNOR2_X1 U643 ( .A(n541), .B(KEYINPUT84), .ZN(n542) );
  NOR2_X1 U644 ( .A1(n542), .A2(n650), .ZN(n619) );
  NAND2_X1 U645 ( .A1(n544), .A2(n543), .ZN(n626) );
  INV_X1 U646 ( .A(n626), .ZN(n636) );
  NOR2_X1 U647 ( .A1(n633), .A2(n636), .ZN(n545) );
  XOR2_X1 U648 ( .A(KEYINPUT101), .B(n545), .Z(n673) );
  XOR2_X1 U649 ( .A(KEYINPUT97), .B(KEYINPUT31), .Z(n549) );
  NAND2_X1 U650 ( .A1(n546), .A2(n399), .ZN(n547) );
  NOR2_X1 U651 ( .A1(n655), .A2(n547), .ZN(n662) );
  NAND2_X1 U652 ( .A1(n343), .A2(n662), .ZN(n548) );
  XNOR2_X1 U653 ( .A(n549), .B(n548), .ZN(n637) );
  INV_X1 U654 ( .A(n399), .ZN(n550) );
  NAND2_X1 U655 ( .A1(n556), .A2(n550), .ZN(n551) );
  NOR2_X1 U656 ( .A1(n552), .A2(n551), .ZN(n621) );
  NOR2_X1 U657 ( .A1(n637), .A2(n621), .ZN(n553) );
  NOR2_X1 U658 ( .A1(n673), .A2(n553), .ZN(n554) );
  NOR2_X1 U659 ( .A1(n619), .A2(n554), .ZN(n555) );
  INV_X1 U660 ( .A(KEYINPUT107), .ZN(n557) );
  NAND2_X1 U661 ( .A1(n660), .A2(n668), .ZN(n562) );
  NAND2_X1 U662 ( .A1(n578), .A2(n564), .ZN(n565) );
  XNOR2_X1 U663 ( .A(KEYINPUT108), .B(n565), .ZN(n739) );
  XOR2_X1 U664 ( .A(n739), .B(KEYINPUT81), .Z(n577) );
  XNOR2_X1 U665 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U666 ( .A(n639), .B(KEYINPUT83), .ZN(n576) );
  NAND2_X1 U667 ( .A1(n577), .A2(n576), .ZN(n590) );
  XNOR2_X1 U668 ( .A(KEYINPUT70), .B(KEYINPUT39), .ZN(n579) );
  NAND2_X1 U669 ( .A1(n668), .A2(n667), .ZN(n672) );
  INV_X1 U670 ( .A(n582), .ZN(n671) );
  XNOR2_X1 U671 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n584) );
  XNOR2_X1 U672 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n586) );
  NOR2_X1 U673 ( .A1(n673), .A2(n630), .ZN(n588) );
  XNOR2_X1 U674 ( .A(n588), .B(KEYINPUT47), .ZN(n589) );
  XNOR2_X1 U675 ( .A(n591), .B(KEYINPUT48), .ZN(n600) );
  INV_X1 U676 ( .A(n668), .ZN(n592) );
  NOR2_X1 U677 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U678 ( .A1(n594), .A2(n655), .ZN(n595) );
  XNOR2_X1 U679 ( .A(n595), .B(KEYINPUT43), .ZN(n596) );
  XNOR2_X1 U680 ( .A(n596), .B(KEYINPUT106), .ZN(n597) );
  NOR2_X1 U681 ( .A1(n598), .A2(n626), .ZN(n641) );
  NOR2_X2 U682 ( .A1(n643), .A2(n601), .ZN(n605) );
  XNOR2_X1 U683 ( .A(n645), .B(KEYINPUT75), .ZN(n602) );
  NOR2_X1 U684 ( .A1(n644), .A2(n602), .ZN(n603) );
  NAND2_X1 U685 ( .A1(n709), .A2(G472), .ZN(n609) );
  XNOR2_X1 U686 ( .A(KEYINPUT112), .B(KEYINPUT62), .ZN(n606) );
  XNOR2_X1 U687 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U688 ( .A(n609), .B(n608), .ZN(n611) );
  INV_X1 U689 ( .A(G952), .ZN(n610) );
  NOR2_X1 U690 ( .A1(n611), .A2(n711), .ZN(n613) );
  XNOR2_X1 U691 ( .A(KEYINPUT113), .B(KEYINPUT63), .ZN(n612) );
  XNOR2_X1 U692 ( .A(n613), .B(n612), .ZN(G57) );
  NAND2_X1 U693 ( .A1(n709), .A2(G469), .ZN(n617) );
  XOR2_X1 U694 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n614) );
  XNOR2_X1 U695 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U696 ( .A(n617), .B(n616), .ZN(n618) );
  NOR2_X1 U697 ( .A1(n618), .A2(n711), .ZN(G54) );
  XOR2_X1 U698 ( .A(G101), .B(n619), .Z(G3) );
  NAND2_X1 U699 ( .A1(n621), .A2(n633), .ZN(n620) );
  XNOR2_X1 U700 ( .A(n620), .B(G104), .ZN(G6) );
  XOR2_X1 U701 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n623) );
  NAND2_X1 U702 ( .A1(n621), .A2(n636), .ZN(n622) );
  XNOR2_X1 U703 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U704 ( .A(G107), .B(n624), .ZN(G9) );
  XNOR2_X1 U705 ( .A(n625), .B(G110), .ZN(G12) );
  NOR2_X1 U706 ( .A1(n626), .A2(n630), .ZN(n628) );
  XNOR2_X1 U707 ( .A(KEYINPUT29), .B(KEYINPUT114), .ZN(n627) );
  XNOR2_X1 U708 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U709 ( .A(G128), .B(n629), .ZN(G30) );
  NOR2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U711 ( .A(G146), .B(n632), .Z(G48) );
  NAND2_X1 U712 ( .A1(n637), .A2(n633), .ZN(n634) );
  XNOR2_X1 U713 ( .A(n634), .B(KEYINPUT116), .ZN(n635) );
  XNOR2_X1 U714 ( .A(G113), .B(n635), .ZN(G15) );
  NAND2_X1 U715 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U716 ( .A(n639), .B(G125), .ZN(n640) );
  XNOR2_X1 U717 ( .A(n640), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U718 ( .A(G134), .B(n641), .Z(G36) );
  XNOR2_X1 U719 ( .A(G140), .B(n642), .ZN(G42) );
  INV_X1 U720 ( .A(n643), .ZN(n649) );
  INV_X1 U721 ( .A(n644), .ZN(n712) );
  NAND2_X1 U722 ( .A1(n712), .A2(n725), .ZN(n647) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(KEYINPUT80), .Z(n646) );
  NAND2_X1 U724 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n690) );
  NAND2_X1 U726 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U727 ( .A(n652), .B(KEYINPUT117), .ZN(n653) );
  XNOR2_X1 U728 ( .A(KEYINPUT49), .B(n653), .ZN(n659) );
  NAND2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(KEYINPUT50), .ZN(n657) );
  XNOR2_X1 U731 ( .A(KEYINPUT118), .B(n657), .ZN(n658) );
  NAND2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n661) );
  NOR2_X1 U733 ( .A1(n661), .A2(n399), .ZN(n663) );
  NOR2_X1 U734 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U735 ( .A(n664), .B(KEYINPUT51), .ZN(n665) );
  XNOR2_X1 U736 ( .A(KEYINPUT119), .B(n665), .ZN(n666) );
  NOR2_X1 U737 ( .A1(n685), .A2(n666), .ZN(n679) );
  NOR2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U739 ( .A(n669), .B(KEYINPUT120), .ZN(n670) );
  NOR2_X1 U740 ( .A1(n671), .A2(n670), .ZN(n675) );
  NOR2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n677) );
  INV_X1 U743 ( .A(n676), .ZN(n684) );
  NOR2_X1 U744 ( .A1(n677), .A2(n684), .ZN(n678) );
  NOR2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U746 ( .A(n680), .B(KEYINPUT52), .Z(n681) );
  XNOR2_X1 U747 ( .A(KEYINPUT121), .B(n681), .ZN(n682) );
  NOR2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n687) );
  NOR2_X1 U749 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U750 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U751 ( .A(n688), .B(KEYINPUT122), .ZN(n689) );
  NAND2_X1 U752 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U753 ( .A1(n691), .A2(n732), .ZN(n692) );
  XNOR2_X1 U754 ( .A(n692), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U755 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n695) );
  XNOR2_X1 U756 ( .A(n693), .B(KEYINPUT79), .ZN(n694) );
  XNOR2_X1 U757 ( .A(n698), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U758 ( .A1(n709), .A2(G475), .ZN(n702) );
  XOR2_X1 U759 ( .A(KEYINPUT59), .B(KEYINPUT86), .Z(n699) );
  XNOR2_X1 U760 ( .A(n704), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U761 ( .A1(n709), .A2(G478), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n705), .B(KEYINPUT123), .ZN(n706) );
  XNOR2_X1 U763 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U764 ( .A1(n711), .A2(n708), .ZN(G63) );
  NAND2_X1 U765 ( .A1(n712), .A2(n726), .ZN(n716) );
  NAND2_X1 U766 ( .A1(n732), .A2(G224), .ZN(n713) );
  XNOR2_X1 U767 ( .A(KEYINPUT61), .B(n713), .ZN(n714) );
  NAND2_X1 U768 ( .A1(n714), .A2(G898), .ZN(n715) );
  NAND2_X1 U769 ( .A1(n716), .A2(n715), .ZN(n722) );
  XNOR2_X1 U770 ( .A(n718), .B(n717), .ZN(n720) );
  NOR2_X1 U771 ( .A1(n726), .A2(G898), .ZN(n719) );
  NOR2_X1 U772 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U773 ( .A(n722), .B(n721), .ZN(n723) );
  XOR2_X1 U774 ( .A(KEYINPUT125), .B(n723), .Z(G69) );
  XNOR2_X1 U775 ( .A(n725), .B(n728), .ZN(n727) );
  NAND2_X1 U776 ( .A1(n727), .A2(n726), .ZN(n734) );
  XOR2_X1 U777 ( .A(G227), .B(n728), .Z(n729) );
  NAND2_X1 U778 ( .A1(n729), .A2(G900), .ZN(n730) );
  XNOR2_X1 U779 ( .A(KEYINPUT126), .B(n730), .ZN(n731) );
  NAND2_X1 U780 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n734), .A2(n733), .ZN(G72) );
  BUF_X1 U782 ( .A(n735), .Z(n736) );
  XOR2_X1 U783 ( .A(G137), .B(n736), .Z(G39) );
  XOR2_X1 U784 ( .A(n342), .B(G119), .Z(n738) );
  XNOR2_X1 U785 ( .A(KEYINPUT127), .B(n738), .ZN(G21) );
  XOR2_X1 U786 ( .A(G143), .B(n739), .Z(n740) );
  XNOR2_X1 U787 ( .A(KEYINPUT115), .B(n740), .ZN(G45) );
endmodule

