//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911;
  XOR2_X1   g000(.A(KEYINPUT91), .B(G29gat), .Z(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G43gat), .B(G50gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT15), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(G29gat), .A2(G36gat), .ZN(new_n209));
  XOR2_X1   g008(.A(new_n209), .B(KEYINPUT14), .Z(new_n210));
  NAND3_X1  g009(.A1(new_n204), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n206), .A2(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n212), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n214), .A2(new_n208), .A3(new_n204), .A4(new_n210), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n213), .A2(KEYINPUT17), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT17), .B1(new_n213), .B2(new_n215), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(G15gat), .B(G22gat), .Z(new_n219));
  INV_X1    g018(.A(G1gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT93), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  AND2_X1   g022(.A1(KEYINPUT92), .A2(G1gat), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT16), .B1(KEYINPUT92), .B2(G1gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OR3_X1    g025(.A1(new_n223), .A2(KEYINPUT93), .A3(G1gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n222), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G8gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT94), .ZN(new_n230));
  INV_X1    g029(.A(G8gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n221), .A2(new_n226), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(KEYINPUT95), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n218), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n229), .A2(KEYINPUT94), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT94), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n236), .B1(new_n228), .B2(G8gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n233), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n213), .A2(new_n215), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n234), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n241), .B(KEYINPUT13), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n239), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n247), .B1(new_n230), .B2(new_n233), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n247), .B(new_n233), .C1(new_n235), .C2(new_n237), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n246), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n234), .A2(new_n240), .A3(KEYINPUT18), .A4(new_n241), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n244), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT11), .B(G169gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(G197gat), .ZN(new_n255));
  XOR2_X1   g054(.A(G113gat), .B(G141gat), .Z(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT12), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n258), .A3(new_n251), .A4(new_n252), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n261), .A2(KEYINPUT96), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(KEYINPUT96), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G99gat), .A2(G106gat), .ZN(new_n266));
  INV_X1    g065(.A(G85gat), .ZN(new_n267));
  INV_X1    g066(.A(G92gat), .ZN(new_n268));
  AOI22_X1  g067(.A1(KEYINPUT8), .A2(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT7), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n270), .B1(new_n267), .B2(new_n268), .ZN(new_n271));
  NAND3_X1  g070(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(G99gat), .B(G106gat), .Z(new_n274));
  AND2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n273), .A2(new_n274), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G57gat), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT98), .B1(new_n278), .B2(G64gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT98), .ZN(new_n280));
  INV_X1    g079(.A(G64gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n281), .A3(G57gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(G64gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n279), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G71gat), .B(G78gat), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT99), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n286), .A2(new_n287), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n284), .B(new_n285), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT105), .ZN(new_n291));
  AND3_X1   g090(.A1(KEYINPUT97), .A2(G71gat), .A3(G78gat), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT97), .B1(G71gat), .B2(G78gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OR2_X1    g093(.A1(G71gat), .A2(G78gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G57gat), .B(G64gat), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n294), .B(new_n295), .C1(new_n286), .C2(new_n296), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n290), .A2(new_n291), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n291), .B1(new_n290), .B2(new_n297), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n277), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT10), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n273), .B(new_n274), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n290), .A2(new_n297), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(KEYINPUT105), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n277), .A2(KEYINPUT10), .A3(new_n290), .A4(new_n297), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G230gat), .ZN(new_n308));
  INV_X1    g107(.A(G233gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n300), .A2(new_n304), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n310), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G120gat), .B(G148gat), .ZN(new_n316));
  INV_X1    g115(.A(G176gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(G204gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n312), .A2(new_n314), .A3(new_n319), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n265), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT32), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT65), .ZN(new_n327));
  OAI211_X1 g126(.A(G183gat), .B(G190gat), .C1(new_n327), .C2(KEYINPUT24), .ZN(new_n328));
  NAND2_X1  g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT24), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(KEYINPUT65), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G183gat), .ZN(new_n332));
  INV_X1    g131(.A(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n328), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G169gat), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT23), .B1(new_n336), .B2(new_n317), .ZN(new_n337));
  NAND2_X1  g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n336), .A2(new_n317), .A3(KEYINPUT23), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n335), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT25), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT64), .B(G176gat), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(KEYINPUT23), .A3(new_n336), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n346));
  NAND3_X1  g145(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(new_n334), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT25), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n345), .A2(new_n348), .A3(new_n349), .A4(new_n340), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n343), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G127gat), .B(G134gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G120gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G113gat), .ZN(new_n355));
  INV_X1    g154(.A(G113gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G120gat), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT1), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT67), .ZN(new_n360));
  INV_X1    g159(.A(G134gat), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n360), .A2(new_n361), .A3(G127gat), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n362), .B1(new_n360), .B2(new_n352), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n359), .B1(new_n363), .B2(new_n358), .ZN(new_n364));
  OR3_X1    g163(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n338), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT27), .B1(new_n332), .B2(KEYINPUT66), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT66), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT27), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n370), .A3(G183gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n368), .A2(new_n371), .A3(new_n333), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT28), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT27), .B(G183gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n373), .A2(G190gat), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n329), .B(new_n367), .C1(new_n374), .C2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n351), .A2(new_n364), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n364), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n343), .A2(new_n350), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n372), .A2(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n382));
  INV_X1    g181(.A(new_n329), .ZN(new_n383));
  INV_X1    g182(.A(new_n367), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n380), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n379), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n326), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G15gat), .B(G43gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(G71gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(G99gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT68), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n393), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT33), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n389), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n387), .A2(new_n388), .B1(new_n326), .B2(KEYINPUT33), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n397), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT34), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(KEYINPUT69), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  OR3_X1    g201(.A1(new_n387), .A2(new_n388), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(KEYINPUT69), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n404), .B(new_n402), .C1(new_n387), .C2(new_n388), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n399), .B(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(G78gat), .B(G106gat), .Z(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(KEYINPUT31), .ZN(new_n409));
  INV_X1    g208(.A(G50gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G155gat), .B(G162gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(KEYINPUT77), .B(KEYINPUT2), .Z(new_n415));
  XNOR2_X1  g214(.A(G141gat), .B(G148gat), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n416), .ZN(new_n418));
  INV_X1    g217(.A(G155gat), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT2), .B1(new_n419), .B2(KEYINPUT78), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n413), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G211gat), .A2(G218gat), .ZN(new_n423));
  INV_X1    g222(.A(G211gat), .ZN(new_n424));
  INV_X1    g223(.A(G218gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G197gat), .B(G204gat), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT70), .B(KEYINPUT22), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n423), .B(new_n426), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n423), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n423), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n427), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT29), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n422), .B1(new_n434), .B2(KEYINPUT3), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT83), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT3), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n417), .A2(new_n421), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT29), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n430), .A2(new_n433), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n444), .B(new_n422), .C1(new_n434), .C2(KEYINPUT3), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n436), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(G228gat), .A2(G233gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT82), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n435), .A2(new_n443), .A3(G228gat), .A4(G233gat), .ZN(new_n450));
  INV_X1    g249(.A(G22gat), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n451), .B1(new_n449), .B2(new_n450), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n412), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(KEYINPUT84), .B(new_n412), .C1(new_n452), .C2(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n449), .A2(new_n451), .A3(new_n450), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n453), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI211_X1 g261(.A(KEYINPUT85), .B(new_n451), .C1(new_n449), .C2(new_n450), .ZN(new_n463));
  OR3_X1    g262(.A1(new_n462), .A2(new_n412), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n407), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G64gat), .B(G92gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT75), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(G8gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(G36gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT72), .B1(new_n381), .B2(new_n385), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT72), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n378), .A2(new_n472), .A3(new_n343), .A4(new_n350), .ZN(new_n473));
  NAND2_X1  g272(.A1(G226gat), .A2(G233gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT71), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n439), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n471), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  OR3_X1    g277(.A1(new_n381), .A2(new_n385), .A3(new_n475), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT73), .B1(new_n480), .B2(new_n441), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT73), .ZN(new_n482));
  AOI211_X1 g281(.A(new_n482), .B(new_n442), .C1(new_n478), .C2(new_n479), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n475), .B1(new_n471), .B2(new_n473), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n476), .B1(new_n351), .B2(new_n378), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n485), .A2(new_n441), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT74), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT74), .ZN(new_n490));
  NOR4_X1   g289(.A1(new_n481), .A2(new_n483), .A3(new_n487), .A4(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n470), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n480), .A2(new_n441), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n482), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n480), .A2(KEYINPUT73), .A3(new_n441), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n494), .A2(new_n488), .A3(new_n495), .A4(new_n469), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT30), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n497), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n492), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT35), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n422), .A2(KEYINPUT3), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n504), .A2(new_n380), .A3(new_n438), .ZN(new_n505));
  NAND2_X1  g304(.A1(G225gat), .A2(G233gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n417), .A2(new_n421), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n364), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT4), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT4), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(new_n364), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(KEYINPUT80), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT80), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n510), .A2(new_n517), .A3(KEYINPUT4), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n508), .A2(new_n514), .A3(new_n516), .A4(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n422), .B(new_n359), .C1(new_n358), .C2(new_n363), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n510), .ZN(new_n521));
  INV_X1    g320(.A(new_n506), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n509), .A2(new_n364), .A3(new_n512), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n512), .B1(new_n509), .B2(new_n364), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n523), .B(new_n515), .C1(new_n526), .C2(new_n507), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT0), .B(G57gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(G85gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(G1gat), .B(G29gat), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n530), .B(new_n531), .Z(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT6), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n527), .A3(new_n532), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n528), .A2(KEYINPUT6), .A3(new_n533), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n465), .A2(new_n502), .A3(new_n503), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT90), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n399), .B(new_n406), .Z(new_n542));
  NOR3_X1   g341(.A1(new_n462), .A2(new_n463), .A3(new_n412), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n542), .B1(new_n458), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(new_n501), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT90), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n545), .A2(new_n546), .A3(new_n503), .A4(new_n539), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n494), .A2(new_n488), .A3(new_n495), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n490), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n484), .A2(KEYINPUT74), .A3(new_n488), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n469), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT76), .B1(new_n551), .B2(new_n498), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT76), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n492), .A2(new_n553), .A3(new_n499), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n534), .B(KEYINPUT81), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n536), .A2(new_n535), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n538), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n552), .A2(new_n554), .A3(new_n557), .A4(new_n500), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT35), .B1(new_n558), .B2(new_n544), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n547), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n549), .B2(new_n550), .ZN(new_n562));
  XOR2_X1   g361(.A(KEYINPUT87), .B(KEYINPUT37), .Z(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n494), .A2(new_n488), .A3(new_n495), .A4(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT38), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n469), .A2(KEYINPUT38), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n537), .A2(new_n496), .A3(new_n538), .A4(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n469), .A2(KEYINPUT38), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n485), .A2(new_n486), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n561), .B1(new_n571), .B2(new_n441), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n480), .A2(new_n442), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n565), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT88), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT88), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n565), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n569), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n567), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n514), .A2(new_n505), .A3(new_n518), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n522), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n582), .A2(KEYINPUT39), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n520), .A2(new_n510), .A3(new_n506), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(KEYINPUT39), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n532), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT40), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n583), .A2(KEYINPUT40), .A3(new_n532), .A4(new_n585), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n588), .A2(new_n534), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n501), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n459), .A2(new_n464), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n580), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT89), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n407), .B(KEYINPUT36), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n464), .A2(KEYINPUT86), .A3(new_n456), .A4(new_n457), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT86), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(new_n458), .B2(new_n543), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n595), .B1(new_n558), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT89), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n580), .A2(new_n591), .A3(new_n601), .A4(new_n592), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n594), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n325), .B1(new_n560), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT21), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n230), .B(new_n233), .C1(new_n605), .C2(new_n303), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G183gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT102), .B(G211gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT103), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT101), .Z(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT100), .B(KEYINPUT21), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n303), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n614), .B(new_n616), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n611), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n620));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n620), .B(new_n621), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n619), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n218), .A2(new_n302), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n625));
  INV_X1    g424(.A(G232gat), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n625), .A2(new_n626), .A3(new_n309), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n627), .B1(new_n239), .B2(new_n277), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(G190gat), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n629), .A2(G190gat), .ZN(new_n632));
  OR3_X1    g431(.A1(new_n631), .A2(new_n425), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n425), .B1(new_n631), .B2(new_n632), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT104), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT104), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n633), .A2(new_n637), .A3(new_n634), .ZN(new_n638));
  XNOR2_X1  g437(.A(G134gat), .B(G162gat), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n625), .B1(new_n626), .B2(new_n309), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n636), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n638), .A2(new_n641), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n623), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n604), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n557), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(new_n220), .ZN(G1324gat));
  NOR2_X1   g447(.A1(new_n646), .A2(new_n502), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(KEYINPUT42), .Z(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(new_n231), .B2(new_n649), .ZN(G1325gat));
  INV_X1    g452(.A(new_n646), .ZN(new_n654));
  AOI21_X1  g453(.A(G15gat), .B1(new_n654), .B2(new_n542), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n595), .A2(G15gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT106), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n654), .B2(new_n657), .ZN(G1326gat));
  INV_X1    g457(.A(new_n599), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n646), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT43), .B(G22gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1327gat));
  NAND2_X1  g461(.A1(new_n642), .A2(new_n643), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n560), .B2(new_n603), .ZN(new_n664));
  INV_X1    g463(.A(new_n623), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n325), .ZN(new_n666));
  INV_X1    g465(.A(new_n557), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n664), .A2(new_n666), .A3(new_n667), .A4(new_n202), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT45), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT109), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n603), .A2(KEYINPUT107), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n594), .A2(new_n600), .A3(new_n672), .A4(new_n602), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n671), .A2(new_n560), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n644), .A3(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n560), .A2(new_n603), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT44), .B1(new_n677), .B2(new_n663), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n670), .B1(new_n679), .B2(new_n666), .ZN(new_n680));
  INV_X1    g479(.A(new_n666), .ZN(new_n681));
  AOI211_X1 g480(.A(KEYINPUT109), .B(new_n681), .C1(new_n676), .C2(new_n678), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n557), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n669), .B1(new_n684), .B2(new_n202), .ZN(G1328gat));
  OAI21_X1  g484(.A(G36gat), .B1(new_n683), .B2(new_n502), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n664), .A2(new_n666), .A3(new_n203), .A4(new_n501), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT46), .Z(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(G1329gat));
  INV_X1    g488(.A(G43gat), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n664), .A2(new_n666), .A3(new_n690), .A4(new_n542), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT110), .Z(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n679), .A2(new_n666), .ZN(new_n694));
  INV_X1    g493(.A(new_n595), .ZN(new_n695));
  OAI21_X1  g494(.A(G43gat), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n693), .A2(KEYINPUT47), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n595), .B1(new_n680), .B2(new_n682), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G43gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n693), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT111), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n692), .B1(new_n698), .B2(G43gat), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT111), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n703), .A2(new_n704), .A3(KEYINPUT47), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n697), .B1(new_n702), .B2(new_n705), .ZN(G1330gat));
  OAI21_X1  g505(.A(G50gat), .B1(new_n694), .B2(new_n592), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n664), .A2(new_n666), .A3(new_n410), .A4(new_n599), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(KEYINPUT48), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n599), .B1(new_n680), .B2(new_n682), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n710), .A2(KEYINPUT112), .A3(G50gat), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT112), .B1(new_n710), .B2(G50gat), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n708), .B(KEYINPUT113), .Z(new_n713));
  NOR3_X1   g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n709), .B1(new_n714), .B2(KEYINPUT48), .ZN(G1331gat));
  AND3_X1   g514(.A1(new_n674), .A2(new_n645), .A3(new_n265), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n323), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n557), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(new_n278), .ZN(G1332gat));
  NOR2_X1   g518(.A1(new_n717), .A2(new_n502), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT49), .B(G64gat), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n720), .B2(new_n723), .ZN(G1333gat));
  OAI21_X1  g523(.A(G71gat), .B1(new_n717), .B2(new_n695), .ZN(new_n725));
  INV_X1    g524(.A(G71gat), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n716), .A2(new_n726), .A3(new_n323), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n407), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT114), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT114), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n725), .B(new_n730), .C1(new_n407), .C2(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n659), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g534(.A1(new_n665), .A2(new_n264), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n674), .A2(new_n644), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(new_n323), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(new_n267), .A3(new_n667), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n679), .A2(new_n323), .A3(new_n736), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n667), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT115), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n741), .B1(new_n745), .B2(new_n267), .ZN(G1336gat));
  INV_X1    g545(.A(KEYINPUT116), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n739), .A2(new_n268), .A3(new_n323), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n502), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT52), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n748), .A2(new_n502), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n268), .B1(new_n743), .B2(new_n501), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n750), .B(new_n753), .ZN(G1337gat));
  INV_X1    g553(.A(G99gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n755), .A3(new_n542), .ZN(new_n756));
  OAI21_X1  g555(.A(G99gat), .B1(new_n742), .B2(new_n695), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT117), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1338gat));
  INV_X1    g559(.A(G106gat), .ZN(new_n761));
  INV_X1    g560(.A(new_n592), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n740), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n761), .B1(new_n743), .B2(new_n599), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT53), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767));
  OAI21_X1  g566(.A(G106gat), .B1(new_n742), .B2(new_n592), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n763), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(G1339gat));
  INV_X1    g569(.A(new_n323), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n645), .A2(new_n771), .A3(new_n265), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n240), .A2(new_n249), .A3(new_n245), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n773), .A2(KEYINPUT119), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(KEYINPUT119), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n241), .B1(new_n234), .B2(new_n240), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n257), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n778), .B(new_n323), .C1(new_n262), .C2(new_n263), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n305), .A2(new_n310), .A3(new_n306), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n312), .A2(KEYINPUT54), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n307), .A2(new_n782), .A3(new_n311), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n783), .A2(KEYINPUT118), .A3(new_n320), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT118), .B1(new_n783), .B2(new_n320), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(KEYINPUT55), .B(new_n781), .C1(new_n784), .C2(new_n785), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n322), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n779), .B1(new_n265), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n663), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n778), .B1(new_n262), .B2(new_n263), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n663), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n623), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n772), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n667), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n799), .A2(new_n659), .A3(new_n542), .A4(new_n502), .ZN(new_n800));
  OAI21_X1  g599(.A(G113gat), .B1(new_n800), .B2(new_n265), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n798), .A2(new_n501), .A3(new_n544), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n356), .A3(new_n264), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(G1340gat));
  OAI21_X1  g603(.A(G120gat), .B1(new_n800), .B2(new_n771), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n354), .A3(new_n323), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(G1341gat));
  AOI21_X1  g606(.A(G127gat), .B1(new_n802), .B2(new_n665), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n800), .A2(new_n623), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(G127gat), .ZN(G1342gat));
  NAND3_X1  g609(.A1(new_n802), .A2(new_n361), .A3(new_n644), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT56), .Z(new_n812));
  OAI21_X1  g611(.A(G134gat), .B1(new_n800), .B2(new_n663), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1343gat));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n762), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n595), .A2(new_n557), .A3(new_n501), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(G141gat), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n819), .A3(new_n264), .ZN(new_n820));
  XNOR2_X1  g619(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n815), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n772), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n790), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n788), .A2(KEYINPUT121), .A3(new_n322), .A4(new_n789), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n264), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n825), .B1(new_n829), .B2(new_n779), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(new_n825), .A3(new_n779), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n663), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n795), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n665), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI211_X1 g634(.A(KEYINPUT57), .B(new_n599), .C1(new_n824), .C2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n817), .B1(new_n823), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(new_n264), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n820), .B1(new_n838), .B2(new_n819), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g639(.A(G148gat), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n818), .A2(new_n841), .A3(new_n323), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n797), .A2(new_n762), .A3(new_n821), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n829), .A2(new_n825), .A3(new_n779), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n846), .A2(new_n830), .A3(new_n644), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n845), .B1(new_n847), .B2(new_n795), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n833), .A2(KEYINPUT123), .A3(new_n834), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n623), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n659), .B1(new_n850), .B2(new_n772), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n844), .B1(new_n851), .B2(KEYINPUT57), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n323), .A3(new_n816), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n843), .B1(new_n853), .B2(G148gat), .ZN(new_n854));
  AOI211_X1 g653(.A(KEYINPUT59), .B(new_n841), .C1(new_n837), .C2(new_n323), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n842), .B1(new_n854), .B2(new_n855), .ZN(G1345gat));
  XOR2_X1   g655(.A(KEYINPUT78), .B(G155gat), .Z(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n818), .B2(new_n665), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n665), .A2(new_n857), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n837), .B2(new_n859), .ZN(G1346gat));
  AOI21_X1  g659(.A(G162gat), .B1(new_n818), .B2(new_n644), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n644), .A2(G162gat), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n837), .B2(new_n862), .ZN(G1347gat));
  NOR2_X1   g662(.A1(new_n502), .A2(new_n667), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n797), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n865), .A2(new_n465), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n336), .A3(new_n264), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n865), .A2(new_n659), .A3(new_n542), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n264), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n869), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT124), .B1(new_n869), .B2(G169gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(G1348gat));
  AOI21_X1  g671(.A(G176gat), .B1(new_n866), .B2(new_n323), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n771), .A2(new_n344), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n868), .B2(new_n874), .ZN(G1349gat));
  NAND2_X1  g674(.A1(new_n868), .A2(new_n665), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G183gat), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n866), .A2(new_n665), .A3(new_n375), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g679(.A1(new_n866), .A2(new_n333), .A3(new_n644), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n868), .A2(new_n644), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G190gat), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(KEYINPUT61), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(KEYINPUT61), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(G1351gat));
  NAND2_X1  g685(.A1(new_n695), .A2(new_n864), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT125), .ZN(new_n888));
  AND4_X1   g687(.A1(G197gat), .A2(new_n852), .A3(new_n264), .A4(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n815), .A2(new_n887), .ZN(new_n890));
  AOI21_X1  g689(.A(G197gat), .B1(new_n890), .B2(new_n264), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n889), .A2(new_n891), .ZN(G1352gat));
  INV_X1    g691(.A(new_n890), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(G204gat), .A3(new_n771), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT62), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n852), .A2(new_n323), .A3(new_n888), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(G204gat), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1353gat));
  NAND3_X1  g697(.A1(new_n890), .A2(new_n424), .A3(new_n665), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n623), .A2(new_n887), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n852), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT63), .B1(new_n901), .B2(G211gat), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT63), .ZN(new_n903));
  AOI211_X1 g702(.A(new_n903), .B(new_n424), .C1(new_n852), .C2(new_n900), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n899), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(KEYINPUT126), .B(new_n899), .C1(new_n902), .C2(new_n904), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1354gat));
  NAND4_X1  g708(.A1(new_n852), .A2(G218gat), .A3(new_n644), .A4(new_n888), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n425), .B1(new_n893), .B2(new_n663), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(G1355gat));
endmodule


