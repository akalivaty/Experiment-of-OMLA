//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1222, new_n1223, new_n1224, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1275,
    new_n1276, new_n1277;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n204), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(G58), .A2(G68), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n227), .A2(G50), .A3(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n209), .B1(KEYINPUT1), .B2(new_n222), .C1(new_n225), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n230), .A2(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G68), .Z(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n223), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G50), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n204), .B1(new_n226), .B2(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n254), .B(KEYINPUT70), .Z(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT69), .A2(G58), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT8), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n257), .A2(new_n259), .B1(G150), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n252), .B1(new_n255), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G13), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n253), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n251), .B1(new_n203), .B2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n267), .B1(new_n269), .B2(new_n253), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT9), .ZN(new_n272));
  XOR2_X1   g0072(.A(new_n272), .B(KEYINPUT71), .Z(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G222), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n258), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G223), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(G1698), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n279), .B1(new_n217), .B2(new_n283), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n223), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT67), .B1(new_n287), .B2(new_n223), .ZN(new_n290));
  AND2_X1   g0090(.A1(G1), .A2(G13), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT67), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G41), .A2(G45), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(G1), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n290), .A2(new_n294), .A3(G274), .A4(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT68), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(new_n295), .B2(G1), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n203), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n300));
  AND4_X1   g0100(.A1(new_n290), .A2(new_n299), .A3(new_n294), .A4(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G226), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n297), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n289), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G200), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n271), .A2(KEYINPUT9), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n289), .A2(new_n304), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G190), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n274), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT10), .B1(new_n273), .B2(new_n310), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n266), .A2(new_n257), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n269), .B2(new_n257), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT16), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT76), .ZN(new_n319));
  AOI21_X1  g0119(.A(KEYINPUT7), .B1(new_n277), .B2(new_n204), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n282), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n319), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n281), .A2(new_n204), .A3(new_n282), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT7), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n319), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n211), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G58), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(new_n211), .ZN(new_n330));
  OAI21_X1  g0130(.A(G20), .B1(new_n330), .B2(new_n226), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n260), .A2(G159), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n318), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n324), .A2(new_n325), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n321), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n333), .B1(new_n336), .B2(G68), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n252), .B1(new_n337), .B2(KEYINPUT16), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n317), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n303), .A2(G1698), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(G223), .B2(G1698), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n341), .A2(new_n277), .B1(new_n258), .B2(new_n213), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n288), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n343), .A2(new_n297), .ZN(new_n344));
  INV_X1    g0144(.A(G190), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n287), .A2(KEYINPUT67), .A3(new_n223), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n292), .B1(new_n291), .B2(new_n293), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n299), .A2(new_n300), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(G232), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n344), .A2(KEYINPUT77), .A3(new_n345), .A4(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT77), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(new_n343), .A3(new_n297), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n353), .A2(G190), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n351), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n339), .A2(new_n357), .ZN(new_n358));
  XOR2_X1   g0158(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(KEYINPUT78), .A2(KEYINPUT17), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n339), .B2(new_n357), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n317), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT76), .B1(new_n335), .B2(new_n321), .ZN(new_n365));
  OAI21_X1  g0165(.A(G68), .B1(new_n365), .B2(new_n326), .ZN(new_n366));
  INV_X1    g0166(.A(new_n333), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT16), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(G68), .B1(new_n320), .B2(new_n322), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(KEYINPUT16), .A3(new_n367), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n251), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n364), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n353), .A2(G169), .ZN(new_n373));
  INV_X1    g0173(.A(G179), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n373), .B1(new_n374), .B2(new_n353), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n376), .B(KEYINPUT18), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n363), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n308), .A2(G169), .ZN(new_n379));
  AOI211_X1 g0179(.A(new_n271), .B(new_n379), .C1(new_n374), .C2(new_n308), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n297), .B1(new_n302), .B2(new_n218), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n277), .A2(G107), .ZN(new_n383));
  INV_X1    g0183(.A(G1698), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n283), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G232), .ZN(new_n386));
  OAI221_X1 g0186(.A(new_n383), .B1(new_n385), .B2(new_n386), .C1(new_n212), .C2(new_n285), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n382), .B1(new_n288), .B2(new_n387), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n388), .A2(G169), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n268), .A2(G77), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT8), .B(G58), .ZN(new_n391));
  INV_X1    g0191(.A(new_n260), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n391), .A2(new_n392), .B1(new_n204), .B2(new_n217), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT15), .B(G87), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n393), .B1(new_n259), .B2(new_n395), .ZN(new_n396));
  OAI221_X1 g0196(.A(new_n390), .B1(G77), .B2(new_n265), .C1(new_n396), .C2(new_n252), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n389), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n388), .A2(new_n374), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n397), .B1(new_n388), .B2(G190), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n354), .B2(new_n388), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n315), .A2(new_n378), .A3(new_n381), .A4(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n348), .A2(KEYINPUT72), .A3(G274), .A4(new_n296), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n348), .A2(new_n349), .A3(G238), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G97), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n303), .A2(new_n384), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n386), .A2(G1698), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n407), .B1(new_n410), .B2(new_n277), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n288), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT72), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n297), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n405), .A2(new_n406), .A3(new_n412), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT13), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n301), .A2(G238), .B1(new_n288), .B2(new_n411), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT13), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(new_n414), .A4(new_n405), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G169), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(KEYINPUT75), .A3(KEYINPUT14), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT75), .ZN(new_n423));
  INV_X1    g0223(.A(G169), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n416), .B2(new_n419), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT14), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n420), .A2(new_n426), .A3(G169), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n416), .A2(G179), .A3(new_n419), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n268), .A2(G68), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT73), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n259), .A2(G77), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n260), .A2(G50), .B1(G20), .B2(new_n211), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n252), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n438), .A2(KEYINPUT11), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n266), .A2(new_n211), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT12), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(KEYINPUT11), .ZN(new_n442));
  AND4_X1   g0242(.A1(new_n435), .A2(new_n439), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n433), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT74), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n416), .A2(G190), .A3(new_n419), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n354), .B1(new_n416), .B2(new_n419), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n449), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(KEYINPUT74), .A3(new_n447), .A4(new_n443), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n445), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n404), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G294), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n385), .A2(new_n214), .B1(new_n258), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n283), .A2(G257), .A3(G1698), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n288), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G41), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT5), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n203), .B(G45), .C1(new_n461), .C2(KEYINPUT5), .ZN(new_n464));
  OR2_X1    g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n348), .A2(new_n465), .A3(G264), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT79), .ZN(new_n467));
  OR2_X1    g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n464), .A2(new_n467), .B1(KEYINPUT5), .B2(new_n461), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n348), .A2(G274), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n460), .A2(G179), .A3(new_n466), .A4(new_n470), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n471), .A2(KEYINPUT85), .ZN(new_n472));
  INV_X1    g0272(.A(new_n288), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n278), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(new_n458), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n466), .ZN(new_n476));
  OAI21_X1  g0276(.A(G169), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(KEYINPUT85), .A3(new_n471), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT23), .B1(new_n204), .B2(G107), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT23), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(new_n219), .A3(G20), .ZN(new_n481));
  INV_X1    g0281(.A(G116), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n204), .A2(G33), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n479), .B(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n484), .B(KEYINPUT84), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n283), .A2(new_n204), .A3(G87), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT22), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT22), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n283), .A2(new_n488), .A3(new_n204), .A4(G87), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT24), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT24), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n485), .A2(new_n493), .A3(new_n490), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n252), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n219), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT25), .B1(new_n266), .B2(new_n219), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n252), .B(new_n265), .C1(G1), .C2(new_n258), .ZN(new_n499));
  OAI22_X1  g0299(.A1(new_n497), .A2(new_n498), .B1(new_n499), .B2(new_n219), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n472), .B(new_n478), .C1(new_n495), .C2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT86), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n494), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n493), .B1(new_n485), .B2(new_n490), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n251), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n500), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n508), .A2(KEYINPUT86), .A3(new_n478), .A4(new_n472), .ZN(new_n509));
  INV_X1    g0309(.A(new_n476), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n460), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G200), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(G190), .A3(new_n460), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n506), .A2(new_n512), .A3(new_n507), .A4(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n503), .A2(new_n509), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n283), .A2(G257), .A3(new_n384), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n277), .A2(G303), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n516), .B(new_n517), .C1(new_n285), .C2(new_n220), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n288), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n348), .A2(new_n465), .A3(G270), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n519), .A2(new_n470), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G179), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT21), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n519), .A2(new_n470), .A3(new_n520), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G169), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n522), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G283), .ZN(new_n527));
  INV_X1    g0327(.A(G97), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(new_n204), .C1(G33), .C2(new_n528), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n529), .B(KEYINPUT81), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT20), .ZN(new_n531));
  AOI22_X1  g0331(.A1(KEYINPUT82), .A2(new_n531), .B1(new_n482), .B2(G20), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n251), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n531), .A2(KEYINPUT82), .ZN(new_n534));
  OR3_X1    g0334(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n499), .A2(G116), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(G116), .B2(new_n266), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n534), .B1(new_n530), .B2(new_n533), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n535), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n526), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n539), .B1(G200), .B2(new_n524), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n345), .B2(new_n524), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT83), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n535), .A2(new_n537), .A3(new_n538), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n523), .C1(new_n544), .C2(new_n525), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n539), .A2(G169), .A3(new_n524), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n547), .B2(new_n523), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n540), .B(new_n542), .C1(new_n546), .C2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n283), .A2(G244), .A3(new_n384), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT4), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n283), .A2(G250), .A3(G1698), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n550), .A2(new_n553), .A3(new_n527), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n288), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n348), .A2(new_n465), .A3(G257), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n470), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n424), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n219), .B1(new_n323), .B2(new_n327), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n219), .A2(KEYINPUT6), .A3(G97), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n528), .A2(new_n219), .ZN(new_n562));
  NOR2_X1   g0362(.A1(G97), .A2(G107), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n561), .B1(new_n564), .B2(KEYINPUT6), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G20), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n217), .B2(new_n392), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n251), .B1(new_n560), .B2(new_n567), .ZN(new_n568));
  MUX2_X1   g0368(.A(new_n265), .B(new_n499), .S(G97), .Z(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n559), .B(new_n570), .C1(G179), .C2(new_n558), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n558), .A2(G200), .ZN(new_n572));
  INV_X1    g0372(.A(new_n557), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n555), .B2(new_n288), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(G190), .A3(new_n470), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n572), .A2(new_n575), .A3(new_n568), .A4(new_n569), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n283), .A2(G238), .A3(new_n384), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G116), .ZN(new_n578));
  OAI211_X1 g0378(.A(G244), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n288), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n203), .A2(G45), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n214), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n348), .B(new_n583), .C1(G274), .C2(new_n582), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(new_n345), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(G200), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT19), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n259), .A2(new_n589), .A3(G97), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n563), .A2(new_n213), .B1(new_n407), .B2(new_n204), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(new_n589), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n283), .A2(KEYINPUT80), .A3(new_n204), .A4(G68), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n204), .B(G68), .C1(new_n275), .C2(new_n276), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT80), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n592), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n597), .A2(new_n251), .B1(new_n266), .B2(new_n394), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n499), .A2(new_n213), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n587), .A2(new_n588), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n581), .A2(new_n584), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n374), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n598), .B1(new_n394), .B2(new_n499), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n585), .A2(new_n424), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n571), .A2(new_n576), .A3(new_n600), .A4(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n549), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n455), .A2(new_n515), .A3(new_n607), .ZN(G372));
  INV_X1    g0408(.A(new_n400), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n453), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n363), .B1(new_n610), .B2(new_n445), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n315), .B1(new_n611), .B2(new_n377), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n612), .A2(new_n381), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT26), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT87), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n598), .A2(new_n599), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n354), .B1(new_n581), .B2(new_n584), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n588), .A2(KEYINPUT87), .A3(new_n598), .A4(new_n599), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n619), .A3(new_n587), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n605), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n614), .B1(new_n621), .B2(new_n571), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT88), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n600), .A2(new_n605), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n624), .A2(new_n571), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT26), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT88), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n627), .B(new_n614), .C1(new_n621), .C2(new_n571), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n623), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n605), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n547), .A2(new_n523), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT83), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n545), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(new_n501), .A3(new_n540), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n571), .A2(new_n576), .A3(new_n514), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n621), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n630), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n629), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n455), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n613), .A2(new_n639), .ZN(G369));
  NAND2_X1  g0440(.A1(new_n633), .A2(new_n540), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n264), .A2(new_n204), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(G213), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n544), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(KEYINPUT89), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n650), .A2(KEYINPUT89), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n549), .A2(new_n649), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G330), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n508), .A2(new_n647), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n515), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n501), .A2(new_n648), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT90), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n647), .B1(new_n633), .B2(new_n540), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n501), .A2(new_n647), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n662), .A2(new_n666), .ZN(G399));
  INV_X1    g0467(.A(new_n207), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G41), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G1), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n563), .A2(new_n213), .A3(new_n482), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n671), .A2(new_n672), .B1(new_n229), .B2(new_n670), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT91), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT28), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT26), .B1(new_n621), .B2(new_n571), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n630), .B1(new_n625), .B2(new_n614), .ZN(new_n677));
  AND4_X1   g0477(.A1(new_n503), .A2(new_n633), .A3(new_n509), .A4(new_n540), .ZN(new_n678));
  INV_X1    g0478(.A(new_n636), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n676), .B(new_n677), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(KEYINPUT29), .A3(new_n648), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n647), .B1(new_n629), .B2(new_n637), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n681), .B1(KEYINPUT29), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G330), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n511), .A2(new_n585), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n524), .A2(new_n374), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n685), .A2(KEYINPUT30), .A3(new_n686), .A4(new_n574), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n574), .A2(new_n460), .A3(new_n510), .A4(new_n601), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n689), .B2(new_n522), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n521), .A2(new_n601), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(new_n374), .A3(new_n511), .A4(new_n558), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n687), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(KEYINPUT31), .B1(new_n693), .B2(new_n647), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n647), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n607), .A2(new_n515), .A3(new_n648), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n684), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n683), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n675), .B1(new_n702), .B2(G1), .ZN(G364));
  NOR2_X1   g0503(.A1(new_n263), .A2(G20), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n203), .B1(new_n704), .B2(G45), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n669), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n655), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n654), .A2(G330), .ZN(new_n710));
  NOR2_X1   g0510(.A1(G13), .A2(G33), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G20), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n654), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(G179), .A2(G200), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(G20), .A3(new_n345), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n718), .A2(KEYINPUT95), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(KEYINPUT95), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR4_X1   g0522(.A1(new_n204), .A2(new_n354), .A3(G179), .A4(G190), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n723), .A2(KEYINPUT93), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(KEYINPUT93), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI22_X1  g0527(.A1(G329), .A2(new_n722), .B1(new_n727), .B2(G283), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n204), .A2(new_n374), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n345), .A3(new_n354), .ZN(new_n730));
  INV_X1    g0530(.A(G311), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n204), .A2(new_n345), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(new_n374), .A3(G200), .ZN(new_n734));
  INV_X1    g0534(.A(G303), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n277), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n733), .A2(G179), .A3(new_n354), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n732), .B(new_n736), .C1(G322), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n729), .A2(G200), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G190), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(KEYINPUT33), .B(G317), .Z(new_n743));
  OAI211_X1 g0543(.A(new_n728), .B(new_n739), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n740), .A2(new_n345), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n204), .B1(new_n716), .B2(G190), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n745), .A2(G326), .B1(G294), .B2(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT94), .Z(new_n749));
  NAND2_X1  g0549(.A1(new_n747), .A2(G97), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n718), .A2(G159), .ZN(new_n751));
  INV_X1    g0551(.A(new_n745), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n750), .B1(new_n751), .B2(KEYINPUT32), .C1(new_n752), .C2(new_n253), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n727), .A2(G107), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n737), .B(KEYINPUT92), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G58), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n283), .B1(new_n730), .B2(new_n217), .ZN(new_n758));
  INV_X1    g0558(.A(new_n734), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n758), .B1(G87), .B2(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(KEYINPUT32), .A2(new_n751), .B1(new_n741), .B2(G68), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n754), .A2(new_n757), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n744), .A2(new_n749), .B1(new_n753), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n223), .B1(G20), .B2(new_n424), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n668), .A2(new_n277), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n766), .A2(G355), .B1(new_n482), .B2(new_n668), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n668), .A2(new_n283), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G45), .B2(new_n229), .ZN(new_n769));
  INV_X1    g0569(.A(G45), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n248), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n767), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n713), .A2(new_n764), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n708), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n765), .A2(new_n774), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n709), .A2(new_n710), .B1(new_n715), .B2(new_n775), .ZN(G396));
  NOR2_X1   g0576(.A1(new_n400), .A2(new_n647), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n397), .A2(new_n647), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n402), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n777), .B1(new_n400), .B2(new_n779), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n682), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n638), .A2(new_n648), .A3(new_n780), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n707), .B1(new_n783), .B2(new_n700), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n700), .B2(new_n783), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n764), .A2(new_n711), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n708), .B1(new_n217), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n764), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n727), .A2(G68), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n283), .B1(new_n734), .B2(new_n253), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(G58), .B2(new_n747), .ZN(new_n791));
  INV_X1    g0591(.A(G132), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n789), .B(new_n791), .C1(new_n792), .C2(new_n721), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT34), .ZN(new_n794));
  INV_X1    g0594(.A(new_n730), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G137), .A2(new_n745), .B1(new_n795), .B2(G159), .ZN(new_n796));
  INV_X1    g0596(.A(G150), .ZN(new_n797));
  INV_X1    g0597(.A(G143), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n796), .B1(new_n797), .B2(new_n742), .C1(new_n755), .C2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n793), .B1(new_n794), .B2(new_n799), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n799), .A2(new_n794), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n283), .B1(new_n795), .B2(G116), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n802), .B1(new_n219), .B2(new_n734), .C1(new_n456), .C2(new_n737), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n721), .A2(new_n731), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n726), .A2(new_n213), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n750), .B1(new_n752), .B2(new_n735), .ZN(new_n806));
  NOR4_X1   g0606(.A1(new_n803), .A2(new_n804), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n741), .A2(KEYINPUT96), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n741), .A2(KEYINPUT96), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G283), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n800), .A2(new_n801), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n787), .B1(new_n788), .B2(new_n813), .C1(new_n780), .C2(new_n712), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n785), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G384));
  AOI211_X1 g0616(.A(new_n482), .B(new_n225), .C1(new_n565), .C2(KEYINPUT35), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(KEYINPUT35), .B2(new_n565), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT36), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n229), .A2(new_n217), .A3(new_n330), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n253), .B2(G68), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n821), .A2(new_n203), .A3(G13), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT97), .Z(new_n823));
  INV_X1    g0623(.A(KEYINPUT100), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n777), .B1(new_n682), .B2(new_n780), .ZN(new_n825));
  INV_X1    g0625(.A(new_n645), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n337), .A2(KEYINPUT16), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n364), .B1(new_n371), .B2(new_n827), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n826), .B(new_n828), .C1(new_n363), .C2(new_n377), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n645), .B(KEYINPUT99), .Z(new_n830));
  NAND2_X1  g0630(.A1(new_n372), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT37), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n358), .A2(new_n376), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n828), .B1(new_n375), .B2(new_n826), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n358), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n833), .B1(new_n835), .B2(new_n832), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n829), .A2(KEYINPUT38), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT38), .B1(new_n829), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n443), .A2(new_n648), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n450), .A2(new_n452), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n841), .B2(new_n433), .ZN(new_n842));
  INV_X1    g0642(.A(new_n840), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n431), .B1(new_n427), .B2(new_n422), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n453), .B(new_n843), .C1(new_n844), .C2(new_n443), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n842), .A2(KEYINPUT98), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT98), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n445), .A2(new_n847), .A3(new_n453), .A4(new_n843), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n825), .A2(new_n839), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n377), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n830), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n824), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n777), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n782), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n837), .A2(new_n838), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n846), .A2(new_n848), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n852), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(KEYINPUT100), .A3(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT39), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n839), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n358), .A2(new_n376), .A3(new_n831), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT37), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT101), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(new_n866), .A3(new_n833), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n864), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(KEYINPUT102), .A3(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n372), .B(new_n830), .C1(new_n363), .C2(new_n377), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT102), .B1(new_n867), .B2(new_n868), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n863), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT103), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT103), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n875), .B(new_n863), .C1(new_n871), .C2(new_n872), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n862), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n445), .A2(new_n647), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n853), .B(new_n860), .C1(new_n879), .C2(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n455), .B(new_n681), .C1(KEYINPUT29), .C2(new_n682), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n883), .A2(new_n613), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n882), .B(new_n884), .Z(new_n885));
  INV_X1    g0685(.A(KEYINPUT104), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n693), .A2(new_n886), .A3(KEYINPUT31), .A4(new_n647), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n696), .B1(new_n694), .B2(KEYINPUT104), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n698), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n780), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n849), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT40), .B1(new_n891), .B2(new_n856), .ZN(new_n892));
  INV_X1    g0692(.A(new_n837), .ZN(new_n893));
  INV_X1    g0693(.A(new_n876), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n867), .A2(new_n868), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT102), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(new_n870), .A3(new_n869), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n875), .B1(new_n898), .B2(new_n863), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n893), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n857), .A2(new_n780), .A3(new_n889), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n892), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n455), .A2(new_n889), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n684), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n905), .B2(new_n904), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n885), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n203), .B2(new_n704), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n885), .A2(new_n907), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n819), .B(new_n823), .C1(new_n909), .C2(new_n910), .ZN(G367));
  OR2_X1    g0711(.A1(new_n571), .A2(new_n648), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n570), .A2(new_n647), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n571), .A2(new_n576), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n664), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n916), .A2(KEYINPUT42), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n503), .A2(new_n509), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n918), .A2(new_n914), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n647), .B1(new_n919), .B2(new_n571), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n916), .B2(KEYINPUT42), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n616), .A2(new_n647), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n620), .A2(new_n605), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n605), .B2(new_n923), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT105), .Z(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n929), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n922), .A2(new_n931), .A3(new_n926), .ZN(new_n932));
  INV_X1    g0732(.A(new_n662), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n930), .A2(new_n932), .B1(new_n933), .B2(new_n915), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n922), .A2(new_n931), .A3(new_n926), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n931), .B1(new_n922), .B2(new_n926), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n933), .A2(new_n915), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n669), .B(KEYINPUT41), .Z(new_n940));
  INV_X1    g0740(.A(KEYINPUT44), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n666), .B2(new_n915), .ZN(new_n942));
  INV_X1    g0742(.A(new_n915), .ZN(new_n943));
  OAI211_X1 g0743(.A(KEYINPUT44), .B(new_n943), .C1(new_n664), .C2(new_n665), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n661), .A2(new_n663), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n946), .B(new_n915), .C1(new_n501), .C2(new_n647), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT45), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n933), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n661), .A2(new_n663), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n946), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(new_n655), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(new_n701), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n945), .A2(new_n949), .A3(new_n662), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n951), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n940), .B1(new_n957), .B2(new_n702), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n939), .B1(new_n958), .B2(new_n706), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT106), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT106), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n939), .B(new_n961), .C1(new_n958), .C2(new_n706), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n773), .B1(new_n207), .B2(new_n394), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n768), .B2(new_n241), .ZN(new_n965));
  INV_X1    g0765(.A(G283), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n277), .B1(new_n730), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G317), .B2(new_n718), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n755), .B2(new_n735), .C1(new_n528), .C2(new_n726), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n734), .A2(new_n482), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(KEYINPUT46), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G311), .B2(new_n745), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n970), .A2(KEYINPUT46), .B1(G107), .B2(new_n747), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(new_n456), .C2(new_n810), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n727), .A2(G77), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n746), .A2(new_n211), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n283), .B1(new_n734), .B2(new_n329), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n976), .B(new_n977), .C1(G143), .C2(new_n745), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n737), .A2(new_n797), .B1(new_n730), .B2(new_n253), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G137), .B2(new_n718), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n975), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(G159), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n810), .A2(new_n982), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n969), .A2(new_n974), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT47), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n708), .B(new_n965), .C1(new_n985), .C2(new_n764), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n925), .B2(new_n714), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n963), .A2(new_n987), .ZN(G387));
  NAND2_X1  g0788(.A1(new_n766), .A2(new_n672), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(G107), .B2(new_n207), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n238), .A2(G45), .ZN(new_n991));
  INV_X1    g0791(.A(new_n768), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n391), .A2(G50), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT50), .ZN(new_n994));
  AOI211_X1 g0794(.A(G45), .B(new_n672), .C1(G68), .C2(G77), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n990), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT107), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n773), .B1(new_n997), .B2(new_n998), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n707), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n746), .A2(new_n394), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n759), .A2(G77), .B1(G150), .B2(new_n718), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1003), .B(new_n283), .C1(new_n253), .C2(new_n737), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1002), .B(new_n1004), .C1(G159), .C2(new_n745), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n257), .A2(new_n741), .B1(new_n795), .B2(G68), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT108), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1005), .B(new_n1007), .C1(new_n528), .C2(new_n726), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n283), .B1(new_n718), .B2(G326), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n734), .A2(new_n456), .B1(new_n746), .B2(new_n966), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT109), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(KEYINPUT110), .B(G322), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n745), .A2(new_n1013), .B1(new_n795), .B2(G303), .ZN(new_n1014));
  INV_X1    g0814(.A(G317), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1014), .B1(new_n1015), .B2(new_n755), .C1(new_n810), .C2(new_n731), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT48), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1011), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT49), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1009), .B1(new_n482), .B2(new_n726), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1008), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1001), .B1(new_n1023), .B2(new_n764), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n661), .B2(new_n714), .ZN(new_n1025));
  OAI21_X1  g0825(.A(KEYINPUT111), .B1(new_n955), .B2(new_n670), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n954), .A2(new_n701), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n955), .A2(KEYINPUT111), .A3(new_n670), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1025), .B1(new_n705), .B2(new_n954), .C1(new_n1028), .C2(new_n1029), .ZN(G393));
  NAND2_X1  g0830(.A1(new_n956), .A2(KEYINPUT112), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(new_n951), .Z(new_n1032));
  OAI211_X1 g0832(.A(new_n669), .B(new_n957), .C1(new_n1032), .C2(new_n955), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n943), .A2(new_n713), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n773), .B1(new_n528), .B2(new_n207), .C1(new_n992), .C2(new_n245), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n707), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n746), .A2(new_n217), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n283), .B1(new_n734), .B2(new_n211), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n730), .A2(new_n391), .B1(new_n717), .B2(new_n798), .ZN(new_n1039));
  OR4_X1    g0839(.A1(new_n805), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G150), .A2(new_n745), .B1(new_n738), .B2(G159), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT51), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1040), .B(new_n1042), .C1(G50), .C2(new_n811), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1044), .A2(KEYINPUT113), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n752), .A2(new_n1015), .B1(new_n731), .B2(new_n737), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT52), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n811), .A2(G303), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n277), .B1(new_n734), .B2(new_n966), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n730), .A2(new_n456), .B1(new_n1012), .B2(new_n717), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G116), .C2(new_n747), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1047), .A2(new_n754), .A3(new_n1048), .A4(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1044), .A2(KEYINPUT113), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1045), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1036), .B1(new_n1054), .B2(new_n764), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1032), .A2(new_n706), .B1(new_n1034), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1033), .A2(new_n1056), .ZN(G390));
  OAI21_X1  g0857(.A(new_n789), .B1(new_n456), .B2(new_n721), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT118), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n810), .A2(new_n219), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n283), .B1(new_n759), .B2(G87), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n528), .B2(new_n730), .C1(new_n482), .C2(new_n737), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n752), .A2(new_n966), .B1(new_n746), .B2(new_n217), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n811), .A2(G137), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n734), .A2(new_n797), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT53), .ZN(new_n1067));
  INV_X1    g0867(.A(G125), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1067), .B1(new_n253), .B2(new_n726), .C1(new_n1068), .C2(new_n721), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT54), .B(G143), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n283), .B1(new_n730), .B2(new_n1070), .C1(new_n792), .C2(new_n737), .ZN(new_n1071));
  INV_X1    g0871(.A(G128), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n752), .A2(new_n1072), .B1(new_n746), .B2(new_n982), .ZN(new_n1073));
  NOR4_X1   g0873(.A1(new_n1065), .A2(new_n1069), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n764), .B1(new_n1064), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n786), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n707), .B1(new_n257), .B2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT117), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT119), .Z(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n879), .B2(new_n711), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT120), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n878), .B1(new_n894), .B2(new_n899), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n862), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n881), .B1(new_n825), .B2(new_n849), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n849), .A2(KEYINPUT114), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT114), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n846), .A2(new_n1088), .A3(new_n848), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n400), .A2(new_n779), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n680), .A2(new_n648), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n854), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n880), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n900), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1086), .A2(new_n1095), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n890), .A2(new_n684), .A3(new_n849), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n857), .A2(new_n699), .A3(new_n780), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1086), .A2(new_n1095), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n706), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n455), .A2(G330), .A3(new_n889), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n883), .A2(new_n613), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n857), .B1(new_n699), .B2(new_n780), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n855), .B1(new_n1104), .B2(new_n1097), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n889), .A2(G330), .A3(new_n780), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1087), .A2(new_n1106), .A3(new_n1089), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1107), .A2(new_n854), .A3(new_n1092), .A4(new_n1099), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1103), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n879), .A2(new_n1085), .B1(new_n900), .B2(new_n1094), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1097), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1100), .B(new_n1109), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(KEYINPUT115), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT115), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1098), .A2(new_n1114), .A3(new_n1100), .A4(new_n1109), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1109), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n670), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1116), .A2(KEYINPUT116), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT116), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1082), .B(new_n1101), .C1(new_n1120), .C2(new_n1121), .ZN(G378));
  XNOR2_X1  g0922(.A(new_n1103), .B(KEYINPUT123), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1116), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT57), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n315), .A2(new_n381), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n271), .A2(new_n645), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1127), .B(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1130), .B(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n904), .A2(G330), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n902), .B1(new_n901), .B2(new_n839), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n837), .B1(new_n874), .B2(new_n876), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n891), .A2(KEYINPUT40), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1134), .B(G330), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1130), .B(new_n1131), .Z(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1133), .A2(new_n1139), .ZN(new_n1140));
  OR2_X1    g0940(.A1(new_n1140), .A2(new_n882), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT100), .B1(new_n858), .B2(new_n859), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n1143), .B2(new_n880), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1133), .A2(new_n1139), .B1(new_n1144), .B2(new_n860), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1126), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1125), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT124), .B1(new_n1148), .B2(new_n669), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1123), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1132), .B1(new_n904), .B2(G330), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1151), .A2(new_n1152), .A3(new_n882), .ZN(new_n1153));
  OAI21_X1  g0953(.A(KEYINPUT57), .B1(new_n1153), .B2(new_n1145), .ZN(new_n1154));
  OAI211_X1 g0954(.A(KEYINPUT124), .B(new_n669), .C1(new_n1150), .C2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1153), .A2(new_n1145), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1126), .B1(new_n1150), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1149), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1138), .A2(new_n711), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n707), .B1(G50), .B2(new_n1076), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n727), .A2(G58), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT121), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n976), .B1(new_n745), .B2(G116), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n528), .B2(new_n742), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n721), .A2(new_n966), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n277), .A2(new_n461), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n795), .B2(new_n395), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n217), .B2(new_n734), .C1(new_n219), .C2(new_n737), .ZN(new_n1170));
  NOR4_X1   g0970(.A1(new_n1164), .A2(new_n1166), .A3(new_n1167), .A4(new_n1170), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1171), .A2(KEYINPUT58), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n1072), .A2(new_n737), .B1(new_n734), .B2(new_n1070), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT122), .Z(new_n1174));
  AOI22_X1  g0974(.A1(G125), .A2(new_n745), .B1(new_n795), .B2(G137), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n741), .A2(G132), .B1(G150), .B2(new_n747), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n727), .A2(G159), .ZN(new_n1180));
  AOI211_X1 g0980(.A(G33), .B(G41), .C1(new_n718), .C2(G124), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1171), .A2(KEYINPUT58), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1168), .B(new_n253), .C1(G33), .C2(G41), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1172), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1161), .B1(new_n1185), .B2(new_n764), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1160), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1156), .B2(new_n705), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1159), .A2(new_n1189), .ZN(G375));
  OAI21_X1  g0990(.A(new_n707), .B1(G68), .B2(new_n1076), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1090), .A2(new_n712), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n283), .B1(new_n738), .B2(G283), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n528), .B2(new_n734), .C1(new_n219), .C2(new_n730), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1002), .B(new_n1194), .C1(G294), .C2(new_n745), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n811), .A2(G116), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n722), .A2(G303), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1195), .A2(new_n975), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n283), .B1(new_n734), .B2(new_n982), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n752), .A2(new_n792), .B1(new_n746), .B2(new_n253), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(G150), .C2(new_n795), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G128), .A2(new_n722), .B1(new_n756), .B2(G137), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n810), .C2(new_n1070), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1198), .B1(new_n1164), .B2(new_n1203), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1191), .B(new_n1192), .C1(new_n764), .C2(new_n1204), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1205), .B1(new_n1207), .B2(new_n706), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1206), .A2(new_n1103), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1109), .A2(new_n940), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1208), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT125), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(G381));
  INV_X1    g1013(.A(G375), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1215), .A2(new_n1082), .A3(new_n1101), .ZN(new_n1216));
  INV_X1    g1016(.A(G390), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(G393), .A2(G396), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1217), .A2(new_n815), .A3(new_n1212), .A4(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1219), .A2(G387), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1214), .A2(new_n1216), .A3(new_n1220), .ZN(G407));
  NAND2_X1  g1021(.A1(new_n646), .A2(G213), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1214), .A2(new_n1216), .A3(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(G407), .A2(new_n1224), .A3(G213), .ZN(G409));
  INV_X1    g1025(.A(KEYINPUT127), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(G387), .A2(new_n1217), .ZN(new_n1227));
  XOR2_X1   g1027(.A(G393), .B(G396), .Z(new_n1228));
  NAND3_X1  g1028(.A1(new_n963), .A2(G390), .A3(new_n987), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1228), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT61), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G378), .B(new_n1189), .C1(new_n1149), .C2(new_n1158), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT126), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1188), .A2(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(KEYINPUT126), .B(new_n1187), .C1(new_n1156), .C2(new_n705), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1150), .A2(new_n940), .A3(new_n1156), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1216), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1223), .B1(new_n1234), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1209), .B1(new_n1118), .B2(KEYINPUT60), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1206), .A2(KEYINPUT60), .A3(new_n1103), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n669), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1208), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n815), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1245), .A2(G384), .A3(new_n1208), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1223), .A2(G2897), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1249), .B(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1233), .B1(new_n1241), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT62), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1249), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1254), .B1(new_n1241), .B2(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1223), .B(new_n1249), .C1(new_n1234), .C2(new_n1240), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1254), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1232), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1241), .A2(KEYINPUT63), .A3(new_n1255), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1261), .B(new_n1233), .C1(new_n1241), .C2(new_n1252), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1232), .B1(new_n1258), .B2(KEYINPUT63), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1226), .B1(new_n1260), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1253), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1241), .A2(new_n1255), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1266), .A2(new_n1269), .A3(new_n1232), .A4(new_n1261), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1267), .A2(KEYINPUT62), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1271), .A2(new_n1253), .A3(new_n1256), .ZN(new_n1272));
  OAI211_X1 g1072(.A(KEYINPUT127), .B(new_n1270), .C1(new_n1272), .C2(new_n1232), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1265), .A2(new_n1273), .ZN(G405));
  NAND2_X1  g1074(.A1(G375), .A2(new_n1216), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1234), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(new_n1249), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(new_n1232), .ZN(G402));
endmodule


