//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT74), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G902), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n194), .B(KEYINPUT75), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G128), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  OAI22_X1  g015(.A1(new_n198), .A2(new_n199), .B1(new_n197), .B2(G128), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n195), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G119), .B(G128), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT24), .B(G110), .Z(new_n205));
  OAI22_X1  g019(.A1(new_n203), .A2(G110), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n207));
  INV_X1    g021(.A(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(G125), .ZN(new_n210));
  INV_X1    g024(.A(G125), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G140), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g027(.A(G146), .B(new_n209), .C1(new_n213), .C2(new_n207), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n210), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT78), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G125), .B(G140), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT78), .A3(new_n215), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n206), .A2(new_n214), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n203), .A2(G110), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n209), .B1(new_n213), .B2(new_n207), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(KEYINPUT77), .A3(new_n215), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n215), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT77), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n227), .A3(new_n214), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n205), .A2(new_n204), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n223), .A2(new_n225), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G953), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(G221), .A3(G234), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n232), .B(KEYINPUT79), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT22), .B(G137), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n233), .B(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n222), .A2(new_n230), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n235), .B1(new_n222), .B2(new_n230), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n192), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n191), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI221_X1 g055(.A(new_n192), .B1(KEYINPUT80), .B2(KEYINPUT25), .C1(new_n237), .C2(new_n238), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n189), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n188), .A2(new_n192), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n237), .B2(new_n238), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT73), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT31), .ZN(new_n250));
  XOR2_X1   g064(.A(KEYINPUT2), .B(G113), .Z(new_n251));
  XNOR2_X1  g065(.A(G116), .B(G119), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n251), .A2(new_n252), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT11), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(G137), .ZN(new_n259));
  AND2_X1   g073(.A1(KEYINPUT65), .A2(G134), .ZN(new_n260));
  NOR2_X1   g074(.A1(KEYINPUT65), .A2(G134), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G137), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT11), .A3(G134), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n258), .A2(G137), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n262), .A2(G131), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G131), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n264), .A2(new_n265), .ZN(new_n269));
  OR2_X1    g083(.A1(KEYINPUT65), .A2(G134), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n263), .A2(KEYINPUT11), .ZN(new_n271));
  NAND2_X1  g085(.A1(KEYINPUT65), .A2(G134), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n268), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n257), .B1(new_n267), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(G143), .B(G146), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT0), .B(G128), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n215), .A2(G143), .ZN(new_n279));
  INV_X1    g093(.A(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G146), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n279), .A2(new_n281), .A3(KEYINPUT0), .A4(G128), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT64), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n276), .A2(KEYINPUT64), .A3(KEYINPUT0), .A4(G128), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n278), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G131), .B1(new_n262), .B2(new_n266), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n269), .A2(new_n268), .A3(new_n273), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(KEYINPUT69), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n275), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n276), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT1), .B1(new_n280), .B2(G146), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n293));
  OAI21_X1  g107(.A(G128), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT68), .B1(new_n279), .B2(KEYINPUT1), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT1), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n276), .A2(new_n297), .A3(G128), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n268), .B1(G134), .B2(G137), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n270), .A2(new_n272), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n300), .B1(new_n301), .B2(G137), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n288), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n290), .A2(KEYINPUT30), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n284), .A2(new_n285), .ZN(new_n305));
  INV_X1    g119(.A(new_n278), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n305), .B(new_n306), .C1(new_n267), .C2(new_n274), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT66), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n287), .A2(new_n288), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT66), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n286), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n288), .A2(KEYINPUT67), .A3(new_n302), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n288), .A2(new_n302), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT67), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n313), .A2(new_n314), .B1(new_n296), .B2(new_n298), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n308), .A2(new_n311), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n256), .B(new_n304), .C1(new_n316), .C2(KEYINPUT30), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n290), .A2(KEYINPUT70), .A3(KEYINPUT30), .A4(new_n303), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n255), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n290), .A2(new_n255), .A3(new_n303), .ZN(new_n320));
  NOR2_X1   g134(.A1(G237), .A2(G953), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G210), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT27), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT26), .B(G101), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n250), .B1(new_n319), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n326), .ZN(new_n328));
  INV_X1    g142(.A(new_n318), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n304), .A2(new_n256), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n313), .A2(new_n314), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n312), .A3(new_n299), .ZN(new_n332));
  INV_X1    g146(.A(new_n311), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n310), .B1(new_n309), .B2(new_n286), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT30), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n329), .B1(new_n330), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(KEYINPUT31), .B(new_n328), .C1(new_n338), .C2(new_n255), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n327), .A2(new_n339), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n325), .B(KEYINPUT71), .Z(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT72), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n308), .A2(new_n311), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n255), .B1(new_n344), .B2(new_n332), .ZN(new_n345));
  INV_X1    g159(.A(new_n320), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT28), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n320), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n343), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n255), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n335), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n348), .B1(new_n352), .B2(new_n320), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n353), .A2(KEYINPUT72), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n342), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n340), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(G472), .A2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT32), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n249), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n360), .ZN(new_n362));
  AOI211_X1 g176(.A(KEYINPUT73), .B(new_n362), .C1(new_n340), .C2(new_n355), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT30), .B1(new_n344), .B2(new_n332), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n304), .A2(new_n256), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n318), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n351), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT31), .B1(new_n368), .B2(new_n328), .ZN(new_n369));
  AOI211_X1 g183(.A(new_n250), .B(new_n326), .C1(new_n367), .C2(new_n351), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n349), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT72), .B1(new_n353), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n347), .A2(new_n343), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n341), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n357), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n255), .B1(new_n290), .B2(new_n303), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT28), .B1(new_n346), .B2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n378), .A2(KEYINPUT29), .A3(new_n349), .A4(new_n325), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n192), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n350), .A2(new_n354), .A3(new_n342), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n346), .B1(new_n367), .B2(new_n351), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(new_n325), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n381), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n376), .A2(new_n359), .B1(new_n386), .B2(G472), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n248), .B1(new_n364), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT9), .B(G234), .ZN(new_n389));
  OAI21_X1  g203(.A(G221), .B1(new_n389), .B2(G902), .ZN(new_n390));
  INV_X1    g204(.A(G469), .ZN(new_n391));
  XNOR2_X1  g205(.A(G110), .B(G140), .ZN(new_n392));
  INV_X1    g206(.A(G227), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(G953), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n392), .B(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n299), .ZN(new_n397));
  INV_X1    g211(.A(G107), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G104), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT82), .B(G107), .ZN(new_n400));
  INV_X1    g214(.A(G104), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(KEYINPUT3), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n399), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT3), .B1(new_n401), .B2(G107), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT81), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT81), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n406), .B(KEYINPUT3), .C1(new_n401), .C2(G107), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G101), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n403), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n400), .A2(G104), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n401), .A2(G107), .ZN(new_n412));
  OAI21_X1  g226(.A(G101), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT10), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n397), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n414), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n193), .B1(new_n279), .B2(KEYINPUT1), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n298), .B1(new_n418), .B2(new_n276), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n416), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n403), .A2(new_n408), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT83), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n403), .A2(new_n408), .A3(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n423), .A2(KEYINPUT84), .A3(G101), .A4(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n403), .A2(new_n408), .A3(new_n424), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n403), .B2(new_n408), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n427), .A2(new_n428), .A3(new_n409), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n410), .A2(KEYINPUT84), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(KEYINPUT4), .B(new_n426), .C1(new_n429), .C2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT85), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT4), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n423), .A2(new_n434), .A3(G101), .A4(new_n425), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n435), .A2(new_n286), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n432), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n433), .B1(new_n432), .B2(new_n436), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n421), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n275), .A2(new_n289), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n440), .B(new_n421), .C1(new_n437), .C2(new_n438), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n396), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n397), .A2(new_n414), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n420), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT12), .A3(new_n309), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n440), .B1(new_n420), .B2(new_n445), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n447), .B1(new_n448), .B2(KEYINPUT12), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n443), .A2(new_n396), .A3(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n391), .B(new_n192), .C1(new_n444), .C2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n442), .A2(new_n443), .A3(new_n396), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n443), .A2(new_n449), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n395), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n455), .A3(G469), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n391), .A2(new_n192), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n390), .B1(new_n452), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT86), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n451), .A2(new_n458), .A3(new_n456), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(KEYINPUT86), .A3(new_n390), .ZN(new_n464));
  OAI21_X1  g278(.A(G210), .B1(G237), .B2(G902), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  OR3_X1    g280(.A1(new_n286), .A2(KEYINPUT88), .A3(new_n211), .ZN(new_n467));
  OAI21_X1  g281(.A(KEYINPUT88), .B1(new_n286), .B2(new_n211), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n397), .A2(new_n211), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G224), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(G953), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n470), .B(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G122), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n435), .A2(new_n351), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n423), .A2(G101), .A3(new_n425), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n434), .B1(new_n478), .B2(new_n430), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n477), .B1(new_n479), .B2(new_n426), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n197), .A2(G116), .ZN(new_n482));
  OAI21_X1  g296(.A(G113), .B1(new_n482), .B2(KEYINPUT5), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n253), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n417), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n476), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n474), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n255), .B1(new_n429), .B2(new_n434), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n488), .B(new_n486), .C1(new_n432), .C2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g306(.A(KEYINPUT6), .B(new_n476), .C1(new_n480), .C2(new_n486), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n473), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT7), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n472), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n470), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n469), .B1(new_n211), .B2(new_n286), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n495), .B2(new_n472), .ZN(new_n499));
  OR2_X1    g313(.A1(new_n483), .A2(KEYINPUT89), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n483), .A2(KEYINPUT89), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n500), .A2(new_n481), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n417), .B1(new_n253), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n414), .A2(new_n485), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n474), .B(KEYINPUT8), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n497), .A2(new_n499), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n432), .A2(new_n489), .ZN(new_n508));
  INV_X1    g322(.A(new_n486), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n474), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n192), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n466), .B1(new_n494), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(G902), .B1(new_n507), .B2(new_n510), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n486), .B1(new_n432), .B2(new_n489), .ZN(new_n515));
  INV_X1    g329(.A(new_n476), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n515), .A2(new_n491), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n517), .B1(new_n487), .B2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n514), .B(new_n465), .C1(new_n519), .C2(new_n473), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(G214), .B1(G237), .B2(G902), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT99), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n228), .A2(new_n225), .ZN(new_n525));
  INV_X1    g339(.A(G237), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n231), .A3(G214), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n280), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n321), .A2(G143), .A3(G214), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G131), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n268), .A3(new_n529), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n530), .A2(KEYINPUT17), .A3(G131), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n525), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(KEYINPUT18), .A2(G131), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n530), .B(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT90), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n213), .A2(G146), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n221), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n539), .B1(new_n221), .B2(new_n540), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n538), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(G113), .B(G122), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(new_n401), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n536), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT91), .B1(new_n219), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT19), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT19), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n219), .B2(KEYINPUT91), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n551), .B(new_n215), .C1(new_n550), .C2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n209), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n219), .B2(KEYINPUT16), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n531), .A2(new_n533), .B1(new_n556), .B2(G146), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n544), .A2(new_n558), .A3(KEYINPUT93), .ZN(new_n559));
  INV_X1    g373(.A(new_n546), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT93), .ZN(new_n562));
  INV_X1    g376(.A(new_n537), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n530), .B(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n221), .A2(new_n540), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT90), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n566), .B2(new_n541), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n554), .A2(new_n557), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n548), .B1(new_n561), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(G475), .A2(G902), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT20), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(new_n560), .A3(new_n559), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n547), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT20), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n571), .ZN(new_n577));
  INV_X1    g391(.A(G475), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n546), .B1(new_n536), .B2(new_n544), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n192), .B1(new_n548), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n578), .B1(new_n580), .B2(KEYINPUT94), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n536), .A2(new_n544), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n560), .ZN(new_n583));
  AOI21_X1  g397(.A(G902), .B1(new_n583), .B2(new_n547), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT94), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n573), .A2(new_n577), .B1(new_n581), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(G116), .B(G122), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n400), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n280), .A2(G128), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n193), .A2(G143), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n301), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n301), .A2(new_n592), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT14), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n588), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n597));
  INV_X1    g411(.A(G122), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(G116), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n398), .B1(new_n599), .B2(KEYINPUT14), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n596), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n597), .B1(new_n596), .B2(new_n600), .ZN(new_n602));
  OAI221_X1 g416(.A(new_n589), .B1(new_n593), .B2(new_n594), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n400), .ZN(new_n604));
  INV_X1    g418(.A(new_n588), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n593), .B1(new_n606), .B2(new_n589), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT13), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT95), .B1(new_n590), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n610), .A2(new_n280), .A3(KEYINPUT13), .A4(G128), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n590), .A2(new_n608), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n609), .A2(new_n611), .A3(new_n612), .A4(new_n591), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(G134), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT96), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n607), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n607), .B2(new_n614), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n603), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(G217), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n389), .A2(new_n619), .A3(G953), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n603), .B(new_n620), .C1(new_n616), .C2(new_n617), .ZN(new_n623));
  AOI21_X1  g437(.A(G902), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(G478), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(KEYINPUT15), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n624), .B(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n587), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(G952), .ZN(new_n631));
  AOI211_X1 g445(.A(G953), .B(new_n631), .C1(G234), .C2(G237), .ZN(new_n632));
  OAI211_X1 g446(.A(G902), .B(G953), .C1(new_n187), .C2(new_n526), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n633), .B(KEYINPUT98), .Z(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT21), .B(G898), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n524), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n636), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n587), .A2(KEYINPUT99), .A3(new_n638), .A4(new_n629), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n523), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n388), .A2(new_n462), .A3(new_n464), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G101), .ZN(G3));
  INV_X1    g456(.A(new_n522), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n513), .B2(new_n520), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n638), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n576), .B1(new_n575), .B2(new_n571), .ZN(new_n646));
  AOI211_X1 g460(.A(KEYINPUT20), .B(new_n572), .C1(new_n574), .C2(new_n547), .ZN(new_n647));
  OAI21_X1  g461(.A(G475), .B1(new_n584), .B2(new_n585), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n580), .A2(KEYINPUT94), .ZN(new_n649));
  OAI22_X1  g463(.A1(new_n646), .A2(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n622), .A2(new_n623), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT33), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT33), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n622), .A2(new_n653), .A3(new_n623), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n652), .A2(G478), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n625), .A2(new_n192), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n624), .B2(new_n625), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n656), .B1(new_n655), .B2(new_n658), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n650), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n645), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(G902), .B1(new_n340), .B2(new_n355), .ZN(new_n663));
  INV_X1    g477(.A(G472), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n663), .B1(KEYINPUT100), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n248), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n664), .A2(KEYINPUT100), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n373), .A2(new_n374), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n668), .A2(new_n342), .B1(new_n327), .B2(new_n339), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n667), .B1(new_n669), .B2(G902), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n665), .A2(new_n666), .A3(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n462), .A2(new_n662), .A3(new_n464), .A4(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT34), .B(G104), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  NAND3_X1  g488(.A1(new_n462), .A2(new_n464), .A3(new_n671), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n580), .A2(KEYINPUT94), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n586), .A3(G475), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n677), .B(new_n628), .C1(new_n646), .C2(new_n647), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n521), .A2(new_n638), .A3(new_n679), .A4(new_n522), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT35), .B(G107), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G9));
  NAND2_X1  g497(.A1(new_n222), .A2(new_n230), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n235), .A2(KEYINPUT36), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n246), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n243), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n665), .A2(new_n670), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n462), .A2(new_n640), .A3(new_n464), .A4(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT37), .B(G110), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G12));
  NAND2_X1  g508(.A1(new_n364), .A2(new_n387), .ZN(new_n695));
  INV_X1    g509(.A(G900), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n632), .B1(new_n634), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n698), .B1(new_n243), .B2(new_n688), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n523), .A2(new_n678), .A3(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n462), .A2(new_n695), .A3(new_n700), .A4(new_n464), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G128), .ZN(G30));
  XNOR2_X1  g516(.A(new_n521), .B(KEYINPUT38), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n359), .B1(new_n669), .B2(new_n358), .ZN(new_n704));
  OAI21_X1  g518(.A(KEYINPUT73), .B1(new_n669), .B2(new_n362), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n356), .A2(new_n249), .A3(new_n360), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n319), .A2(new_n326), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n346), .A2(new_n377), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n341), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n192), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G472), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n704), .A2(new_n705), .A3(new_n706), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n650), .A2(new_n628), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n690), .A2(new_n713), .A3(new_n643), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n703), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT102), .ZN(new_n716));
  INV_X1    g530(.A(new_n390), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n443), .A2(new_n396), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n718), .A2(new_n442), .B1(new_n454), .B2(new_n395), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n457), .B1(new_n719), .B2(G469), .ZN(new_n720));
  AOI211_X1 g534(.A(new_n461), .B(new_n717), .C1(new_n720), .C2(new_n451), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT86), .B1(new_n463), .B2(new_n390), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT40), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n697), .B(KEYINPUT39), .Z(new_n725));
  NAND3_X1  g539(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n725), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT40), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n716), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT103), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT103), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n716), .A2(new_n731), .A3(new_n726), .A4(new_n728), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n280), .ZN(G45));
  NOR2_X1   g548(.A1(new_n661), .A2(new_n699), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n735), .A2(new_n644), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n462), .A2(new_n695), .A3(new_n464), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G146), .ZN(G48));
  OAI21_X1  g552(.A(new_n192), .B1(new_n444), .B2(new_n450), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(G469), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n390), .A3(new_n451), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT104), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n740), .A2(new_n743), .A3(new_n390), .A4(new_n451), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n388), .A2(new_n662), .A3(new_n742), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT41), .B(G113), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT105), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n745), .B(new_n747), .ZN(G15));
  INV_X1    g562(.A(new_n680), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n388), .A2(new_n749), .A3(new_n742), .A4(new_n744), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G116), .ZN(G18));
  NOR2_X1   g565(.A1(new_n741), .A2(new_n523), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n689), .B1(new_n637), .B2(new_n639), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n753), .A3(new_n695), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G119), .ZN(G21));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n756), .B1(new_n663), .B2(new_n664), .ZN(new_n757));
  OAI211_X1 g571(.A(KEYINPUT106), .B(G472), .C1(new_n669), .C2(G902), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n341), .B1(new_n378), .B2(new_n349), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n357), .B1(new_n371), .B2(new_n759), .ZN(new_n760));
  AND4_X1   g574(.A1(new_n666), .A2(new_n757), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n645), .A2(new_n713), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n742), .A3(new_n744), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G122), .ZN(G24));
  AND4_X1   g578(.A1(new_n690), .A2(new_n757), .A3(new_n758), .A4(new_n760), .ZN(new_n765));
  INV_X1    g579(.A(new_n660), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n650), .A3(new_n698), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n765), .A2(new_n752), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G125), .ZN(G27));
  AOI21_X1  g586(.A(new_n717), .B1(new_n720), .B2(new_n451), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n513), .A2(new_n520), .A3(new_n522), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT107), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n513), .A2(new_n520), .A3(KEYINPUT107), .A4(new_n522), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n769), .A2(KEYINPUT42), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n388), .A2(new_n773), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n386), .A2(G472), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n356), .A2(new_n360), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n704), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n770), .A3(new_n666), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n776), .A2(new_n463), .A3(new_n390), .A4(new_n777), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT42), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n780), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n268), .ZN(G33));
  NOR2_X1   g602(.A1(new_n678), .A2(new_n697), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n388), .A2(new_n773), .A3(new_n778), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  OAI21_X1  g605(.A(new_n587), .B1(new_n659), .B2(new_n660), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n792), .A2(new_n793), .A3(KEYINPUT43), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT43), .B1(new_n792), .B2(new_n793), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n689), .B1(new_n665), .B2(new_n670), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(KEYINPUT44), .A3(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n798), .A2(KEYINPUT110), .A3(new_n778), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT110), .B1(new_n798), .B2(new_n778), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n796), .A2(new_n797), .ZN(new_n801));
  OAI22_X1  g615(.A1(new_n799), .A2(new_n800), .B1(KEYINPUT44), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n453), .A2(new_n455), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n391), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n719), .A2(KEYINPUT45), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n457), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT46), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n451), .B1(new_n807), .B2(KEYINPUT46), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n390), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n725), .ZN(new_n812));
  OR3_X1    g626(.A1(new_n811), .A2(KEYINPUT108), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT108), .B1(new_n811), .B2(new_n812), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n802), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(new_n263), .ZN(G39));
  NAND2_X1  g630(.A1(new_n776), .A2(new_n777), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n695), .A2(new_n817), .A3(new_n666), .A4(new_n769), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT47), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n811), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n805), .A2(new_n806), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n458), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT46), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n451), .A3(new_n808), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT47), .B1(new_n825), .B2(new_n390), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n818), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  NAND4_X1  g642(.A1(new_n745), .A2(new_n750), .A3(new_n763), .A4(new_n754), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT113), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n757), .A2(new_n735), .A3(new_n758), .A4(new_n760), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n785), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n705), .A2(new_n706), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n358), .B1(new_n340), .B2(new_n355), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n320), .B1(new_n338), .B2(new_n255), .ZN(new_n835));
  INV_X1    g649(.A(new_n325), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT29), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n373), .A2(new_n374), .A3(new_n341), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n380), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI22_X1  g653(.A1(KEYINPUT32), .A2(new_n834), .B1(new_n839), .B2(new_n664), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n666), .B1(new_n833), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n785), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n832), .B1(new_n842), .B2(new_n789), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n630), .A2(new_n699), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n776), .A2(new_n777), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n462), .A3(new_n695), .A4(new_n464), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n843), .A2(new_n786), .A3(new_n780), .A4(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n680), .B(KEYINPUT111), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n723), .A3(new_n671), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n641), .A3(new_n672), .A4(new_n692), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n847), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n523), .A2(new_n713), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n690), .A2(new_n697), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n712), .A3(new_n773), .A4(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n701), .A2(new_n737), .A3(new_n771), .A4(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n856), .B(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n830), .A2(new_n852), .A3(new_n858), .ZN(new_n859));
  XOR2_X1   g673(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n860));
  XNOR2_X1  g674(.A(new_n856), .B(KEYINPUT52), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n785), .A2(new_n831), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n790), .A2(new_n846), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n787), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT111), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n680), .B(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n692), .B1(new_n675), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n641), .A2(new_n672), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n745), .A2(new_n750), .A3(new_n763), .A4(new_n754), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n864), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n860), .B1(new_n861), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n859), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n851), .B1(new_n861), .B2(new_n871), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n847), .A2(new_n850), .A3(new_n829), .ZN(new_n876));
  INV_X1    g690(.A(new_n860), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n858), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n873), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n761), .A2(new_n796), .A3(new_n632), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n820), .A2(new_n826), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n740), .A2(new_n451), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n390), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n778), .B(new_n881), .C1(new_n882), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n796), .A2(new_n632), .ZN(new_n886));
  INV_X1    g700(.A(new_n741), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n778), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n765), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n703), .A2(new_n522), .A3(new_n741), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n881), .A2(KEYINPUT50), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT50), .B1(new_n881), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n712), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n666), .A3(new_n632), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n897));
  OR3_X1    g711(.A1(new_n896), .A2(new_n888), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n897), .B1(new_n896), .B2(new_n888), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n768), .A2(new_n650), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n894), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n885), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT51), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n898), .A2(new_n650), .A3(new_n768), .A4(new_n899), .ZN(new_n905));
  AOI211_X1 g719(.A(new_n631), .B(G953), .C1(new_n881), .C2(new_n752), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT115), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n248), .B1(new_n387), .B2(new_n782), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n889), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT48), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT115), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n905), .A2(new_n912), .A3(new_n906), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n908), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n880), .B(new_n904), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n631), .A2(new_n231), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT117), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n703), .B1(KEYINPUT49), .B2(new_n883), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n666), .A2(new_n390), .A3(new_n522), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n712), .A2(new_n792), .A3(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n922), .B(new_n924), .C1(KEYINPUT49), .C2(new_n883), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n921), .A2(new_n925), .ZN(G75));
  NOR2_X1   g740(.A1(new_n231), .A2(G952), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n859), .A2(new_n872), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n929), .A2(KEYINPUT120), .A3(G210), .A4(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n519), .B(new_n473), .Z(new_n931));
  XNOR2_X1  g745(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n931), .B(new_n932), .Z(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(KEYINPUT56), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n192), .B1(new_n859), .B2(new_n872), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT120), .B1(new_n936), .B2(G210), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n928), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT56), .B1(new_n936), .B2(G210), .ZN(new_n940));
  INV_X1    g754(.A(new_n933), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n936), .A2(G210), .ZN(new_n943));
  OAI211_X1 g757(.A(KEYINPUT119), .B(new_n933), .C1(new_n943), .C2(KEYINPUT56), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n938), .B1(new_n942), .B2(new_n944), .ZN(G51));
  AOI21_X1  g759(.A(new_n873), .B1(new_n859), .B2(new_n872), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n874), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n457), .B(KEYINPUT57), .Z(new_n948));
  OAI22_X1  g762(.A1(new_n947), .A2(new_n948), .B1(new_n444), .B2(new_n450), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n936), .A2(new_n806), .A3(new_n805), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n927), .B1(new_n949), .B2(new_n950), .ZN(G54));
  NAND2_X1  g765(.A1(KEYINPUT58), .A2(G475), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT121), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n936), .A2(new_n575), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n575), .B1(new_n936), .B2(new_n953), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n954), .A2(new_n955), .A3(new_n927), .ZN(G60));
  INV_X1    g770(.A(KEYINPUT123), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n657), .B(KEYINPUT59), .ZN(new_n958));
  INV_X1    g772(.A(new_n878), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT53), .B1(new_n876), .B2(new_n858), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT54), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n859), .A2(new_n872), .A3(new_n873), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n652), .A2(new_n654), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n957), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n964), .ZN(new_n966));
  OAI211_X1 g780(.A(KEYINPUT123), .B(new_n966), .C1(new_n880), .C2(new_n958), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT122), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n966), .A2(new_n958), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n745), .A2(new_n754), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n971), .A2(KEYINPUT113), .A3(new_n750), .A4(new_n763), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n867), .A2(new_n868), .A3(new_n851), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT113), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n829), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n972), .A2(new_n973), .A3(new_n864), .A4(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n976), .A2(new_n861), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n877), .B1(new_n876), .B2(new_n858), .ZN(new_n978));
  OAI21_X1  g792(.A(KEYINPUT54), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n970), .B1(new_n979), .B2(new_n962), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n968), .B1(new_n980), .B2(new_n927), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n969), .B1(new_n874), .B2(new_n946), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n982), .A2(KEYINPUT122), .A3(new_n928), .ZN(new_n983));
  AOI22_X1  g797(.A1(new_n965), .A2(new_n967), .B1(new_n981), .B2(new_n983), .ZN(G63));
  NAND2_X1  g798(.A1(G217), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT60), .Z(new_n986));
  NAND2_X1  g800(.A1(new_n929), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n238), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n987), .A2(new_n236), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n929), .A2(new_n686), .A3(new_n986), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n989), .A2(new_n928), .A3(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT61), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n989), .A2(KEYINPUT61), .A3(new_n928), .A4(new_n990), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(G66));
  NAND2_X1  g809(.A1(new_n869), .A2(new_n870), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n231), .ZN(new_n997));
  OAI21_X1  g811(.A(G953), .B1(new_n635), .B2(new_n471), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n519), .B1(G898), .B2(new_n231), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(G69));
  OAI21_X1  g815(.A(G953), .B1(new_n393), .B2(new_n696), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n909), .A2(new_n853), .ZN(new_n1003));
  AOI22_X1  g817(.A1(new_n802), .A2(new_n1003), .B1(new_n813), .B2(new_n814), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n701), .A2(new_n737), .A3(new_n771), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT124), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n787), .B1(new_n842), .B2(new_n789), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n827), .A2(new_n1007), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n231), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n696), .A2(G953), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n1011), .A2(KEYINPUT125), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(KEYINPUT125), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n551), .B1(new_n550), .B2(new_n553), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n367), .B(new_n1015), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1016), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1018), .A2(G953), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1005), .B(KEYINPUT124), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n730), .A2(new_n1021), .A3(new_n732), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT62), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n661), .A2(new_n678), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n388), .A2(new_n778), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n827), .B1(new_n727), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n815), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1020), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1002), .B1(new_n1017), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1013), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1034), .A2(new_n1019), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1002), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1030), .A2(new_n1037), .ZN(G72));
  NAND2_X1  g852(.A1(new_n384), .A2(new_n836), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1039), .B(KEYINPUT126), .ZN(new_n1040));
  NOR3_X1   g854(.A1(new_n1004), .A2(new_n1010), .A3(new_n996), .ZN(new_n1041));
  NAND2_X1  g855(.A1(G472), .A2(G902), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1042), .B(KEYINPUT63), .Z(new_n1043));
  INV_X1    g857(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1040), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n959), .A2(new_n960), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n835), .A2(new_n836), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n707), .B1(new_n1047), .B2(KEYINPUT127), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1048), .B1(KEYINPUT127), .B2(new_n1047), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1049), .A2(new_n1043), .ZN(new_n1050));
  OAI211_X1 g864(.A(new_n1045), .B(new_n928), .C1(new_n1046), .C2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1043), .B1(new_n1034), .B2(new_n996), .ZN(new_n1052));
  NOR2_X1   g866(.A1(new_n384), .A2(new_n836), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(G57));
endmodule


