//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n794, new_n795, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n202), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(G8gat), .Z(new_n207));
  NOR2_X1   g006(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n210), .A2(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT15), .ZN(new_n213));
  XOR2_X1   g012(.A(G43gat), .B(G50gat), .Z(new_n214));
  OR3_X1    g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(new_n213), .ZN(new_n216));
  NAND2_X1  g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n208), .A2(KEYINPUT91), .A3(new_n209), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT91), .B1(new_n208), .B2(new_n209), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n211), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(new_n213), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n216), .A2(new_n217), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n207), .B1(new_n215), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n215), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT92), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n223), .B1(new_n227), .B2(new_n207), .ZN(new_n228));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT18), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n207), .B(new_n224), .Z(new_n231));
  XOR2_X1   g030(.A(new_n229), .B(KEYINPUT13), .Z(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT93), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n233), .A2(KEYINPUT93), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n230), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT89), .B(G197gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(KEYINPUT11), .B(G169gat), .Z(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT90), .B(KEYINPUT12), .Z(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n228), .A2(KEYINPUT18), .A3(new_n229), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n236), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n244), .B1(new_n236), .B2(new_n245), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G64gat), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n250), .A2(G57gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(G57gat), .ZN(new_n252));
  AND2_X1   g051(.A1(G71gat), .A2(G78gat), .ZN(new_n253));
  OAI22_X1  g052(.A1(new_n251), .A2(new_n252), .B1(KEYINPUT9), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(G71gat), .A2(G78gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n254), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT94), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT95), .B(KEYINPUT21), .Z(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G231gat), .A2(G233gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G127gat), .B(G155gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT20), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n262), .B(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(G183gat), .B(G211gat), .Z(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT21), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n207), .B1(new_n258), .B2(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(KEYINPUT96), .B(KEYINPUT19), .Z(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n267), .B(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT98), .B(KEYINPUT7), .ZN(new_n274));
  INV_X1    g073(.A(G85gat), .ZN(new_n275));
  INV_X1    g074(.A(G92gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n274), .A2(new_n277), .ZN(new_n279));
  NAND2_X1  g078(.A1(G99gat), .A2(G106gat), .ZN(new_n280));
  AOI22_X1  g079(.A1(KEYINPUT8), .A2(new_n280), .B1(new_n275), .B2(new_n276), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G99gat), .B(G106gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT99), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n224), .ZN(new_n287));
  NAND3_X1  g086(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT102), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(KEYINPUT102), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT100), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n286), .B(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT101), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(new_n227), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G190gat), .B(G218gat), .Z(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n296), .B1(new_n295), .B2(new_n227), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n298), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n304), .B(KEYINPUT97), .Z(new_n305));
  XNOR2_X1  g104(.A(G134gat), .B(G162gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n293), .A2(new_n297), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n299), .B1(new_n308), .B2(new_n301), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n303), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n307), .B1(new_n303), .B2(new_n309), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G230gat), .A2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n284), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n258), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT103), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n282), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n257), .B1(new_n317), .B2(new_n283), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(new_n283), .B2(new_n317), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n313), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n320), .B(KEYINPUT105), .Z(new_n321));
  XNOR2_X1  g120(.A(G120gat), .B(G148gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(G176gat), .B(G204gat), .ZN(new_n323));
  XOR2_X1   g122(.A(new_n322), .B(new_n323), .Z(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT10), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n258), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n286), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n315), .A2(new_n327), .A3(new_n319), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT104), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n331), .A2(new_n332), .B1(G230gat), .B2(G233gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n329), .A2(KEYINPUT104), .A3(new_n330), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n326), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n313), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n325), .B1(new_n321), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n273), .A2(new_n312), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n343));
  OR2_X1    g142(.A1(G197gat), .A2(G204gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(G197gat), .A2(G204gat), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(G211gat), .B(G218gat), .Z(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n349), .B1(new_n346), .B2(new_n347), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n354));
  INV_X1    g153(.A(G148gat), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(G141gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(G141gat), .ZN(new_n357));
  INV_X1    g156(.A(G141gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n356), .A2(new_n359), .A3(KEYINPUT78), .A4(new_n357), .ZN(new_n363));
  NAND2_X1  g162(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT2), .ZN(new_n365));
  INV_X1    g164(.A(G162gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G155gat), .ZN(new_n367));
  INV_X1    g166(.A(G155gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G162gat), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n365), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n362), .A2(new_n363), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n373));
  INV_X1    g172(.A(new_n357), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n355), .A2(G141gat), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n367), .A2(new_n369), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n371), .A2(new_n372), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n353), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n370), .A2(new_n363), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n382), .A2(new_n362), .B1(new_n376), .B2(new_n377), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n351), .A2(new_n384), .A3(new_n352), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n385), .B2(new_n372), .ZN(new_n386));
  OAI211_X1 g185(.A(G228gat), .B(G233gat), .C1(new_n381), .C2(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n346), .A2(new_n349), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n380), .B1(new_n346), .B2(new_n349), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n372), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n371), .A2(new_n378), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n390), .A2(new_n391), .B1(G228gat), .B2(G233gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n381), .B2(KEYINPUT83), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n394));
  AOI211_X1 g193(.A(new_n394), .B(new_n353), .C1(new_n379), .C2(new_n380), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n387), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT31), .B(G50gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G78gat), .B(G106gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(G22gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n397), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n387), .B(new_n401), .C1(new_n393), .C2(new_n395), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n398), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n400), .B1(new_n398), .B2(new_n402), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT0), .ZN(new_n407));
  XNOR2_X1  g206(.A(G57gat), .B(G85gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g208(.A(KEYINPUT39), .ZN(new_n410));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G120gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(G113gat), .ZN(new_n414));
  INV_X1    g213(.A(G113gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G120gat), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT1), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G127gat), .B(G134gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G134gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G127gat), .ZN(new_n421));
  INV_X1    g220(.A(G127gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G134gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n423), .A3(KEYINPUT65), .ZN(new_n424));
  OR3_X1    g223(.A1(new_n422), .A2(KEYINPUT65), .A3(G134gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n426), .A2(KEYINPUT66), .A3(new_n417), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT66), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n422), .A2(KEYINPUT65), .A3(G134gat), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n418), .B2(KEYINPUT65), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n416), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT1), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n428), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n419), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n435), .A2(KEYINPUT4), .A3(new_n391), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT66), .B1(new_n426), .B2(new_n417), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n430), .A2(new_n428), .A3(new_n433), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n438), .A2(new_n439), .B1(new_n417), .B2(new_n418), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n437), .B1(new_n440), .B2(new_n383), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n436), .A2(new_n441), .A3(KEYINPUT81), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(KEYINPUT81), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n391), .A2(KEYINPUT3), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(new_n435), .A3(new_n379), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n410), .B(new_n412), .C1(new_n442), .C2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n442), .ZN(new_n448));
  INV_X1    g247(.A(new_n446), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n411), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n391), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n440), .A2(new_n383), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT39), .B1(new_n453), .B2(new_n412), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n409), .B(new_n447), .C1(new_n450), .C2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(KEYINPUT40), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n412), .A2(KEYINPUT5), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n448), .A2(new_n449), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT5), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n453), .B2(new_n412), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n411), .B(new_n445), .C1(new_n436), .C2(new_n441), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT80), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT80), .B1(new_n462), .B2(new_n463), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n409), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n455), .A2(new_n457), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT75), .ZN(new_n469));
  INV_X1    g268(.A(new_n380), .ZN(new_n470));
  NAND2_X1  g269(.A1(G169gat), .A2(G176gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(G183gat), .A2(G190gat), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n471), .B1(new_n472), .B2(KEYINPUT24), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT23), .ZN(new_n475));
  INV_X1    g274(.A(G169gat), .ZN(new_n476));
  INV_X1    g275(.A(G176gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G183gat), .ZN(new_n481));
  INV_X1    g280(.A(G190gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(KEYINPUT24), .A3(new_n472), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n474), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT25), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n474), .A2(new_n480), .A3(new_n484), .A4(KEYINPUT25), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT26), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT26), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n471), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(G169gat), .A2(G176gat), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n472), .B(new_n490), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT64), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n493), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n476), .A2(new_n477), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n500), .A3(KEYINPUT64), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n481), .A2(KEYINPUT27), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT27), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G183gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n504), .A3(new_n482), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT28), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT27), .B(G183gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT28), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n508), .A3(new_n482), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n496), .A2(new_n501), .A3(new_n506), .A4(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n470), .B1(new_n489), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G226gat), .A2(G233gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT72), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(KEYINPUT73), .Z(new_n514));
  OAI21_X1  g313(.A(new_n469), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n514), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n501), .A2(new_n506), .A3(new_n509), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n517), .A2(new_n496), .B1(new_n487), .B2(new_n488), .ZN(new_n518));
  OAI211_X1 g317(.A(KEYINPUT75), .B(new_n516), .C1(new_n518), .C2(new_n470), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n473), .B1(new_n479), .B2(new_n478), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT25), .B1(new_n520), .B2(new_n484), .ZN(new_n521));
  INV_X1    g320(.A(new_n488), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n501), .A2(new_n506), .A3(new_n509), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT64), .B1(new_n497), .B2(new_n500), .ZN(new_n524));
  OAI22_X1  g323(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n513), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n515), .A2(new_n519), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n353), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(KEYINPUT76), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n518), .A2(KEYINPUT29), .ZN(new_n530));
  OAI221_X1 g329(.A(new_n353), .B1(new_n516), .B2(new_n518), .C1(new_n530), .C2(new_n513), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n527), .A2(new_n528), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT76), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G8gat), .B(G36gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(G64gat), .B(G92gat), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n538), .B(new_n539), .Z(new_n540));
  NAND4_X1  g339(.A1(new_n533), .A2(new_n534), .A3(new_n537), .A4(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n540), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT76), .B1(new_n527), .B2(new_n528), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n542), .B1(new_n532), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n537), .A2(new_n531), .A3(new_n529), .A4(new_n540), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(KEYINPUT30), .A3(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n458), .A2(new_n468), .A3(new_n541), .A4(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n527), .A2(new_n528), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT85), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI22_X1  g350(.A1(new_n530), .A2(new_n513), .B1(new_n516), .B2(new_n518), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n550), .B1(new_n552), .B2(new_n528), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(new_n528), .B2(new_n527), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT38), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n533), .A2(new_n537), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n555), .B(new_n542), .C1(new_n556), .C2(KEYINPUT37), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n462), .A2(new_n463), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT80), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT80), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n563));
  NAND4_X1  g362(.A1(new_n562), .A2(new_n460), .A3(new_n563), .A4(new_n467), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n467), .A2(new_n563), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n467), .A2(new_n563), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n466), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n557), .A2(new_n564), .A3(new_n567), .A4(new_n545), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT38), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n544), .B1(new_n548), .B2(new_n540), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n556), .A2(KEYINPUT37), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n405), .B(new_n547), .C1(new_n568), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n518), .A2(new_n435), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n525), .A2(new_n440), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(G227gat), .ZN(new_n577));
  INV_X1    g376(.A(G233gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT68), .ZN(new_n585));
  XNOR2_X1  g384(.A(G15gat), .B(G43gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(G71gat), .B(G99gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n574), .A2(new_n579), .A3(new_n575), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n588), .B1(new_n589), .B2(KEYINPUT32), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n589), .A2(KEYINPUT67), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT67), .B1(new_n589), .B2(new_n591), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n585), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n596), .A2(KEYINPUT68), .A3(new_n592), .A4(new_n590), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n589), .B(KEYINPUT32), .C1(new_n591), .C2(new_n588), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n584), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n599), .ZN(new_n601));
  AOI211_X1 g400(.A(new_n601), .B(new_n583), .C1(new_n595), .C2(new_n597), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n604));
  OR3_X1    g403(.A1(new_n603), .A2(KEYINPUT70), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n546), .A2(new_n541), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n567), .A2(new_n564), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n405), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n604), .B1(new_n603), .B2(KEYINPUT70), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n573), .A2(new_n605), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n598), .A2(new_n599), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n583), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n599), .A3(new_n584), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(new_n405), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT35), .B1(new_n616), .B2(new_n608), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT35), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n606), .A2(new_n618), .A3(new_n607), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n614), .A2(KEYINPUT86), .A3(new_n615), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT86), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(new_n600), .B2(new_n602), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n619), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT87), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n617), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n606), .A2(new_n607), .A3(new_n618), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT86), .B1(new_n614), .B2(new_n615), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n600), .A2(new_n602), .A3(new_n621), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(KEYINPUT87), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n612), .B1(new_n625), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT88), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT88), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n612), .B(new_n633), .C1(new_n625), .C2(new_n630), .ZN(new_n634));
  AOI211_X1 g433(.A(new_n249), .B(new_n342), .C1(new_n632), .C2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n607), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G1gat), .ZN(G1324gat));
  INV_X1    g437(.A(KEYINPUT42), .ZN(new_n639));
  INV_X1    g438(.A(new_n606), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT106), .Z(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT16), .B(G8gat), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(G8gat), .ZN(new_n645));
  OR3_X1    g444(.A1(new_n641), .A2(new_n639), .A3(new_n643), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(G1325gat));
  NAND2_X1  g446(.A1(new_n620), .A2(new_n622), .ZN(new_n648));
  AOI21_X1  g447(.A(G15gat), .B1(new_n635), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n605), .A2(new_n611), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(G15gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT107), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n649), .B1(new_n635), .B2(new_n652), .ZN(G1326gat));
  NAND2_X1  g452(.A1(new_n635), .A2(new_n609), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT43), .B(G22gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1327gat));
  NAND2_X1  g455(.A1(new_n632), .A2(new_n634), .ZN(new_n657));
  NOR4_X1   g456(.A1(new_n273), .A2(new_n312), .A3(new_n249), .A4(new_n340), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(G29gat), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(new_n660), .A3(new_n636), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT45), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n312), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n634), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n629), .A2(KEYINPUT87), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n623), .A2(new_n624), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n667), .A3(new_n617), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n633), .B1(new_n668), .B2(new_n612), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n664), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n310), .A2(new_n311), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n631), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n663), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n273), .A2(new_n249), .A3(new_n340), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT108), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n670), .A2(new_n677), .A3(new_n673), .A4(new_n674), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n676), .A2(new_n636), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n662), .B1(new_n679), .B2(new_n660), .ZN(G1328gat));
  NAND3_X1  g479(.A1(new_n676), .A2(new_n640), .A3(new_n678), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n209), .B1(new_n681), .B2(KEYINPUT109), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(KEYINPUT109), .B2(new_n681), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n659), .A2(new_n209), .A3(new_n640), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT46), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(G1329gat));
  INV_X1    g485(.A(new_n650), .ZN(new_n687));
  OAI21_X1  g486(.A(G43gat), .B1(new_n675), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT47), .ZN(new_n689));
  INV_X1    g488(.A(new_n648), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(G43gat), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n658), .B(new_n691), .C1(new_n665), .C2(new_n669), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n657), .A2(KEYINPUT110), .A3(new_n658), .A4(new_n691), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n689), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n688), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n676), .A2(new_n650), .A3(new_n678), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G43gat), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT111), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n694), .A2(new_n700), .A3(new_n695), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n694), .B2(new_n695), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT112), .B1(new_n704), .B2(new_n689), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT112), .ZN(new_n706));
  AOI211_X1 g505(.A(new_n706), .B(KEYINPUT47), .C1(new_n699), .C2(new_n703), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n697), .B1(new_n705), .B2(new_n707), .ZN(G1330gat));
  OAI21_X1  g507(.A(G50gat), .B1(new_n675), .B2(new_n405), .ZN(new_n709));
  INV_X1    g508(.A(G50gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n659), .A2(new_n710), .A3(new_n609), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(KEYINPUT48), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n711), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n676), .A2(new_n609), .A3(new_n678), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(G50gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n712), .B1(new_n715), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g515(.A1(new_n671), .A2(new_n272), .ZN(new_n717));
  AND4_X1   g516(.A1(new_n631), .A2(new_n249), .A3(new_n717), .A4(new_n340), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n636), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT113), .B(G57gat), .Z(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1332gat));
  AOI21_X1  g520(.A(new_n606), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT114), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1333gat));
  NAND2_X1  g525(.A1(new_n718), .A2(new_n650), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n690), .A2(G71gat), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n727), .A2(G71gat), .B1(new_n718), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1334gat));
  NAND2_X1  g530(.A1(new_n718), .A2(new_n609), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G78gat), .ZN(G1335gat));
  INV_X1    g532(.A(new_n249), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n273), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n631), .A2(new_n671), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n736), .A2(KEYINPUT51), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(KEYINPUT51), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n737), .A2(new_n738), .A3(new_n341), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n739), .A2(new_n275), .A3(new_n636), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n670), .A2(new_n340), .A3(new_n673), .A4(new_n735), .ZN(new_n741));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741), .B2(new_n607), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(G1336gat));
  OAI21_X1  g542(.A(G92gat), .B1(new_n741), .B2(new_n606), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n739), .A2(new_n276), .A3(new_n640), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g546(.A(G99gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n739), .A2(new_n748), .A3(new_n648), .ZN(new_n749));
  OAI21_X1  g548(.A(G99gat), .B1(new_n741), .B2(new_n687), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(G1338gat));
  OAI21_X1  g550(.A(G106gat), .B1(new_n741), .B2(new_n405), .ZN(new_n752));
  INV_X1    g551(.A(G106gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n739), .A2(new_n753), .A3(new_n609), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g555(.A1(new_n717), .A2(new_n249), .A3(new_n341), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n325), .B1(new_n337), .B2(KEYINPUT54), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n335), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT54), .B1(new_n331), .B2(new_n313), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n759), .B(KEYINPUT55), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n761), .B1(new_n333), .B2(new_n334), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(new_n758), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n762), .A2(new_n765), .A3(new_n336), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n310), .B2(new_n311), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n228), .A2(new_n229), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n231), .A2(new_n232), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n241), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n246), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n340), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n766), .B2(new_n249), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n769), .A2(new_n773), .B1(new_n775), .B2(new_n312), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n757), .B1(new_n776), .B2(new_n273), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n636), .ZN(new_n778));
  OR3_X1    g577(.A1(new_n778), .A2(new_n640), .A3(new_n616), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(G113gat), .B1(new_n780), .B2(new_n734), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n769), .A2(new_n773), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n775), .A2(new_n312), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n273), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n757), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n786), .A2(new_n609), .A3(new_n690), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n787), .A2(new_n636), .A3(new_n606), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n788), .A2(new_n415), .A3(new_n249), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n781), .A2(new_n789), .ZN(G1340gat));
  AOI21_X1  g589(.A(G120gat), .B1(new_n780), .B2(new_n340), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n788), .A2(new_n413), .A3(new_n341), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(G1341gat));
  OAI21_X1  g592(.A(G127gat), .B1(new_n788), .B2(new_n272), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n273), .A2(new_n422), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n779), .B2(new_n795), .ZN(G1342gat));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n420), .A3(new_n671), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n797), .A2(KEYINPUT56), .ZN(new_n798));
  OAI21_X1  g597(.A(G134gat), .B1(new_n788), .B2(new_n312), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(KEYINPUT56), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(G1343gat));
  NOR3_X1   g600(.A1(new_n650), .A2(new_n607), .A3(new_n640), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT57), .B1(new_n777), .B2(new_n609), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n609), .A2(KEYINPUT57), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n769), .A2(new_n773), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n766), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n762), .A2(new_n765), .A3(KEYINPUT116), .A4(new_n336), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n734), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n671), .B1(new_n809), .B2(new_n774), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n272), .B1(new_n805), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n804), .B1(new_n811), .B2(new_n757), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n734), .B(new_n802), .C1(new_n803), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G141gat), .ZN(new_n814));
  XOR2_X1   g613(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n815));
  NAND4_X1  g614(.A1(new_n777), .A2(new_n636), .A3(new_n609), .A4(new_n687), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n816), .A2(KEYINPUT118), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(KEYINPUT118), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n606), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n734), .A2(new_n358), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n814), .B(new_n815), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n814), .A2(KEYINPUT117), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n813), .B2(G141gat), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n816), .A2(new_n640), .A3(new_n820), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n821), .B1(new_n826), .B2(new_n827), .ZN(G1344gat));
  NOR2_X1   g627(.A1(new_n355), .A2(KEYINPUT59), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n802), .B1(new_n803), .B2(new_n812), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n341), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(KEYINPUT120), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(KEYINPUT120), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n671), .A2(new_n835), .A3(new_n767), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n768), .A2(KEYINPUT121), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(new_n837), .A3(new_n773), .ZN(new_n838));
  INV_X1    g637(.A(new_n810), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n273), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n609), .B1(new_n840), .B2(new_n785), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n777), .A2(KEYINPUT57), .A3(new_n609), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n802), .A2(new_n340), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n355), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI22_X1  g646(.A1(new_n832), .A2(new_n833), .B1(new_n834), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n819), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n355), .A3(new_n340), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(G1345gat));
  OAI21_X1  g650(.A(G155gat), .B1(new_n830), .B2(new_n272), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n273), .A2(new_n368), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n819), .B2(new_n853), .ZN(G1346gat));
  XOR2_X1   g653(.A(KEYINPUT79), .B(G162gat), .Z(new_n855));
  NAND3_X1  g654(.A1(new_n849), .A2(new_n671), .A3(new_n855), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n830), .A2(new_n312), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(KEYINPUT122), .ZN(new_n858));
  INV_X1    g657(.A(new_n855), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n857), .B2(KEYINPUT122), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n856), .B1(new_n858), .B2(new_n860), .ZN(G1347gat));
  NOR2_X1   g660(.A1(new_n636), .A2(new_n606), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n787), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n863), .A2(new_n476), .A3(new_n249), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n786), .A2(new_n636), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n865), .A2(new_n405), .A3(new_n640), .A4(new_n603), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n734), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n864), .B1(new_n868), .B2(new_n476), .ZN(G1348gat));
  OAI21_X1  g668(.A(G176gat), .B1(new_n863), .B2(new_n341), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n340), .A2(new_n477), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n866), .B2(new_n871), .ZN(G1349gat));
  OAI21_X1  g671(.A(G183gat), .B1(new_n863), .B2(new_n272), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n273), .A2(new_n507), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n866), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g675(.A(G190gat), .B1(new_n863), .B2(new_n312), .ZN(new_n877));
  XOR2_X1   g676(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n878));
  XNOR2_X1  g677(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n867), .A2(new_n482), .A3(new_n671), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1351gat));
  NOR3_X1   g680(.A1(new_n650), .A2(new_n405), .A3(new_n606), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n865), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(G197gat), .B1(new_n883), .B2(new_n734), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n845), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n786), .A2(new_n804), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n887), .B1(new_n841), .B2(new_n842), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT124), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n650), .A2(new_n636), .A3(new_n606), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n886), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n734), .A2(G197gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n884), .B1(new_n892), .B2(new_n893), .ZN(G1352gat));
  OAI21_X1  g693(.A(G204gat), .B1(new_n891), .B2(new_n341), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n341), .A2(G204gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n865), .A2(new_n882), .A3(new_n896), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n897), .A2(KEYINPUT125), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(KEYINPUT125), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(KEYINPUT62), .ZN(new_n902));
  XOR2_X1   g701(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n903));
  NAND3_X1  g702(.A1(new_n898), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n895), .A2(new_n902), .A3(new_n904), .ZN(G1353gat));
  INV_X1    g704(.A(G211gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n883), .A2(new_n906), .A3(new_n273), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n273), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT127), .B1(new_n888), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n910));
  INV_X1    g709(.A(new_n908), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n845), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AND4_X1   g711(.A1(KEYINPUT63), .A2(new_n909), .A3(new_n912), .A4(G211gat), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n908), .B1(new_n843), .B2(new_n844), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n906), .B1(new_n914), .B2(new_n910), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT63), .B1(new_n915), .B2(new_n909), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n907), .B1(new_n913), .B2(new_n916), .ZN(G1354gat));
  AOI21_X1  g716(.A(G218gat), .B1(new_n883), .B2(new_n671), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n671), .A2(G218gat), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n892), .B2(new_n919), .ZN(G1355gat));
endmodule


