//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n562, new_n564, new_n565, new_n566, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT64), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n465), .A2(KEYINPUT65), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT66), .Z(new_n482));
  NOR2_X1   g057(.A1(new_n479), .A2(new_n472), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n490), .A2(new_n462), .A3(new_n464), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT68), .B(KEYINPUT4), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT69), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT68), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n499), .A2(new_n476), .A3(new_n500), .A4(new_n490), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n493), .A2(new_n494), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n476), .A2(G126), .A3(G2105), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n472), .A2(G114), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  OR3_X1    g080(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT67), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT67), .B1(new_n504), .B2(new_n505), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n502), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n511), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT6), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G651), .ZN(new_n523));
  AND3_X1   g098(.A1(new_n521), .A2(new_n523), .A3(G543), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n519), .A2(G651), .B1(G50), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n521), .A2(new_n523), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(new_n516), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT71), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n527), .A2(new_n530), .A3(new_n516), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n525), .B1(new_n526), .B2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  INV_X1    g109(.A(new_n532), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G89), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n524), .A2(G51), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  AOI22_X1  g118(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n520), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT73), .ZN(new_n546));
  XOR2_X1   g121(.A(KEYINPUT74), .B(G52), .Z(new_n547));
  NAND2_X1  g122(.A1(new_n524), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n535), .A2(G90), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  NAND2_X1  g126(.A1(new_n524), .A2(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n532), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n520), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT75), .Z(new_n559));
  AND2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  XOR2_X1   g138(.A(KEYINPUT77), .B(KEYINPUT8), .Z(new_n564));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(new_n535), .A2(G91), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(new_n520), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n524), .A2(G53), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT9), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(G299));
  NAND2_X1  g148(.A1(new_n535), .A2(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n524), .A2(G49), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(new_n535), .A2(G86), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT78), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n517), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(G651), .B1(G48), .B2(new_n524), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n579), .A2(new_n584), .ZN(G305));
  XOR2_X1   g160(.A(KEYINPUT79), .B(G85), .Z(new_n586));
  NAND2_X1  g161(.A1(new_n535), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(G72), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n517), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G47), .B2(new_n524), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  XNOR2_X1  g169(.A(KEYINPUT80), .B(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n517), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(G54), .B2(new_n524), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(KEYINPUT10), .B1(new_n532), .B2(new_n600), .ZN(new_n601));
  OR3_X1    g176(.A1(new_n532), .A2(KEYINPUT10), .A3(new_n600), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n593), .B1(new_n604), .B2(G868), .ZN(G284));
  XOR2_X1   g180(.A(G284), .B(KEYINPUT82), .Z(G321));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  OR3_X1    g182(.A1(G168), .A2(KEYINPUT83), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT83), .B1(G168), .B2(new_n607), .ZN(new_n609));
  AND3_X1   g184(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n608), .B(new_n609), .C1(G868), .C2(new_n610), .ZN(G297));
  XNOR2_X1  g186(.A(G297), .B(KEYINPUT84), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n604), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n556), .A2(new_n559), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(new_n607), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n603), .A2(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n607), .ZN(G323));
  XOR2_X1   g193(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n619));
  XNOR2_X1  g194(.A(G323), .B(new_n619), .ZN(G282));
  NAND2_X1  g195(.A1(new_n483), .A2(G123), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n480), .A2(G135), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n472), .A2(G111), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  XOR2_X1   g201(.A(KEYINPUT86), .B(KEYINPUT12), .Z(new_n627));
  NOR3_X1   g202(.A1(new_n463), .A2(new_n461), .A3(G2105), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT13), .B(G2100), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n626), .A2(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT15), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2435), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n637));
  XOR2_X1   g212(.A(G2443), .B(G2446), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G1341), .B(G1348), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n642), .B(new_n643), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G14), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n649), .A2(KEYINPUT17), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  AOI21_X1  g226(.A(KEYINPUT18), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n649), .B2(KEYINPUT18), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2096), .B(G2100), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT87), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n660), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n669), .B(new_n670), .C1(new_n668), .C2(new_n667), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT88), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1981), .B(G1986), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(G229));
  NOR2_X1   g253(.A1(G16), .A2(G23), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n577), .B2(G16), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT33), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G6), .ZN(new_n684));
  INV_X1    g259(.A(G305), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT93), .B(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT32), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n683), .A2(G22), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n683), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(G1971), .Z(new_n692));
  NAND3_X1  g267(.A1(new_n682), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(KEYINPUT94), .B1(new_n693), .B2(KEYINPUT34), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n695));
  AND2_X1   g270(.A1(KEYINPUT89), .A2(G29), .ZN(new_n696));
  NOR2_X1   g271(.A1(KEYINPUT89), .A2(G29), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n699), .A2(G25), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n701));
  INV_X1    g276(.A(new_n483), .ZN(new_n702));
  INV_X1    g277(.A(G119), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n472), .A2(G107), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n480), .A2(G131), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n483), .A2(KEYINPUT91), .A3(G119), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n704), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI211_X1 g285(.A(new_n695), .B(new_n700), .C1(new_n710), .C2(new_n698), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n695), .B2(new_n700), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT35), .B(G1991), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT92), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n712), .B(new_n714), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n694), .B(new_n715), .C1(KEYINPUT34), .C2(new_n693), .ZN(new_n716));
  NOR2_X1   g291(.A1(G16), .A2(G24), .ZN(new_n717));
  INV_X1    g292(.A(G290), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(G16), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1986), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT36), .Z(new_n722));
  AOI21_X1  g297(.A(KEYINPUT28), .B1(new_n699), .B2(G26), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n699), .A2(KEYINPUT28), .A3(G26), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n483), .A2(G128), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n480), .A2(G140), .ZN(new_n727));
  OAI21_X1  g302(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n472), .A2(G116), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n726), .B(new_n727), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT95), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(KEYINPUT95), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI211_X1 g308(.A(new_n723), .B(new_n725), .C1(new_n733), .C2(G29), .ZN(new_n734));
  INV_X1    g309(.A(G2067), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n699), .A2(G27), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G164), .B2(new_n699), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G2078), .ZN(new_n739));
  NAND2_X1  g314(.A1(G171), .A2(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G5), .B2(G16), .ZN(new_n741));
  INV_X1    g316(.A(G1961), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n739), .B1(new_n743), .B2(KEYINPUT99), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n738), .A2(G2078), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n736), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G29), .ZN(new_n747));
  AND2_X1   g322(.A1(KEYINPUT30), .A2(G28), .ZN(new_n748));
  NOR2_X1   g323(.A1(KEYINPUT30), .A2(G28), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT31), .B(G11), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n750), .B(new_n751), .C1(new_n625), .C2(new_n699), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT98), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n683), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n683), .ZN(new_n755));
  INV_X1    g330(.A(G1966), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G2072), .ZN(new_n758));
  OR2_X1    g333(.A1(G29), .A2(G33), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n480), .A2(G139), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT25), .Z(new_n762));
  AOI22_X1  g337(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n760), .B(new_n762), .C1(new_n472), .C2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n759), .B1(new_n764), .B2(new_n747), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n741), .A2(new_n742), .B1(new_n758), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n746), .A2(new_n753), .A3(new_n757), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n743), .A2(KEYINPUT99), .ZN(new_n768));
  NOR2_X1   g343(.A1(G4), .A2(G16), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n604), .B2(G16), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n768), .B1(G1348), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(G1348), .ZN(new_n772));
  NAND2_X1  g347(.A1(G160), .A2(G29), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT24), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(G34), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(G34), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n699), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n773), .A2(new_n777), .B1(KEYINPUT100), .B2(G2084), .ZN(new_n778));
  NOR2_X1   g353(.A1(KEYINPUT100), .A2(G2084), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n778), .B(new_n779), .Z(new_n780));
  OAI211_X1 g355(.A(new_n772), .B(new_n780), .C1(new_n758), .C2(new_n765), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT23), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n683), .A2(G20), .ZN(new_n783));
  AOI22_X1  g358(.A1(G299), .A2(G16), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n782), .B2(new_n783), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1956), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n767), .A2(new_n771), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n683), .A2(G19), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n560), .B2(new_n683), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G1341), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n699), .A2(G35), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G162), .B2(new_n699), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT101), .B(KEYINPUT29), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2090), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n792), .B(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n722), .A2(new_n787), .A3(new_n790), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n747), .A2(G32), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n483), .A2(G129), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n480), .A2(G141), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n800));
  NAND3_X1  g375(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT26), .Z(new_n802));
  NAND4_X1  g377(.A1(new_n798), .A2(new_n799), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT96), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n797), .B1(new_n804), .B2(new_n747), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n806));
  INV_X1    g381(.A(G1996), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n805), .B(new_n808), .Z(new_n809));
  NOR2_X1   g384(.A1(new_n796), .A2(new_n809), .ZN(G311));
  OR2_X1    g385(.A1(new_n796), .A2(new_n809), .ZN(G150));
  NAND2_X1  g386(.A1(new_n524), .A2(G55), .ZN(new_n812));
  INV_X1    g387(.A(G93), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n532), .B2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT102), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(new_n520), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G860), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT37), .Z(new_n821));
  INV_X1    g396(.A(new_n819), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(new_n615), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n560), .A2(new_n819), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT39), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n604), .A2(G559), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT38), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n821), .B1(new_n829), .B2(G860), .ZN(G145));
  XNOR2_X1  g405(.A(new_n804), .B(new_n509), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n629), .B(KEYINPUT104), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n710), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n831), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n480), .A2(G142), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n472), .A2(G118), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT103), .Z(new_n838));
  OAI21_X1  g413(.A(new_n835), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G130), .B2(new_n483), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n733), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n834), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n625), .B(G160), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n487), .B(new_n843), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n764), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G37), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n842), .A2(new_n845), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g425(.A(new_n825), .B(new_n617), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n604), .A2(G299), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n603), .A2(new_n610), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n603), .B(G299), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(KEYINPUT105), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT105), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(new_n603), .B2(new_n610), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n856), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n854), .A2(new_n856), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n855), .B1(new_n865), .B2(new_n851), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(KEYINPUT42), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n577), .B(G166), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(G305), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G290), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n866), .A2(KEYINPUT42), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n867), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n867), .B2(new_n871), .ZN(new_n873));
  OAI21_X1  g448(.A(G868), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(G868), .B2(new_n822), .ZN(G295));
  OAI21_X1  g450(.A(new_n874), .B1(G868), .B2(new_n822), .ZN(G331));
  XNOR2_X1  g451(.A(G301), .B(G286), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n822), .A2(new_n615), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n560), .A2(new_n819), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n823), .A2(new_n824), .A3(new_n877), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n854), .A2(new_n859), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT107), .ZN(new_n886));
  INV_X1    g461(.A(new_n860), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT41), .A4(new_n887), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT106), .A4(new_n877), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n884), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT41), .B1(new_n852), .B2(new_n853), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n860), .B1(new_n854), .B2(new_n859), .ZN(new_n892));
  AOI211_X1 g467(.A(new_n886), .B(new_n891), .C1(new_n892), .C2(KEYINPUT41), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n881), .A2(new_n883), .ZN(new_n894));
  OAI22_X1  g469(.A1(new_n890), .A2(new_n893), .B1(new_n857), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n870), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n857), .B1(new_n884), .B2(new_n889), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n864), .A2(new_n894), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n901), .A3(new_n870), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n897), .A2(new_n898), .A3(new_n847), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT108), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n861), .A2(new_n863), .B1(new_n881), .B2(new_n883), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n896), .B1(new_n905), .B2(new_n899), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(new_n902), .A3(new_n847), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT43), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n905), .A2(new_n899), .ZN(new_n909));
  AOI21_X1  g484(.A(G37), .B1(new_n909), .B2(new_n870), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n910), .A2(new_n911), .A3(new_n898), .A4(new_n897), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n904), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n910), .A2(KEYINPUT43), .A3(new_n897), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT43), .B1(new_n910), .B2(new_n906), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT44), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(G397));
  XNOR2_X1  g494(.A(new_n733), .B(new_n735), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n804), .ZN(new_n921));
  INV_X1    g496(.A(G1384), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n509), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g498(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n468), .A2(new_n473), .A3(G40), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  AOI22_X1  g504(.A1(new_n921), .A2(new_n929), .B1(KEYINPUT125), .B2(KEYINPUT46), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n807), .ZN(new_n931));
  NOR2_X1   g506(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n931), .B(new_n932), .Z(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT126), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT47), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n804), .B(G1996), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n920), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n710), .A2(new_n713), .ZN(new_n939));
  OAI22_X1  g514(.A1(new_n938), .A2(new_n939), .B1(G2067), .B2(new_n733), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n929), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n938), .B1(new_n713), .B2(new_n710), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n939), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n929), .ZN(new_n944));
  NOR2_X1   g519(.A1(G290), .A2(G1986), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n929), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT48), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n936), .A2(new_n941), .A3(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(G305), .B(G1981), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT49), .ZN(new_n951));
  OR3_X1    g526(.A1(new_n950), .A2(KEYINPUT111), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT111), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  INV_X1    g528(.A(G8), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n509), .A2(new_n922), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n955), .B2(new_n927), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n950), .A2(new_n951), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n952), .A2(new_n953), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n577), .A2(G1976), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n959), .A2(new_n956), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n960), .B(new_n961), .C1(G1976), .C2(new_n577), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n958), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n955), .A2(KEYINPUT45), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n965), .A2(new_n926), .A3(new_n927), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n955), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n968), .B1(new_n509), .B2(new_n922), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n927), .A3(new_n971), .ZN(new_n972));
  OAI22_X1  g547(.A1(new_n967), .A2(G1971), .B1(G2090), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(G303), .A2(G8), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n974), .B(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n973), .A2(G8), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n964), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1976), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n958), .A2(new_n979), .A3(new_n577), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(G1981), .B2(G305), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n956), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n976), .B1(new_n973), .B2(G8), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n977), .A2(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n964), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n509), .A2(new_n922), .A3(new_n924), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n927), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT45), .B1(new_n509), .B2(new_n922), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n756), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(KEYINPUT112), .B(new_n756), .C1(new_n987), .C2(new_n988), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT113), .B(G2084), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n969), .A2(new_n927), .A3(new_n971), .A4(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(G8), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(G286), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n985), .A2(KEYINPUT63), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT63), .B1(new_n985), .B2(new_n997), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n978), .B(new_n982), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(KEYINPUT117), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n1002));
  NOR2_X1   g577(.A1(G168), .A2(new_n954), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n995), .A2(new_n1005), .A3(G8), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(KEYINPUT51), .B(G8), .C1(new_n995), .C2(G286), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT116), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT51), .B1(new_n996), .B2(KEYINPUT117), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1012), .A2(KEYINPUT118), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1009), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n995), .A2(new_n1003), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT62), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n966), .B2(G2078), .ZN(new_n1019));
  XOR2_X1   g594(.A(new_n1019), .B(KEYINPUT120), .Z(new_n1020));
  NOR2_X1   g595(.A1(new_n987), .A2(new_n988), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1018), .A2(G2078), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT119), .B(G1961), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n972), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1020), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1026), .A2(G171), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT62), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1014), .A2(new_n1028), .A3(new_n1015), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1017), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n927), .B(KEYINPUT122), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1031), .A2(new_n926), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT123), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1032), .A2(new_n1033), .B1(KEYINPUT45), .B2(new_n955), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1034), .B(new_n1022), .C1(new_n1033), .C2(new_n1032), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT124), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(G301), .B(KEYINPUT54), .ZN(new_n1038));
  XOR2_X1   g613(.A(new_n1025), .B(KEYINPUT121), .Z(new_n1039));
  NAND2_X1  g614(.A1(new_n1020), .A2(new_n1039), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n923), .A2(KEYINPUT50), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1042), .A2(new_n928), .A3(new_n970), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n955), .A2(new_n927), .ZN(new_n1044));
  OAI22_X1  g619(.A1(new_n1043), .A2(G1348), .B1(G2067), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT114), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n1047));
  OAI221_X1 g622(.A(new_n1047), .B1(G2067), .B2(new_n1044), .C1(new_n1043), .C2(G1348), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n603), .B1(new_n1049), .B2(KEYINPUT60), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT60), .ZN(new_n1051));
  AOI211_X1 g626(.A(new_n1051), .B(new_n604), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1052));
  OAI22_X1  g627(.A1(new_n1050), .A2(new_n1052), .B1(KEYINPUT60), .B2(new_n1049), .ZN(new_n1053));
  INV_X1    g628(.A(G1956), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n972), .A2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT56), .B(G2072), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n965), .A2(new_n926), .A3(new_n927), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(G299), .B(KEYINPUT57), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n610), .B(KEYINPUT57), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1060), .A2(KEYINPUT61), .A3(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT115), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n967), .A2(new_n807), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT58), .B(G1341), .Z(new_n1066));
  NAND2_X1  g641(.A1(new_n1044), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n615), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1068), .A2(KEYINPUT59), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT61), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1068), .A2(KEYINPUT59), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1053), .A2(new_n1064), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1060), .B1(new_n1049), .B2(new_n603), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1062), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1041), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1026), .A2(new_n1038), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n1016), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1030), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1000), .B1(new_n1079), .B2(new_n985), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n943), .B1(G1986), .B2(G290), .ZN(new_n1081));
  INV_X1    g656(.A(new_n945), .ZN(new_n1082));
  AOI211_X1 g657(.A(new_n926), .B(new_n928), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n949), .B1(new_n1080), .B2(new_n1083), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g659(.A(G229), .ZN(new_n1086));
  AND2_X1   g660(.A1(new_n849), .A2(new_n645), .ZN(new_n1087));
  INV_X1    g661(.A(G319), .ZN(new_n1088));
  NOR2_X1   g662(.A1(G227), .A2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g663(.A(new_n1089), .B(KEYINPUT127), .Z(new_n1090));
  AND4_X1   g664(.A1(new_n1086), .A2(new_n913), .A3(new_n1087), .A4(new_n1090), .ZN(G308));
  NAND4_X1  g665(.A1(new_n913), .A2(new_n1086), .A3(new_n1087), .A4(new_n1090), .ZN(G225));
endmodule


