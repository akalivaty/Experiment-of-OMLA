//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT79), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT78), .ZN(new_n193));
  INV_X1    g007(.A(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G125), .ZN(new_n195));
  INV_X1    g009(.A(G125), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G140), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n197), .A3(KEYINPUT16), .ZN(new_n198));
  OR3_X1    g012(.A1(new_n196), .A2(KEYINPUT16), .A3(G140), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n193), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n196), .A2(KEYINPUT16), .A3(G140), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT78), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n192), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n202), .ZN(new_n204));
  XNOR2_X1  g018(.A(G125), .B(G140), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n201), .B1(new_n205), .B2(KEYINPUT16), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n204), .B(G146), .C1(new_n206), .C2(new_n193), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G119), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT24), .B(G110), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n211), .B2(G128), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n212), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G110), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT77), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(KEYINPUT77), .A3(G110), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n215), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n208), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n213), .A2(new_n214), .ZN(new_n226));
  INV_X1    g040(.A(G110), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n217), .A2(new_n218), .A3(new_n227), .A4(new_n212), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n226), .A2(new_n228), .B1(new_n192), .B2(new_n205), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n207), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n191), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT80), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n208), .A2(new_n224), .B1(new_n207), .B2(new_n229), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n231), .A2(new_n232), .B1(new_n233), .B2(new_n190), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT80), .B1(new_n233), .B2(new_n191), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G217), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(G234), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(G902), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n240), .B(KEYINPUT81), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT82), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n225), .A2(new_n230), .ZN(new_n245));
  INV_X1    g059(.A(new_n191), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n232), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n233), .A2(new_n190), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n247), .A2(new_n235), .A3(new_n238), .A4(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT25), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n234), .A2(KEYINPUT25), .A3(new_n238), .A4(new_n235), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n239), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  OR2_X1    g069(.A1(new_n244), .A2(new_n255), .ZN(new_n256));
  XOR2_X1   g070(.A(G116), .B(G119), .Z(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT2), .B(G113), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XOR2_X1   g073(.A(KEYINPUT2), .B(G113), .Z(new_n260));
  XNOR2_X1  g074(.A(G116), .B(G119), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(G143), .B(G146), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT65), .B1(new_n266), .B2(G146), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(new_n192), .A3(G143), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(G146), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT1), .B1(new_n266), .B2(G146), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G128), .ZN(new_n273));
  AOI221_X4 g087(.A(KEYINPUT69), .B1(new_n264), .B2(new_n265), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n273), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n264), .A2(new_n265), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G134), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G137), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n280), .A2(G137), .ZN(new_n283));
  OAI21_X1  g097(.A(G131), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT11), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n280), .B2(G137), .ZN(new_n286));
  INV_X1    g100(.A(G137), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT11), .A3(G134), .ZN(new_n288));
  INV_X1    g102(.A(G131), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n286), .A2(new_n288), .A3(new_n289), .A4(new_n281), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n263), .B1(new_n279), .B2(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(KEYINPUT0), .A2(G128), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT0), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n209), .A3(KEYINPUT64), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT64), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(KEYINPUT0), .B2(G128), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n294), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n271), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n264), .A2(new_n294), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT67), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n286), .A2(new_n288), .A3(new_n281), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G131), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n290), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n299), .A2(new_n271), .B1(new_n264), .B2(new_n294), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT67), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n303), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT28), .B1(new_n293), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT26), .B(G101), .Z(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(G237), .A2(G953), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G210), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n315), .B(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n321), .A2(KEYINPUT29), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT68), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n310), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n303), .A2(KEYINPUT68), .A3(new_n306), .A4(new_n309), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n293), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT70), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n324), .A2(new_n293), .A3(KEYINPUT70), .A4(new_n325), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n329), .B1(new_n328), .B2(new_n330), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n279), .A2(new_n292), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n324), .A2(new_n333), .A3(new_n325), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n263), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n331), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n312), .B(new_n322), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n328), .A2(new_n330), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n192), .A2(G143), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n265), .A2(new_n341), .A3(new_n270), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n342), .B1(new_n271), .B2(new_n273), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(new_n291), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n302), .A2(KEYINPUT66), .B1(new_n290), .B2(new_n305), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT66), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n307), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n344), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n348), .A2(KEYINPUT30), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n324), .A2(KEYINPUT30), .A3(new_n333), .A4(new_n325), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n263), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n340), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT29), .B1(new_n352), .B2(new_n320), .ZN(new_n353));
  INV_X1    g167(.A(new_n263), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT75), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT75), .ZN(new_n356));
  INV_X1    g170(.A(new_n347), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n306), .B1(new_n307), .B2(new_n346), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n356), .B(new_n263), .C1(new_n359), .C2(new_n344), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(new_n328), .B2(new_n330), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n321), .B(new_n312), .C1(new_n362), .C2(new_n338), .ZN(new_n363));
  AOI21_X1  g177(.A(G902), .B1(new_n353), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n339), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n340), .A2(new_n321), .A3(new_n351), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT31), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT74), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n361), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n338), .B1(new_n340), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n320), .B1(new_n371), .B2(new_n311), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n366), .A2(KEYINPUT74), .A3(KEYINPUT31), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT31), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n340), .A2(new_n374), .A3(new_n321), .A4(new_n351), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n369), .A2(new_n372), .A3(new_n373), .A4(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(G472), .A2(G902), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT32), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n365), .A2(G472), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n377), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n379), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n256), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT9), .B(G234), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(KEYINPUT83), .ZN(new_n386));
  OAI21_X1  g200(.A(G221), .B1(new_n386), .B2(G902), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G469), .ZN(new_n389));
  XNOR2_X1  g203(.A(G110), .B(G140), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n188), .A2(G227), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n390), .B(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G104), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT3), .B1(new_n393), .B2(G107), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT3), .ZN(new_n395));
  INV_X1    g209(.A(G107), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n396), .A3(G104), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n393), .A2(G107), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n399), .A2(G101), .ZN(new_n400));
  INV_X1    g214(.A(G101), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n394), .A2(new_n397), .A3(new_n401), .A4(new_n398), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT4), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT85), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n399), .A2(G101), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT85), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT4), .A4(new_n402), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n399), .A2(new_n409), .A3(G101), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n303), .A2(new_n309), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n276), .A2(new_n277), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT69), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n276), .A2(new_n275), .A3(new_n277), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n393), .A2(G107), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n396), .A2(G104), .ZN(new_n417));
  OAI21_X1  g231(.A(G101), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n402), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n414), .A2(KEYINPUT10), .A3(new_n415), .A4(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n264), .B1(G128), .B2(new_n272), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n402), .B(new_n418), .C1(new_n422), .C2(new_n342), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT86), .B(KEYINPUT10), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT87), .B1(new_n412), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n404), .A2(new_n407), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n428), .A2(new_n303), .A3(new_n309), .A4(new_n410), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n420), .A2(KEYINPUT10), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n279), .A2(new_n430), .B1(new_n423), .B2(new_n424), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT87), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n427), .A2(new_n306), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n306), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n429), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n392), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n419), .A2(new_n276), .A3(new_n277), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n423), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n306), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT12), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(KEYINPUT12), .A3(new_n306), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n436), .A2(new_n392), .A3(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n389), .B(new_n238), .C1(new_n437), .C2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n392), .B(KEYINPUT84), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n436), .B2(new_n444), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n436), .A2(new_n392), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n434), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G469), .B1(new_n450), .B2(G902), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n388), .B1(new_n446), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G116), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G122), .ZN(new_n454));
  INV_X1    g268(.A(G122), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G116), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n456), .A3(new_n396), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n209), .A2(G143), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n266), .A2(G128), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n280), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n280), .B1(new_n458), .B2(new_n459), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n457), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n454), .A2(new_n456), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(KEYINPUT14), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT14), .ZN(new_n466));
  OAI21_X1  g280(.A(G107), .B1(new_n454), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT92), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n454), .A2(new_n456), .A3(new_n396), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n396), .B1(new_n454), .B2(new_n456), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n464), .A2(G107), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(KEYINPUT92), .A3(new_n457), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n461), .A2(KEYINPUT95), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT95), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n460), .A2(new_n477), .ZN(new_n478));
  AND4_X1   g292(.A1(new_n473), .A2(new_n475), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n266), .A2(KEYINPUT13), .A3(G128), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT93), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT13), .B1(new_n266), .B2(G128), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n459), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT93), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n484), .A3(new_n459), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G134), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT94), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n482), .A2(new_n459), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(KEYINPUT93), .A3(new_n480), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT94), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n489), .A2(new_n490), .A3(G134), .A4(new_n485), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n469), .B1(new_n479), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n188), .A2(G217), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n386), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  AOI211_X1 g311(.A(new_n469), .B(new_n495), .C1(new_n479), .C2(new_n492), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n238), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT96), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G478), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(KEYINPUT15), .ZN(new_n503));
  OAI211_X1 g317(.A(KEYINPUT96), .B(new_n238), .C1(new_n497), .C2(new_n498), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n499), .A2(new_n503), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT20), .ZN(new_n508));
  XNOR2_X1  g322(.A(G113), .B(G122), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(new_n393), .ZN(new_n510));
  INV_X1    g324(.A(G237), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n188), .A3(G214), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n266), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n316), .A2(G143), .A3(G214), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(KEYINPUT18), .A2(G131), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n195), .A2(new_n197), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n205), .A2(KEYINPUT89), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n521), .A3(G146), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(G146), .B2(new_n518), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n515), .A2(KEYINPUT91), .A3(G131), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT91), .B1(new_n515), .B2(G131), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT17), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n203), .A3(new_n207), .ZN(new_n529));
  INV_X1    g343(.A(new_n514), .ZN(new_n530));
  AOI21_X1  g344(.A(G143), .B1(new_n316), .B2(G214), .ZN(new_n531));
  OAI21_X1  g345(.A(G131), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT91), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT90), .B1(new_n515), .B2(G131), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT90), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n513), .A2(new_n536), .A3(new_n289), .A4(new_n514), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n534), .A2(new_n535), .A3(new_n525), .A4(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(KEYINPUT17), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n510), .B(new_n524), .C1(new_n529), .C2(new_n539), .ZN(new_n540));
  AND4_X1   g354(.A1(new_n534), .A2(new_n535), .A3(new_n525), .A4(new_n537), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT19), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n518), .A2(KEYINPUT19), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n207), .B1(new_n544), .B2(G146), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n524), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n510), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(G475), .A2(G902), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n508), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n550), .ZN(new_n552));
  AOI211_X1 g366(.A(KEYINPUT20), .B(new_n552), .C1(new_n540), .C2(new_n548), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n524), .B1(new_n529), .B2(new_n539), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n547), .ZN(new_n555));
  AOI21_X1  g369(.A(G902), .B1(new_n555), .B2(new_n540), .ZN(new_n556));
  INV_X1    g370(.A(G475), .ZN(new_n557));
  OAI22_X1  g371(.A1(new_n551), .A2(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n507), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n452), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n263), .A2(new_n410), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n428), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT5), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(new_n211), .A3(G116), .ZN(new_n565));
  OAI211_X1 g379(.A(G113), .B(new_n565), .C1(new_n257), .C2(new_n564), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n420), .A2(new_n262), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(G110), .B(G122), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n568), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n561), .B1(new_n404), .B2(new_n407), .ZN(new_n571));
  INV_X1    g385(.A(new_n567), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(KEYINPUT6), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT6), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n575), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n307), .A2(G125), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(G125), .B2(new_n343), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n188), .A2(G224), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(KEYINPUT88), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n578), .B(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n574), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(KEYINPUT7), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n583), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n577), .B(new_n585), .C1(G125), .C2(new_n343), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n566), .A2(new_n262), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n419), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n567), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n568), .B(KEYINPUT8), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n584), .A2(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(G902), .B1(new_n591), .B2(new_n569), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n582), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(G210), .B1(G237), .B2(G902), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n582), .A2(new_n594), .A3(new_n592), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n188), .A2(G952), .ZN(new_n599));
  NAND2_X1  g413(.A1(G234), .A2(G237), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(G902), .A3(G953), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT21), .B(G898), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G214), .B1(G237), .B2(G902), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n598), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n560), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n384), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  AND2_X1   g426(.A1(new_n376), .A2(new_n377), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n244), .A2(new_n255), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n452), .ZN(new_n615));
  INV_X1    g429(.A(G472), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n376), .B2(new_n238), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n613), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n479), .A2(new_n492), .ZN(new_n619));
  INV_X1    g433(.A(new_n469), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n620), .A3(new_n496), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n619), .A2(new_n620), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n495), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n493), .A2(KEYINPUT98), .A3(new_n496), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n623), .A2(new_n625), .A3(KEYINPUT33), .A4(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT97), .B(KEYINPUT33), .Z(new_n628));
  OAI21_X1  g442(.A(new_n628), .B1(new_n497), .B2(new_n498), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n502), .A2(G902), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n627), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT99), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n627), .A2(new_n634), .A3(new_n629), .A4(new_n630), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n558), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n609), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n618), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G104), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  INV_X1    g456(.A(new_n558), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n507), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n609), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n618), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NOR2_X1   g462(.A1(new_n613), .A2(new_n617), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n246), .A2(KEYINPUT36), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n233), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n233), .A2(new_n652), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n651), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n655), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n657), .A2(new_n650), .A3(new_n653), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n253), .A2(new_n239), .B1(new_n659), .B2(new_n241), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n560), .A2(new_n609), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n649), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  NAND2_X1  g478(.A1(new_n381), .A2(new_n383), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n446), .A2(new_n451), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n387), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n659), .A2(new_n241), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n254), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n608), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n596), .B2(new_n597), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n603), .A2(G900), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n601), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n643), .A2(new_n507), .A3(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n667), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n665), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XNOR2_X1  g492(.A(new_n674), .B(KEYINPUT39), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n452), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n680), .A2(new_n681), .ZN(new_n684));
  OAI21_X1  g498(.A(KEYINPUT40), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n684), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT40), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n687), .A3(new_n682), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n376), .A2(new_n380), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n352), .A2(new_n321), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n336), .B1(new_n340), .B2(KEYINPUT76), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n238), .B(new_n690), .C1(new_n693), .C2(new_n321), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G472), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n383), .A2(new_n689), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT38), .B1(new_n596), .B2(new_n597), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n596), .A2(KEYINPUT38), .A3(new_n597), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n507), .A2(new_n558), .A3(new_n608), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n700), .A2(new_n669), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n685), .A2(new_n688), .A3(new_n696), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  NAND3_X1  g518(.A1(new_n636), .A2(new_n558), .A3(new_n674), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n667), .A2(new_n672), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n665), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  OAI21_X1  g522(.A(new_n238), .B1(new_n437), .B2(new_n445), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G469), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n387), .A3(new_n446), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n256), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n665), .A2(new_n638), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND3_X1  g529(.A1(new_n665), .A2(new_n645), .A3(new_n712), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  NAND4_X1  g531(.A1(new_n710), .A2(new_n671), .A3(new_n387), .A4(new_n446), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n559), .A2(new_n607), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n718), .A2(new_n719), .A3(new_n660), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n665), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  AOI21_X1  g536(.A(new_n338), .B1(new_n691), .B2(new_n692), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n320), .B1(new_n723), .B2(new_n311), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n367), .A2(new_n375), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n378), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n617), .A2(new_n726), .A3(new_n256), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n710), .A2(new_n607), .A3(new_n387), .A4(new_n446), .ZN(new_n728));
  INV_X1    g542(.A(new_n597), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n594), .B1(new_n582), .B2(new_n592), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT103), .B1(new_n701), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n670), .B1(new_n505), .B2(new_n506), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n598), .A3(new_n734), .A4(new_n558), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n728), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n727), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR2_X1   g552(.A1(new_n617), .A2(new_n726), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n718), .A2(new_n660), .A3(new_n705), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  NOR3_X1   g556(.A1(new_n729), .A2(new_n730), .A3(new_n670), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n452), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n705), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n384), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n384), .A2(KEYINPUT42), .A3(new_n745), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G131), .ZN(G33));
  NOR2_X1   g565(.A1(new_n744), .A2(new_n675), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n384), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G134), .ZN(G36));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n649), .B2(new_n660), .ZN(new_n756));
  OAI211_X1 g570(.A(KEYINPUT105), .B(new_n669), .C1(new_n613), .C2(new_n617), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n558), .A2(KEYINPUT104), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT104), .ZN(new_n760));
  OAI221_X1 g574(.A(new_n760), .B1(new_n556), .B2(new_n557), .C1(new_n551), .C2(new_n553), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n761), .A3(new_n636), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT43), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n558), .A2(KEYINPUT43), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n636), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n758), .A2(KEYINPUT44), .A3(new_n767), .ZN(new_n771));
  NAND2_X1  g585(.A1(G469), .A2(G902), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n450), .A2(KEYINPUT45), .ZN(new_n773));
  OAI21_X1  g587(.A(G469), .B1(new_n450), .B2(KEYINPUT45), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(KEYINPUT46), .B(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n446), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n387), .A3(new_n679), .ZN(new_n780));
  INV_X1    g594(.A(new_n743), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n770), .A2(new_n771), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  NOR4_X1   g598(.A1(new_n665), .A2(new_n614), .A3(new_n705), .A4(new_n781), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n779), .A2(new_n387), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n779), .A2(KEYINPUT47), .A3(new_n387), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  NOR2_X1   g606(.A1(G952), .A2(G953), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n638), .A2(KEYINPUT106), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT106), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n609), .B2(new_n637), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n795), .B(new_n797), .C1(new_n609), .C2(new_n644), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n618), .A2(new_n798), .B1(new_n727), .B2(new_n736), .ZN(new_n799));
  AOI22_X1  g613(.A1(new_n720), .A2(new_n665), .B1(new_n649), .B2(new_n661), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n665), .B(new_n712), .C1(new_n638), .C2(new_n645), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n799), .A2(new_n611), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n384), .A2(KEYINPUT42), .A3(new_n745), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT42), .B1(new_n384), .B2(new_n745), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n617), .A2(new_n726), .A3(new_n660), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n745), .ZN(new_n807));
  INV_X1    g621(.A(new_n674), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n507), .A2(new_n558), .A3(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(new_n452), .A3(new_n669), .A4(new_n743), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT107), .B1(new_n665), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT107), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n813), .B(new_n810), .C1(new_n381), .C2(new_n383), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n753), .B(new_n807), .C1(new_n812), .C2(new_n814), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n802), .A2(new_n805), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n365), .A2(G472), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n689), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT32), .B1(new_n376), .B2(new_n377), .ZN(new_n819));
  OAI22_X1  g633(.A1(new_n818), .A2(new_n819), .B1(new_n676), .B2(new_n706), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n660), .A2(new_n674), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT108), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n821), .B(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n667), .B1(new_n732), .B2(new_n735), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n689), .A2(new_n695), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n823), .B(new_n824), .C1(new_n825), .C2(new_n819), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n820), .A2(new_n741), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT52), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n820), .A2(new_n826), .A3(new_n829), .A4(new_n741), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT53), .B1(new_n816), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n812), .ZN(new_n834));
  INV_X1    g648(.A(new_n814), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n753), .A2(new_n807), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n750), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n839), .A2(new_n831), .A3(new_n840), .A4(new_n802), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n794), .B1(new_n833), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n618), .A2(new_n798), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n801), .A2(new_n843), .A3(new_n737), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n800), .A2(new_n611), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n815), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n750), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n840), .B1(new_n848), .B2(new_n831), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n816), .A2(KEYINPUT53), .A3(new_n832), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(KEYINPUT54), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n842), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n853));
  AOI221_X4 g667(.A(new_n601), .B1(new_n764), .B2(new_n636), .C1(new_n762), .C2(KEYINPUT43), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n739), .A2(new_n854), .A3(new_n614), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT109), .B1(new_n855), .B2(new_n781), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT109), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n727), .A2(new_n857), .A3(new_n743), .A4(new_n854), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n710), .A2(new_n446), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n860), .A2(new_n388), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n790), .B2(KEYINPUT110), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT110), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n788), .A2(new_n863), .A3(new_n789), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n859), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n710), .A2(new_n743), .A3(new_n387), .A4(new_n446), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT112), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n763), .A2(new_n602), .A3(new_n765), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n860), .A2(KEYINPUT112), .A3(new_n387), .A4(new_n743), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT112), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(KEYINPUT113), .A3(new_n854), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n806), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n608), .B1(new_n698), .B2(new_n699), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT111), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n860), .A3(new_n879), .A4(new_n387), .ZN(new_n880));
  INV_X1    g694(.A(new_n699), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n670), .B1(new_n881), .B2(new_n697), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT111), .B1(new_n882), .B2(new_n711), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(KEYINPUT50), .A3(new_n727), .A4(new_n854), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT50), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n880), .A2(new_n883), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n886), .B1(new_n855), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n696), .A2(new_n256), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n601), .B1(new_n871), .B2(new_n873), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n636), .A2(new_n558), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n877), .A2(new_n889), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n853), .B1(new_n865), .B2(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n890), .A2(new_n891), .ZN(new_n896));
  AOI22_X1  g710(.A1(new_n896), .A2(new_n892), .B1(new_n876), .B2(new_n806), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n856), .B(new_n858), .C1(new_n790), .C2(new_n861), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(KEYINPUT51), .A3(new_n889), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT48), .B1(new_n876), .B2(new_n384), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT48), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n665), .A2(new_n614), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n902), .B(new_n903), .C1(new_n870), .C2(new_n875), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n825), .A2(new_n819), .ZN(new_n906));
  INV_X1    g720(.A(new_n637), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n891), .A2(new_n614), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n718), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n727), .A2(new_n909), .A3(new_n854), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n599), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT114), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT114), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n908), .A2(new_n913), .A3(new_n599), .A4(new_n910), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT115), .B1(new_n905), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n905), .A2(new_n915), .A3(KEYINPUT115), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n900), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n793), .B1(new_n852), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n860), .B(KEYINPUT49), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n762), .A2(new_n670), .A3(new_n388), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n890), .A2(new_n700), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(KEYINPUT116), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT116), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n905), .A2(KEYINPUT115), .A3(new_n915), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n895), .B(new_n899), .C1(new_n927), .C2(new_n916), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n842), .B2(new_n851), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n926), .B(new_n923), .C1(new_n929), .C2(new_n793), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n930), .ZN(G75));
  AOI21_X1  g745(.A(new_n238), .B1(new_n849), .B2(new_n850), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(G210), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n574), .A2(new_n576), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n581), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT55), .ZN(new_n936));
  XOR2_X1   g750(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n937));
  AND3_X1   g751(.A1(new_n933), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT56), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n936), .B1(new_n933), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n188), .A2(G952), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n938), .A2(new_n940), .A3(new_n941), .ZN(G51));
  NOR2_X1   g756(.A1(new_n773), .A2(new_n774), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT118), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n932), .A2(KEYINPUT119), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT119), .B1(new_n932), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n772), .B(KEYINPUT57), .ZN(new_n948));
  OAI22_X1  g762(.A1(new_n852), .A2(new_n948), .B1(new_n437), .B2(new_n445), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n941), .B1(new_n947), .B2(new_n949), .ZN(G54));
  NAND3_X1  g764(.A1(new_n932), .A2(KEYINPUT58), .A3(G475), .ZN(new_n951));
  INV_X1    g765(.A(new_n549), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n951), .A2(KEYINPUT120), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n941), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n951), .B2(new_n952), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT120), .B1(new_n951), .B2(new_n952), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(G60));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT59), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n842), .A2(new_n851), .A3(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n627), .A2(new_n629), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n954), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n960), .B2(new_n962), .ZN(G63));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT60), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(new_n849), .B2(new_n850), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n967), .A2(new_n236), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n941), .B1(new_n967), .B2(new_n659), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT121), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n967), .B2(new_n659), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n972), .A2(KEYINPUT61), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n968), .B(new_n969), .C1(new_n972), .C2(KEYINPUT61), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(G66));
  INV_X1    g790(.A(G224), .ZN(new_n977));
  OAI21_X1  g791(.A(G953), .B1(new_n605), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n846), .B2(G953), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n934), .B1(G898), .B2(new_n188), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(G69));
  NAND2_X1  g795(.A1(new_n349), .A2(new_n350), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT122), .Z(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(new_n544), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT123), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n781), .B1(new_n644), .B2(new_n637), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n384), .A2(new_n682), .A3(new_n686), .A4(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n820), .A2(new_n741), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n703), .A2(new_n988), .A3(KEYINPUT62), .ZN(new_n989));
  AOI21_X1  g803(.A(KEYINPUT62), .B1(new_n703), .B2(new_n988), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n791), .B(new_n987), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n770), .A2(new_n771), .A3(new_n782), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n985), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n791), .A2(new_n987), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n703), .A2(new_n988), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT62), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n703), .A2(new_n988), .A3(KEYINPUT62), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n994), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(KEYINPUT123), .A3(new_n783), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n993), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n984), .B1(new_n1001), .B2(G953), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT124), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT126), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n732), .A2(new_n735), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n384), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(KEYINPUT125), .B1(new_n1008), .B2(new_n780), .ZN(new_n1009));
  INV_X1    g823(.A(new_n780), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT125), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1010), .A2(new_n1011), .A3(new_n384), .A4(new_n1007), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g827(.A1(new_n785), .A2(new_n790), .B1(new_n384), .B2(new_n752), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1013), .A2(new_n1014), .A3(new_n750), .A4(new_n988), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1006), .B1(new_n992), .B2(new_n1015), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n1014), .A2(new_n750), .A3(new_n988), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1017), .A2(new_n783), .A3(KEYINPUT126), .A4(new_n1013), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1016), .A2(new_n188), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n984), .B1(G900), .B2(G953), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .A4(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(G953), .B1(new_n993), .B2(new_n1000), .ZN(new_n1023));
  INV_X1    g837(.A(new_n984), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1003), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1021), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1004), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1022), .A2(new_n1027), .ZN(G72));
  NAND3_X1  g842(.A1(new_n1016), .A2(new_n846), .A3(new_n1018), .ZN(new_n1029));
  NAND2_X1  g843(.A1(G472), .A2(G902), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT63), .Z(new_n1031));
  NAND2_X1  g845(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n352), .A2(new_n321), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n833), .A2(new_n841), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(new_n690), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1031), .ZN(new_n1038));
  NOR3_X1   g852(.A1(new_n1037), .A2(new_n1033), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n941), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1034), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n993), .A2(new_n846), .A3(new_n1000), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1042), .A2(new_n1031), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(new_n1037), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1044), .A2(KEYINPUT127), .ZN(new_n1045));
  INV_X1    g859(.A(KEYINPUT127), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1043), .A2(new_n1046), .A3(new_n1037), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1041), .B1(new_n1045), .B2(new_n1047), .ZN(G57));
endmodule


