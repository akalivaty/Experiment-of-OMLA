//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT66), .B(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n465), .B(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n462), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  OR2_X1    g047(.A1(G100), .A2(G2105), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n473), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT68), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT3), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n475), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND3_X1  g061(.A1(new_n477), .A2(new_n479), .A3(G126), .ZN(new_n487));
  NAND2_X1  g062(.A1(G114), .A2(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n476), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G102), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n477), .A2(new_n479), .A3(G138), .A4(new_n462), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n463), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n490), .A2(new_n492), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT69), .A3(G543), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n501), .A2(new_n503), .B1(KEYINPUT5), .B2(new_n500), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(G543), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n507), .A2(new_n513), .ZN(G166));
  AND2_X1   g089(.A1(new_n508), .A2(G543), .ZN(new_n515));
  XOR2_X1   g090(.A(KEYINPUT70), .B(G51), .Z(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND3_X1   g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  INV_X1    g093(.A(G89), .ZN(new_n519));
  OAI221_X1 g094(.A(new_n517), .B1(KEYINPUT7), .B2(new_n518), .C1(new_n519), .C2(new_n509), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n504), .A2(G63), .ZN(new_n521));
  NAND3_X1  g096(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n506), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n520), .A2(new_n523), .ZN(G168));
  AOI22_X1  g099(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n506), .ZN(new_n526));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  INV_X1    g102(.A(G52), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n509), .A2(new_n527), .B1(new_n528), .B2(new_n512), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n526), .A2(new_n529), .ZN(G301));
  INV_X1    g105(.A(G301), .ZN(G171));
  AOI22_X1  g106(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(new_n506), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n515), .A2(G43), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n504), .A2(G81), .A3(new_n508), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n535), .B1(new_n534), .B2(new_n536), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n533), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT72), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT72), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n533), .B(new_n541), .C1(new_n537), .C2(new_n538), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT73), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(G188));
  INV_X1    g125(.A(G53), .ZN(new_n551));
  OAI211_X1 g126(.A(KEYINPUT74), .B(KEYINPUT9), .C1(new_n512), .C2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n554));
  AND4_X1   g129(.A1(G53), .A2(new_n508), .A3(G543), .A4(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT75), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n555), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n557), .A2(new_n552), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n501), .A2(new_n503), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n566), .A2(KEYINPUT76), .A3(G651), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n504), .A2(new_n508), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G91), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n560), .A2(new_n571), .A3(new_n573), .ZN(G299));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(G166), .ZN(G303));
  AOI22_X1  g151(.A1(new_n572), .A2(G87), .B1(G49), .B2(new_n515), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g155(.A(KEYINPUT77), .B(G651), .C1(new_n504), .C2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n577), .A2(new_n580), .A3(new_n581), .ZN(G288));
  NAND4_X1  g157(.A1(new_n562), .A2(G86), .A3(new_n563), .A4(new_n508), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n515), .A2(G48), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n506), .ZN(G305));
  AOI22_X1  g161(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT78), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  XNOR2_X1  g164(.A(KEYINPUT79), .B(G85), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n572), .A2(new_n590), .B1(G47), .B2(new_n515), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n572), .A2(KEYINPUT81), .A3(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n509), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n595), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n596), .B1(new_n595), .B2(new_n599), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n594), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n602), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n600), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n564), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n515), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n603), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(KEYINPUT82), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n603), .A2(new_n605), .A3(new_n612), .A4(new_n609), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n593), .B1(new_n615), .B2(G868), .ZN(G284));
  OAI21_X1  g191(.A(new_n593), .B1(new_n615), .B2(G868), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(G299), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G297));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND3_X1  g198(.A1(new_n611), .A2(new_n622), .A3(new_n613), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n463), .A2(new_n491), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g205(.A(G2100), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n481), .A2(G123), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n483), .A2(G135), .ZN(new_n634));
  NOR2_X1   g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n632), .A2(new_n638), .ZN(G156));
  XOR2_X1   g214(.A(KEYINPUT85), .B(G2438), .Z(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT15), .B(G2435), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT84), .B(KEYINPUT14), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2451), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n650), .A2(new_n651), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n650), .A2(new_n651), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(G14), .A3(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT86), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n662), .A2(new_n663), .ZN(new_n668));
  INV_X1    g243(.A(new_n664), .ZN(new_n669));
  INV_X1    g244(.A(new_n662), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n663), .B(KEYINPUT17), .Z(new_n671));
  OAI211_X1 g246(.A(new_n668), .B(new_n669), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n670), .A2(new_n671), .A3(new_n664), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n667), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2096), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n631), .ZN(G227));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n678), .A2(new_n681), .A3(new_n683), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n686), .B(new_n687), .C1(new_n685), .C2(new_n684), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(G1986), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT22), .B(G1981), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G229));
  NAND2_X1  g269(.A1(new_n481), .A2(G119), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n483), .A2(G131), .ZN(new_n696));
  NOR2_X1   g271(.A1(G95), .A2(G2105), .ZN(new_n697));
  OAI21_X1  g272(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n695), .B(new_n696), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT87), .B(G29), .ZN(new_n700));
  MUX2_X1   g275(.A(G25), .B(new_n699), .S(new_n700), .Z(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT35), .B(G1991), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  AND2_X1   g278(.A1(KEYINPUT88), .A2(G16), .ZN(new_n704));
  NOR2_X1   g279(.A1(KEYINPUT88), .A2(G16), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(G290), .A2(KEYINPUT89), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT89), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n589), .A2(new_n709), .A3(new_n591), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n707), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n706), .A2(G24), .ZN(new_n712));
  OR3_X1    g287(.A1(new_n711), .A2(G1986), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(G1986), .B1(new_n711), .B2(new_n712), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n703), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(G166), .A2(new_n707), .ZN(new_n716));
  INV_X1    g291(.A(G22), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n706), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(G1971), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G1971), .ZN(new_n720));
  INV_X1    g295(.A(new_n718), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n720), .B(new_n721), .C1(G166), .C2(new_n707), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G6), .A2(G16), .ZN(new_n724));
  INV_X1    g299(.A(G48), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n583), .B1(new_n725), .B2(new_n512), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n562), .A2(G61), .A3(new_n563), .ZN(new_n727));
  NAND2_X1  g302(.A1(G73), .A2(G543), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n506), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n724), .B1(new_n730), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT32), .B(G1981), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n577), .A2(G16), .A3(new_n580), .A4(new_n581), .ZN(new_n735));
  OR2_X1    g310(.A1(G16), .A2(G23), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT33), .B(G1976), .Z(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n735), .B2(new_n736), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n723), .A2(new_n734), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n719), .B(new_n722), .C1(new_n739), .C2(new_n740), .ZN(new_n744));
  OAI21_X1  g319(.A(KEYINPUT90), .B1(new_n744), .B2(new_n733), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT34), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n743), .A2(new_n745), .A3(KEYINPUT34), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n715), .A2(new_n748), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(KEYINPUT91), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT91), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n715), .A2(new_n748), .A3(new_n753), .A4(new_n750), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n752), .A2(KEYINPUT36), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n751), .A2(KEYINPUT91), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT97), .ZN(new_n759));
  OAI21_X1  g334(.A(G16), .B1(new_n520), .B2(new_n523), .ZN(new_n760));
  INV_X1    g335(.A(G16), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G21), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n759), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n760), .A2(new_n759), .A3(new_n762), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n764), .A2(G1966), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT98), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n707), .B1(new_n540), .B2(new_n542), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n706), .A2(G19), .ZN(new_n769));
  OR3_X1    g344(.A1(new_n768), .A2(G1341), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(G1341), .B1(new_n768), .B2(new_n769), .ZN(new_n771));
  INV_X1    g346(.A(new_n700), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G27), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G164), .B2(new_n772), .ZN(new_n774));
  MUX2_X1   g349(.A(new_n773), .B(new_n774), .S(KEYINPUT99), .Z(new_n775));
  AOI22_X1  g350(.A1(new_n770), .A2(new_n771), .B1(G2078), .B2(new_n775), .ZN(new_n776));
  OAI22_X1  g351(.A1(new_n775), .A2(G2078), .B1(new_n637), .B2(new_n772), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n772), .A2(G35), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G162), .B2(new_n772), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT29), .B(G2090), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G1966), .ZN(new_n783));
  INV_X1    g358(.A(new_n765), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n763), .ZN(new_n785));
  INV_X1    g360(.A(G34), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n700), .B1(KEYINPUT24), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT96), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n786), .A2(KEYINPUT24), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n788), .A2(new_n789), .B1(G160), .B2(G29), .ZN(new_n790));
  INV_X1    g365(.A(G2084), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n483), .A2(G141), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n481), .A2(G129), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n491), .A2(G105), .ZN(new_n796));
  NAND3_X1  g371(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT26), .Z(new_n798));
  NAND4_X1  g373(.A1(new_n794), .A2(new_n795), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G29), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G29), .B2(G32), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT27), .B(G1996), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n792), .A2(new_n793), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G5), .A2(G16), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G171), .B2(G16), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G1961), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT31), .B(G11), .ZN(new_n808));
  AND4_X1   g383(.A1(new_n785), .A2(new_n804), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n767), .A2(new_n776), .A3(new_n782), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n707), .A2(G20), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT100), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT23), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n619), .B2(new_n761), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT101), .B(G1956), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G33), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(G29), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT25), .Z(new_n820));
  NAND2_X1  g395(.A1(new_n483), .A2(G139), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n820), .B(new_n821), .C1(new_n462), .C2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT95), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n818), .B1(new_n824), .B2(G29), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G2072), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT30), .B(G28), .Z(new_n827));
  OAI221_X1 g402(.A(new_n826), .B1(G29), .B2(new_n827), .C1(new_n802), .C2(new_n803), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n481), .A2(G128), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n483), .A2(G140), .ZN(new_n830));
  NOR2_X1   g405(.A1(G104), .A2(G2105), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n829), .B(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n772), .A2(G26), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n833), .A2(G29), .B1(KEYINPUT28), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(KEYINPUT28), .B2(new_n834), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G2067), .ZN(new_n837));
  NOR4_X1   g412(.A1(new_n810), .A2(new_n816), .A3(new_n828), .A4(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n806), .A2(G1961), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n758), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT93), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G4), .B2(G16), .ZN(new_n842));
  OR3_X1    g417(.A1(new_n841), .A2(G4), .A3(G16), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n842), .B(new_n843), .C1(new_n614), .C2(new_n761), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(KEYINPUT94), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(KEYINPUT94), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G1348), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n845), .A2(G1348), .A3(new_n846), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n756), .A2(new_n840), .A3(new_n851), .ZN(G311));
  INV_X1    g427(.A(new_n851), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n758), .A2(new_n838), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n853), .A2(new_n854), .A3(new_n839), .A4(new_n755), .ZN(G150));
  AOI22_X1  g430(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(new_n506), .ZN(new_n857));
  INV_X1    g432(.A(G93), .ZN(new_n858));
  INV_X1    g433(.A(G55), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n509), .A2(new_n858), .B1(new_n859), .B2(new_n512), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G860), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT37), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n615), .A2(G559), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT39), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n861), .B1(new_n540), .B2(new_n542), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n539), .A2(new_n861), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n866), .B(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n864), .B1(new_n873), .B2(G860), .ZN(G145));
  NAND2_X1  g449(.A1(new_n481), .A2(G130), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n483), .A2(G142), .ZN(new_n876));
  NOR2_X1   g451(.A1(G106), .A2(G2105), .ZN(new_n877));
  OAI21_X1  g452(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n875), .B(new_n876), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n699), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT104), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n629), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n880), .B(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n629), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n824), .B(new_n833), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n799), .B(new_n497), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n887), .A2(new_n888), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n637), .B(KEYINPUT103), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(G160), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(G162), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n882), .A2(new_n886), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n891), .A2(new_n892), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n887), .A2(new_n892), .A3(new_n891), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT105), .ZN(new_n902));
  AOI21_X1  g477(.A(G37), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n901), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n904), .A2(new_n896), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g482(.A1(new_n624), .A2(new_n870), .ZN(new_n908));
  INV_X1    g483(.A(new_n870), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n909), .A2(new_n622), .A3(new_n611), .A4(new_n613), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n610), .A2(G299), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n619), .A2(new_n609), .A3(new_n605), .A4(new_n603), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(new_n912), .B2(new_n913), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n912), .A2(new_n913), .A3(new_n920), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n908), .B(new_n910), .C1(new_n919), .C2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n916), .A2(KEYINPUT106), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n911), .A2(new_n924), .A3(new_n915), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n589), .A2(G288), .A3(new_n591), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(G288), .B1(new_n589), .B2(new_n591), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT108), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(G166), .B(new_n730), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n928), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n934), .A3(new_n926), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n929), .A2(new_n935), .A3(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT42), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n923), .A2(new_n925), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n938), .B1(new_n923), .B2(new_n925), .ZN(new_n940));
  OAI21_X1  g515(.A(G868), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n861), .A2(G868), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(G295));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n942), .ZN(G331));
  INV_X1    g519(.A(new_n937), .ZN(new_n945));
  XNOR2_X1  g520(.A(G168), .B(G301), .ZN(new_n946));
  OR3_X1    g521(.A1(new_n946), .A2(new_n867), .A3(new_n869), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n946), .B1(new_n867), .B2(new_n869), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(new_n921), .B2(new_n919), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n915), .A2(new_n947), .A3(new_n948), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n945), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n914), .A2(new_n920), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n949), .B(new_n955), .C1(new_n914), .C2(new_n918), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n945), .B1(new_n956), .B2(new_n951), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT43), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n950), .A2(new_n951), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n937), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n960), .A2(new_n961), .A3(new_n953), .A4(new_n952), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n958), .A2(KEYINPUT44), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n954), .B2(new_n957), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n960), .A2(KEYINPUT43), .A3(new_n953), .A4(new_n952), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n963), .A2(new_n967), .ZN(G397));
  NAND2_X1  g543(.A1(G305), .A2(G1981), .ZN(new_n969));
  XOR2_X1   g544(.A(KEYINPUT114), .B(G1981), .Z(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT115), .B1(new_n730), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT115), .ZN(new_n973));
  NOR4_X1   g548(.A1(new_n726), .A2(new_n729), .A3(new_n973), .A4(new_n970), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n969), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT49), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n495), .A2(new_n496), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n489), .A2(G2105), .B1(G102), .B2(new_n491), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G40), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n468), .A2(new_n471), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n978), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n973), .B1(G305), .B2(new_n970), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n730), .A2(KEYINPUT115), .A3(new_n971), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(KEYINPUT49), .A3(new_n969), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n977), .A2(new_n984), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n981), .A2(new_n983), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(G8), .ZN(new_n992));
  INV_X1    g567(.A(G1976), .ZN(new_n993));
  NAND2_X1  g568(.A1(G288), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n990), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n577), .A2(G1976), .A3(new_n580), .A4(new_n581), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n984), .A2(KEYINPUT113), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n996), .A2(KEYINPUT113), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n999), .A2(new_n990), .A3(new_n984), .A4(new_n994), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n989), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(G166), .A2(new_n978), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT55), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n464), .A2(new_n467), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(G2105), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n469), .A2(new_n470), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n462), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1008), .A3(G40), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n981), .B2(KEYINPUT45), .ZN(new_n1010));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  AOI211_X1 g586(.A(KEYINPUT112), .B(KEYINPUT45), .C1(new_n497), .C2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n1013));
  INV_X1    g588(.A(new_n488), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n463), .B2(G126), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n492), .B1(new_n1015), .B2(new_n462), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n495), .A2(new_n496), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1011), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1013), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1010), .B1(new_n1012), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G2090), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1018), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(KEYINPUT50), .B(new_n1011), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1009), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1021), .A2(new_n720), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(new_n978), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1002), .A2(new_n1004), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G288), .A2(G1976), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT116), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(new_n977), .B2(new_n988), .ZN(new_n1032));
  INV_X1    g607(.A(new_n987), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n984), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n977), .A2(new_n984), .A3(new_n988), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(new_n998), .A3(new_n1000), .ZN(new_n1036));
  OAI211_X1 g611(.A(KEYINPUT45), .B(new_n1011), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n983), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT112), .B1(new_n981), .B2(KEYINPUT45), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1018), .A2(new_n1013), .A3(new_n1019), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1025), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT50), .B1(new_n497), .B2(new_n1011), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n983), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI22_X1  g619(.A1(new_n1041), .A2(G1971), .B1(G2090), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1004), .B1(new_n1045), .B2(G8), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n791), .B(new_n983), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT45), .B1(new_n497), .B2(new_n1011), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n783), .B1(new_n1038), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(G8), .A3(G168), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1036), .A2(new_n1046), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT63), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1029), .B(new_n1034), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n1050), .B2(G286), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1047), .A2(new_n1049), .A3(G168), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G8), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1055), .B1(new_n1057), .B2(G8), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT62), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G2078), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1062), .B(new_n1010), .C1(new_n1012), .C2(new_n1020), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1038), .A2(new_n1064), .A3(G2078), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(KEYINPUT45), .B2(new_n981), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT124), .B(G1961), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1044), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1065), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1058), .A2(KEYINPUT51), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT62), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1073), .B(new_n1074), .C1(new_n1058), .C2(new_n1056), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1061), .A2(new_n1072), .A3(new_n1075), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1051), .A2(KEYINPUT63), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n989), .B2(new_n1001), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1035), .A2(KEYINPUT117), .A3(new_n998), .A4(new_n1000), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1028), .A2(new_n1004), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1046), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1054), .B1(new_n1078), .B2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n569), .A2(new_n570), .B1(G91), .B2(new_n572), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT57), .B1(new_n557), .B2(new_n552), .ZN(new_n1088));
  AOI22_X1  g663(.A1(G299), .A2(KEYINPUT57), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT56), .B(G2072), .Z(new_n1090));
  XNOR2_X1  g665(.A(new_n1090), .B(KEYINPUT118), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1010), .B(new_n1091), .C1(new_n1012), .C2(new_n1020), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n1026), .A2(G1956), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1096), .A2(KEYINPUT119), .A3(new_n1010), .A4(new_n1091), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1089), .A2(new_n1094), .A3(new_n1095), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  OAI22_X1  g674(.A1(new_n1026), .A2(G1348), .B1(G2067), .B2(new_n991), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n615), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT120), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1089), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .A4(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1099), .B1(new_n1101), .B2(new_n1107), .ZN(new_n1108));
  OAI221_X1 g683(.A(KEYINPUT60), .B1(G2067), .B2(new_n991), .C1(new_n1026), .C2(G1348), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n614), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT60), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1100), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n611), .A2(new_n1113), .A3(new_n613), .A4(new_n1109), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1116), .A2(KEYINPUT123), .A3(new_n1095), .A4(new_n1089), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1098), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(KEYINPUT61), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT61), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1121), .A2(new_n1118), .A3(new_n1098), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1115), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT58), .B(G1341), .Z(new_n1124));
  NAND2_X1  g699(.A1(new_n991), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT121), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1021), .A2(G1996), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1126), .A2(new_n1127), .B1(new_n540), .B2(new_n542), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT59), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1128), .B(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1108), .B1(new_n1123), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1044), .A2(KEYINPUT125), .A3(new_n1068), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT125), .B1(new_n1044), .B2(new_n1068), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT110), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n981), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1018), .A2(KEYINPUT110), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1138), .A2(new_n1139), .A3(new_n1019), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1063), .A2(new_n1064), .B1(new_n1066), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1136), .A2(G301), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT54), .B1(new_n1142), .B2(new_n1071), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1084), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1135), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1141), .A2(new_n1145), .A3(new_n1133), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(G171), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1065), .A2(new_n1067), .A3(G301), .A4(new_n1069), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1147), .A2(KEYINPUT126), .A3(KEYINPUT54), .A4(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n1150));
  AOI21_X1  g725(.A(G301), .B1(new_n1136), .B2(new_n1141), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1148), .A2(KEYINPUT54), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1149), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1073), .B1(new_n1058), .B2(new_n1056), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1144), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1086), .B1(new_n1132), .B2(new_n1156), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1138), .A2(new_n1019), .A3(new_n1139), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n983), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1159), .A2(G1996), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT111), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT111), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(new_n1159), .B2(G1996), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n799), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n799), .A2(G1996), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n833), .B(G2067), .Z(new_n1166));
  AOI21_X1  g741(.A(new_n1159), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n699), .B(new_n702), .Z(new_n1169));
  OR2_X1    g744(.A1(new_n1159), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  OR2_X1    g746(.A1(G290), .A2(G1986), .ZN(new_n1172));
  NAND2_X1  g747(.A1(G290), .A2(G1986), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1159), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1157), .A2(new_n1175), .ZN(new_n1176));
  NOR4_X1   g751(.A1(new_n1164), .A2(new_n702), .A3(new_n699), .A4(new_n1167), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n833), .A2(G2067), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n983), .B(new_n1158), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1172), .A2(new_n1159), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n1180), .B(KEYINPUT48), .Z(new_n1181));
  NAND3_X1  g756(.A1(new_n1168), .A2(new_n1181), .A3(new_n1170), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1159), .B1(new_n800), .B2(new_n1166), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT46), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1161), .A2(KEYINPUT46), .A3(new_n1163), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1183), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT47), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1179), .B(new_n1182), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1176), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g769(.A1(G227), .A2(new_n460), .ZN(new_n1196));
  OAI21_X1  g770(.A(new_n659), .B1(new_n1196), .B2(KEYINPUT127), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n1197), .B1(new_n903), .B2(new_n905), .ZN(new_n1198));
  AOI21_X1  g772(.A(G229), .B1(KEYINPUT127), .B2(new_n1196), .ZN(new_n1199));
  AND4_X1   g773(.A1(new_n964), .A2(new_n1198), .A3(new_n965), .A4(new_n1199), .ZN(G308));
  NAND4_X1  g774(.A1(new_n1198), .A2(new_n964), .A3(new_n965), .A4(new_n1199), .ZN(G225));
endmodule


