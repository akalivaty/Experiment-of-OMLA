//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n543, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n462), .A2(new_n464), .A3(G137), .A4(new_n460), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n461), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n462), .A2(new_n464), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n460), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n460), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n475), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT69), .ZN(G162));
  NAND4_X1  g056(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n460), .ZN(new_n482));
  XNOR2_X1  g057(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(KEYINPUT3), .B(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n485), .A2(G138), .A3(new_n460), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT70), .B1(new_n460), .B2(G114), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n490), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n462), .A2(new_n464), .A3(G126), .A4(G2105), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n488), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  XNOR2_X1  g074(.A(KEYINPUT5), .B(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT72), .A2(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT72), .A3(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n502), .A2(new_n504), .A3(G543), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n509), .A2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  NAND2_X1  g089(.A1(new_n502), .A2(new_n504), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n521), .A2(G89), .ZN(new_n522));
  AND2_X1   g097(.A1(G63), .A2(G651), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT7), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n500), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n526), .B1(new_n524), .B2(new_n525), .ZN(new_n527));
  INV_X1    g102(.A(new_n508), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  OR3_X1    g104(.A1(new_n522), .A2(new_n527), .A3(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  AND2_X1   g106(.A1(new_n521), .A2(G90), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n528), .A2(G52), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n511), .ZN(new_n535));
  NOR3_X1   g110(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(G171));
  AND2_X1   g111(.A1(new_n521), .A2(G81), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n528), .A2(G43), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n511), .ZN(new_n540));
  NOR3_X1   g115(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G188));
  AOI22_X1  g122(.A1(new_n500), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n511), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT73), .B(KEYINPUT9), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n528), .A2(G53), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OAI211_X1 g128(.A(KEYINPUT73), .B(new_n552), .C1(new_n508), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n521), .A2(G91), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n549), .A2(new_n551), .A3(new_n554), .A4(new_n555), .ZN(G299));
  INV_X1    g131(.A(G171), .ZN(G301));
  NAND4_X1  g132(.A1(new_n502), .A2(new_n504), .A3(G49), .A4(G543), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n500), .A2(G87), .A3(new_n502), .A4(new_n504), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n558), .A2(new_n559), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT75), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n558), .A2(new_n559), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n560), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(G288));
  NAND4_X1  g145(.A1(new_n502), .A2(new_n504), .A3(G48), .A4(G543), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n500), .A2(G86), .A3(new_n502), .A4(new_n504), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n500), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n511), .ZN(G305));
  NAND4_X1  g149(.A1(new_n500), .A2(G85), .A3(new_n502), .A4(new_n504), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n502), .A2(new_n504), .A3(G47), .A4(G543), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n511), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT76), .ZN(new_n579));
  NAND2_X1  g154(.A1(G72), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G60), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n520), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n583), .A2(new_n584), .A3(new_n575), .A4(new_n576), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n579), .A2(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n521), .A2(new_n588), .A3(G92), .ZN(new_n589));
  INV_X1    g164(.A(G92), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT77), .B1(new_n505), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n591), .A3(KEYINPUT10), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n520), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(G651), .A2(new_n595), .B1(new_n528), .B2(G54), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(KEYINPUT10), .B1(new_n589), .B2(new_n591), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n587), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n587), .B1(new_n599), .B2(G868), .ZN(G321));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(G299), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G168), .B2(new_n602), .ZN(G280));
  XOR2_X1   g179(.A(G280), .B(KEYINPUT78), .Z(G297));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  INV_X1    g182(.A(new_n541), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(new_n602), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n599), .A2(new_n606), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n609), .B1(new_n611), .B2(new_n602), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n476), .A2(G135), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G111), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n617), .A2(new_n618), .B1(new_n620), .B2(G2105), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n474), .A2(G123), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2096), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n485), .A2(new_n469), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  AND2_X1   g203(.A1(KEYINPUT80), .A2(G2100), .ZN(new_n629));
  NOR2_X1   g204(.A1(KEYINPUT80), .A2(G2100), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n624), .B(new_n631), .C1(new_n629), .C2(new_n628), .ZN(G156));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2435), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT16), .B(G1341), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n641), .B(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(G14), .B1(new_n638), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n638), .B2(new_n644), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT83), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n650), .A2(new_n651), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n653), .B1(new_n658), .B2(new_n652), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(G227));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT85), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(new_n663), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n668), .A2(new_n666), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n667), .B1(KEYINPUT20), .B2(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(KEYINPUT20), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n664), .A2(new_n668), .A3(new_n666), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(G1991), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G1996), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n678), .ZN(new_n682));
  AND3_X1   g257(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n681), .B1(new_n679), .B2(new_n682), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(G229));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G5), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G171), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G1961), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n469), .A2(G103), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT25), .ZN(new_n691));
  AOI22_X1  g266(.A1(new_n485), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n692), .A2(new_n460), .ZN(new_n693));
  AOI211_X1 g268(.A(new_n691), .B(new_n693), .C1(G139), .C2(new_n476), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n695), .B2(G33), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n697), .A2(G2072), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(G2072), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n689), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n623), .A2(G29), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT96), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G1961), .B2(new_n688), .ZN(new_n704));
  AND2_X1   g279(.A1(KEYINPUT24), .A2(G34), .ZN(new_n705));
  NOR2_X1   g280(.A1(KEYINPUT24), .A2(G34), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n695), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT93), .ZN(new_n708));
  INV_X1    g283(.A(G160), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n695), .ZN(new_n710));
  INV_X1    g285(.A(G2084), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT30), .B(G28), .ZN(new_n714));
  OR2_X1    g289(.A1(KEYINPUT31), .A2(G11), .ZN(new_n715));
  NAND2_X1  g290(.A1(KEYINPUT31), .A2(G11), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n714), .A2(new_n695), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n712), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n700), .A2(new_n704), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n686), .A2(G4), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n599), .B2(new_n686), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT91), .B(G1348), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G164), .A2(new_n695), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G27), .B2(new_n695), .ZN(new_n725));
  INV_X1    g300(.A(G2078), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n541), .A2(G16), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G16), .B2(G19), .ZN(new_n729));
  INV_X1    g304(.A(G1341), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n725), .A2(new_n726), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(new_n730), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n727), .A2(new_n731), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(G168), .A2(G16), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G16), .B2(G21), .ZN(new_n736));
  INV_X1    g311(.A(G1966), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n474), .A2(G128), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n476), .A2(G140), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n460), .A2(G116), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n740), .B(new_n741), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G29), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n695), .A2(G26), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT92), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2067), .ZN(new_n750));
  NOR4_X1   g325(.A1(new_n734), .A2(new_n738), .A3(new_n739), .A4(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n719), .A2(new_n723), .A3(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G2090), .ZN(new_n753));
  NOR2_X1   g328(.A1(G162), .A2(new_n695), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n695), .A2(G35), .ZN(new_n755));
  OAI21_X1  g330(.A(KEYINPUT97), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(KEYINPUT97), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n758), .A2(new_n759), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n753), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n758), .A2(new_n759), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n764), .A2(G2090), .A3(new_n760), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  AOI22_X1  g341(.A1(G129), .A2(new_n474), .B1(new_n476), .B2(G141), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT26), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n770), .A2(new_n771), .B1(G105), .B2(new_n469), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT94), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT95), .ZN(new_n776));
  OR2_X1    g351(.A1(G29), .A2(G32), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT27), .B(G1996), .Z(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT23), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n686), .A2(G20), .ZN(new_n783));
  AOI211_X1 g358(.A(new_n782), .B(new_n783), .C1(G299), .C2(G16), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n782), .B2(new_n783), .ZN(new_n785));
  INV_X1    g360(.A(G1956), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n776), .A2(new_n779), .A3(new_n777), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n781), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n752), .A2(new_n766), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT36), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n476), .A2(G131), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n474), .A2(G119), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT88), .ZN(new_n794));
  OR3_X1    g369(.A1(new_n794), .A2(G95), .A3(G2105), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(G95), .B2(G2105), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n460), .A2(G107), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n795), .A2(new_n796), .A3(G2104), .A4(new_n797), .ZN(new_n798));
  AND3_X1   g373(.A1(new_n792), .A2(new_n793), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G29), .ZN(new_n800));
  OR2_X1    g375(.A1(G25), .A2(G29), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n800), .A2(KEYINPUT89), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(KEYINPUT89), .B1(new_n800), .B2(new_n801), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT35), .B(G1991), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NOR3_X1   g381(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n800), .A2(new_n801), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT89), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n805), .B1(new_n810), .B2(new_n802), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  MUX2_X1   g387(.A(G24), .B(G290), .S(G16), .Z(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(G1986), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(G1986), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n686), .A2(G22), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G166), .B2(new_n686), .ZN(new_n819));
  INV_X1    g394(.A(G1971), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n686), .A2(G6), .ZN(new_n822));
  INV_X1    g397(.A(new_n572), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n517), .A2(new_n519), .A3(G61), .ZN(new_n824));
  NAND2_X1  g399(.A1(G73), .A2(G543), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n511), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n571), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n823), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n822), .B1(new_n828), .B2(new_n686), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT32), .B(G1981), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(G16), .A2(G23), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n563), .A2(new_n564), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(G16), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT33), .B(G1976), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n821), .A2(new_n831), .A3(new_n836), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n817), .B(KEYINPUT90), .C1(KEYINPUT34), .C2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT90), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n837), .A2(KEYINPUT34), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(new_n816), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n837), .A2(KEYINPUT34), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n791), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n843), .ZN(new_n845));
  AOI211_X1 g420(.A(KEYINPUT36), .B(new_n845), .C1(new_n838), .C2(new_n841), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n790), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n790), .B(KEYINPUT99), .C1(new_n844), .C2(new_n846), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(G311));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n790), .B(KEYINPUT100), .C1(new_n844), .C2(new_n846), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(G150));
  NAND2_X1  g430(.A1(new_n521), .A2(G93), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n528), .A2(G55), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n856), .B(new_n857), .C1(new_n511), .C2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G860), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n608), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n541), .A2(new_n859), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT39), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n599), .A2(G559), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT38), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n862), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n868), .A2(new_n870), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n864), .B1(new_n872), .B2(new_n873), .ZN(G145));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n694), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n627), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n495), .A2(new_n878), .A3(new_n496), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n878), .B1(new_n495), .B2(new_n496), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n488), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n877), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n799), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n774), .B(new_n623), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(G162), .B(KEYINPUT102), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(G160), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n888), .A2(G160), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n888), .A2(G160), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n889), .A3(new_n886), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n474), .A2(G130), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n476), .A2(G142), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n460), .A2(G118), .ZN(new_n897));
  OAI21_X1  g472(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n895), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n744), .B(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n892), .A2(new_n894), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n901), .B1(new_n892), .B2(new_n894), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n885), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n883), .B(new_n799), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n892), .A2(new_n894), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n900), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n908), .A3(new_n902), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g487(.A1(new_n833), .A2(new_n579), .A3(new_n585), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n833), .B1(new_n579), .B2(new_n585), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n828), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n833), .ZN(new_n917));
  NAND2_X1  g492(.A1(G290), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n918), .A2(G305), .A3(new_n913), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n920));
  XNOR2_X1  g495(.A(G303), .B(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n916), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(new_n916), .B2(new_n919), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT42), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT106), .ZN(new_n925));
  INV_X1    g500(.A(new_n921), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n914), .A2(new_n915), .A3(new_n828), .ZN(new_n927));
  AOI21_X1  g502(.A(G305), .B1(new_n918), .B2(new_n913), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n916), .A2(new_n919), .A3(new_n921), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT42), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n922), .A2(new_n923), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT42), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(KEYINPUT107), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n931), .B2(KEYINPUT42), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n610), .B1(new_n865), .B2(new_n866), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n865), .A2(new_n610), .A3(new_n866), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n599), .B(G299), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT41), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n599), .A2(G299), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n599), .A2(G299), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT41), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n942), .B(new_n943), .C1(new_n946), .C2(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n942), .A2(new_n943), .ZN(new_n951));
  INV_X1    g526(.A(new_n944), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n934), .A2(new_n940), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n934), .B2(new_n940), .ZN(new_n955));
  OAI21_X1  g530(.A(G868), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n861), .A2(G868), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(G295));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n956), .A2(new_n960), .A3(new_n958), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(new_n956), .B2(new_n958), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(G331));
  NAND2_X1  g538(.A1(new_n952), .A2(KEYINPUT41), .ZN(new_n964));
  INV_X1    g539(.A(new_n949), .ZN(new_n965));
  XNOR2_X1  g540(.A(G286), .B(G171), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(new_n865), .A3(new_n866), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n867), .A2(new_n966), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n964), .A2(new_n965), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n944), .A3(new_n969), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n935), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n969), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(new_n949), .B2(new_n946), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(new_n931), .A3(new_n971), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n976), .A3(new_n910), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n970), .A2(new_n972), .ZN(new_n980));
  AOI21_X1  g555(.A(G37), .B1(new_n980), .B2(new_n931), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n973), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g558(.A(KEYINPUT109), .B(new_n935), .C1(new_n970), .C2(new_n972), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n979), .B1(new_n985), .B2(new_n978), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT44), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n981), .A2(new_n983), .A3(new_n978), .A4(new_n984), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n987), .A2(new_n992), .ZN(G397));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  INV_X1    g569(.A(G40), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n467), .A2(new_n471), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n881), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n566), .A2(G1976), .A3(new_n568), .A4(new_n560), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n997), .A2(G8), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1976), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT52), .B1(G288), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n495), .A2(new_n496), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT103), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n495), .A2(new_n878), .A3(new_n496), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1384), .B1(new_n1007), .B2(new_n488), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1003), .B1(new_n1008), .B2(new_n996), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n1010));
  INV_X1    g585(.A(G1981), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n828), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  AND3_X1   g588(.A1(G305), .A2(new_n1013), .A3(G1981), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(G305), .B2(G1981), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT49), .B1(new_n828), .B2(new_n1011), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT115), .B1(G305), .B2(G1981), .ZN(new_n1018));
  NAND3_X1  g593(.A1(G305), .A2(new_n1013), .A3(G1981), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1009), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n997), .A2(G8), .ZN(new_n1022));
  INV_X1    g597(.A(new_n998), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT52), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1002), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1002), .A2(new_n1021), .A3(new_n1024), .A4(KEYINPUT118), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n881), .A2(KEYINPUT45), .A3(new_n994), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n488), .B2(new_n497), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n996), .B1(new_n1031), .B2(KEYINPUT45), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n820), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n498), .A2(new_n994), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT50), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n881), .A2(new_n1036), .A3(new_n994), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1035), .A2(new_n1037), .A3(new_n753), .A4(new_n996), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1003), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(G303), .A2(G8), .ZN(new_n1040));
  XOR2_X1   g615(.A(new_n1040), .B(KEYINPUT55), .Z(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1040), .B(KEYINPUT55), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n881), .A2(new_n994), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT50), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G160), .A2(G40), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n753), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1033), .A2(new_n1048), .A3(KEYINPUT117), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT117), .B1(new_n1033), .B2(new_n1048), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1043), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1029), .A2(new_n1042), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1035), .A2(new_n1037), .A3(new_n996), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(G2084), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT45), .B1(new_n881), .B2(new_n994), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT119), .B1(new_n1056), .B2(new_n1046), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(new_n996), .C1(new_n1008), .C2(KEYINPUT45), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1031), .A2(KEYINPUT45), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1055), .B1(new_n1061), .B2(new_n737), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1003), .B1(new_n1062), .B2(G168), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(G286), .A2(G8), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT51), .B(new_n1066), .C1(new_n1062), .C2(new_n1003), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT45), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1046), .B1(new_n1034), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n881), .A2(KEYINPUT45), .A3(new_n994), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n726), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n1072));
  INV_X1    g647(.A(G1961), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1071), .A2(new_n1072), .B1(new_n1054), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n726), .A2(KEYINPUT53), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1074), .B1(new_n1061), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(KEYINPUT62), .A3(G171), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1065), .A2(new_n1067), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1065), .A2(new_n1067), .A3(new_n1078), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT62), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1076), .A2(new_n1081), .A3(G171), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  XOR2_X1   g658(.A(G171), .B(KEYINPUT54), .Z(new_n1084));
  INV_X1    g659(.A(new_n1056), .ZN(new_n1085));
  INV_X1    g660(.A(new_n471), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT123), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(KEYINPUT123), .ZN(new_n1088));
  NOR4_X1   g663(.A1(new_n1088), .A2(new_n995), .A3(new_n467), .A4(new_n1075), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1085), .A2(new_n1070), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1084), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1092), .B(new_n1074), .C1(new_n1091), .C2(new_n1090), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1076), .A2(new_n1084), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G1348), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n881), .A2(new_n1036), .A3(new_n994), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n996), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n997), .ZN(new_n1100));
  INV_X1    g675(.A(G2067), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n599), .ZN(new_n1103));
  AND4_X1   g678(.A1(KEYINPUT60), .A2(new_n1099), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1103), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1054), .A2(new_n1096), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT60), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1104), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1996), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1069), .A2(new_n1111), .A3(new_n1070), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT58), .B(G1341), .Z(new_n1113));
  NAND2_X1  g688(.A1(new_n997), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n608), .A2(KEYINPUT122), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT59), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1115), .A2(new_n1119), .A3(new_n1116), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT56), .B(G2072), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1069), .A2(new_n1070), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(G1956), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1126));
  XNOR2_X1  g701(.A(G299), .B(KEYINPUT57), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n1129));
  XNOR2_X1  g704(.A(G299), .B(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1047), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1036), .B1(new_n881), .B2(new_n994), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n786), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1130), .B1(new_n1133), .B2(new_n1124), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1122), .B1(new_n1128), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1127), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1130), .A3(new_n1124), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(KEYINPUT61), .A3(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1110), .A2(new_n1121), .A3(new_n1135), .A4(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1108), .A2(new_n1103), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1137), .B1(new_n1140), .B2(new_n1134), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1095), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1053), .B(new_n1079), .C1(new_n1083), .C2(new_n1142), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1062), .A2(new_n1003), .A3(G286), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1144), .A2(new_n1029), .A3(new_n1042), .A4(new_n1052), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1025), .A2(KEYINPUT116), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1149), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1038), .ZN(new_n1151));
  AOI21_X1  g726(.A(G1971), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1152));
  OAI21_X1  g727(.A(G8), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n1043), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT116), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1002), .A2(new_n1021), .A3(new_n1024), .A4(new_n1155), .ZN(new_n1156));
  AND4_X1   g731(.A1(new_n1148), .A2(new_n1150), .A3(new_n1154), .A4(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1144), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1147), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1148), .A2(new_n1041), .A3(new_n1039), .A4(new_n1156), .ZN(new_n1161));
  AND4_X1   g736(.A1(new_n1000), .A2(new_n1021), .A3(new_n565), .A4(new_n569), .ZN(new_n1162));
  NOR2_X1   g737(.A1(G305), .A2(G1981), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1009), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1159), .A2(new_n1160), .A3(new_n1166), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1145), .A2(new_n1146), .B1(new_n1157), .B2(new_n1144), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT121), .B1(new_n1168), .B2(new_n1165), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1143), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1056), .A2(new_n996), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT112), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1171), .B(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n744), .B(new_n1101), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT113), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1171), .B(KEYINPUT112), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1178), .A2(new_n1111), .A3(new_n774), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1171), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1111), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT111), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1179), .B1(new_n774), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n884), .A2(new_n805), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n799), .A2(new_n806), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1173), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OR2_X1    g761(.A1(G290), .A2(G1986), .ZN(new_n1187));
  NAND2_X1  g762(.A1(G290), .A2(G1986), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1187), .A2(KEYINPUT110), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT110), .ZN(new_n1190));
  NAND3_X1  g765(.A1(G290), .A2(new_n1190), .A3(G1986), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1189), .A2(new_n1180), .A3(new_n1191), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1177), .A2(new_n1183), .A3(new_n1186), .A4(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT114), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1170), .A2(new_n1194), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1177), .A2(new_n1183), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1186), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1187), .A2(new_n1171), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT125), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT48), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT47), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1178), .B1(new_n774), .B2(new_n1174), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1202), .B1(KEYINPUT46), .B2(new_n1182), .ZN(new_n1203));
  OR2_X1    g778(.A1(new_n1182), .A2(KEYINPUT46), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1201), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AND3_X1   g780(.A1(new_n1203), .A2(new_n1204), .A3(new_n1201), .ZN(new_n1206));
  OAI22_X1  g781(.A1(new_n1197), .A2(new_n1200), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1196), .A2(new_n1184), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n744), .A2(G2067), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1178), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1207), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1195), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g787(.A(new_n458), .ZN(new_n1214));
  NOR2_X1   g788(.A1(G227), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g789(.A1(new_n647), .A2(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g790(.A(new_n1216), .B(KEYINPUT126), .ZN(new_n1217));
  OAI21_X1  g791(.A(KEYINPUT127), .B1(G229), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n1219));
  XNOR2_X1  g793(.A(new_n1216), .B(new_n1219), .ZN(new_n1220));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n1221));
  OAI211_X1 g795(.A(new_n1220), .B(new_n1221), .C1(new_n683), .C2(new_n684), .ZN(new_n1222));
  NAND4_X1  g796(.A1(new_n990), .A2(new_n1218), .A3(new_n1222), .A4(new_n911), .ZN(G225));
  INV_X1    g797(.A(G225), .ZN(G308));
endmodule


