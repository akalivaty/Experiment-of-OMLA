

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591;

  XOR2_X1 U324 ( .A(G22GAT), .B(G155GAT), .Z(n436) );
  XNOR2_X1 U325 ( .A(n415), .B(KEYINPUT9), .ZN(n417) );
  INV_X1 U326 ( .A(n489), .ZN(n447) );
  XNOR2_X1 U327 ( .A(n380), .B(n379), .ZN(n385) );
  XNOR2_X1 U328 ( .A(n308), .B(n307), .ZN(n539) );
  AND2_X1 U329 ( .A1(G228GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U330 ( .A(n329), .B(KEYINPUT33), .ZN(n330) );
  XNOR2_X1 U331 ( .A(KEYINPUT114), .B(KEYINPUT47), .ZN(n461) );
  XNOR2_X1 U332 ( .A(n426), .B(n330), .ZN(n336) );
  XNOR2_X1 U333 ( .A(n417), .B(n416), .ZN(n421) );
  XNOR2_X1 U334 ( .A(n462), .B(n461), .ZN(n469) );
  NAND2_X1 U335 ( .A1(n587), .A2(n563), .ZN(n446) );
  XNOR2_X1 U336 ( .A(n378), .B(n292), .ZN(n379) );
  XNOR2_X1 U337 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U338 ( .A(n405), .B(KEYINPUT94), .ZN(n574) );
  XOR2_X1 U339 ( .A(KEYINPUT36), .B(n566), .Z(n587) );
  XNOR2_X1 U340 ( .A(n344), .B(n343), .ZN(n350) );
  INV_X1 U341 ( .A(n574), .ZN(n555) );
  XNOR2_X1 U342 ( .A(n429), .B(n428), .ZN(n566) );
  XOR2_X1 U343 ( .A(n474), .B(KEYINPUT28), .Z(n537) );
  XNOR2_X1 U344 ( .A(KEYINPUT38), .B(n451), .ZN(n509) );
  XNOR2_X1 U345 ( .A(n484), .B(KEYINPUT58), .ZN(n485) );
  XNOR2_X1 U346 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U347 ( .A(n486), .B(n485), .ZN(G1351GAT) );
  XNOR2_X1 U348 ( .A(n455), .B(n454), .ZN(G1330GAT) );
  XOR2_X1 U349 ( .A(G71GAT), .B(G176GAT), .Z(n294) );
  XNOR2_X1 U350 ( .A(G190GAT), .B(G183GAT), .ZN(n293) );
  XNOR2_X1 U351 ( .A(n294), .B(n293), .ZN(n308) );
  XOR2_X1 U352 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n296) );
  NAND2_X1 U353 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U354 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U355 ( .A(n297), .B(KEYINPUT20), .Z(n303) );
  XOR2_X1 U356 ( .A(G120GAT), .B(KEYINPUT0), .Z(n299) );
  XNOR2_X1 U357 ( .A(G113GAT), .B(G134GAT), .ZN(n298) );
  XNOR2_X1 U358 ( .A(n299), .B(n298), .ZN(n362) );
  XOR2_X1 U359 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n301) );
  XNOR2_X1 U360 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n300) );
  XNOR2_X1 U361 ( .A(n301), .B(n300), .ZN(n392) );
  XNOR2_X1 U362 ( .A(n362), .B(n392), .ZN(n302) );
  XNOR2_X1 U363 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U364 ( .A(G15GAT), .B(G127GAT), .Z(n437) );
  XOR2_X1 U365 ( .A(n304), .B(n437), .Z(n306) );
  XNOR2_X1 U366 ( .A(G43GAT), .B(G99GAT), .ZN(n305) );
  XNOR2_X1 U367 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U368 ( .A(G29GAT), .B(G43GAT), .Z(n310) );
  XNOR2_X1 U369 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n309) );
  XNOR2_X1 U370 ( .A(n310), .B(n309), .ZN(n427) );
  XOR2_X1 U371 ( .A(G1GAT), .B(KEYINPUT68), .Z(n443) );
  XOR2_X1 U372 ( .A(n427), .B(n443), .Z(n312) );
  NAND2_X1 U373 ( .A1(G229GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U374 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U375 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n314) );
  XNOR2_X1 U376 ( .A(G15GAT), .B(KEYINPUT67), .ZN(n313) );
  XNOR2_X1 U377 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U378 ( .A(n316), .B(n315), .Z(n324) );
  XOR2_X1 U379 ( .A(G141GAT), .B(G113GAT), .Z(n318) );
  XNOR2_X1 U380 ( .A(G50GAT), .B(G36GAT), .ZN(n317) );
  XNOR2_X1 U381 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U382 ( .A(G22GAT), .B(G197GAT), .Z(n320) );
  XNOR2_X1 U383 ( .A(G169GAT), .B(G8GAT), .ZN(n319) );
  XNOR2_X1 U384 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U386 ( .A(n324), .B(n323), .Z(n577) );
  INV_X1 U387 ( .A(n577), .ZN(n569) );
  INV_X1 U388 ( .A(G85GAT), .ZN(n328) );
  XOR2_X1 U389 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n326) );
  XNOR2_X1 U390 ( .A(G99GAT), .B(G92GAT), .ZN(n325) );
  XNOR2_X1 U391 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U392 ( .A(n328), .B(n327), .ZN(n426) );
  XOR2_X1 U393 ( .A(KEYINPUT31), .B(KEYINPUT76), .Z(n329) );
  INV_X1 U394 ( .A(n336), .ZN(n335) );
  XOR2_X1 U395 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n332) );
  XNOR2_X1 U396 ( .A(G148GAT), .B(G106GAT), .ZN(n331) );
  XNOR2_X1 U397 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U398 ( .A(G204GAT), .B(n333), .Z(n378) );
  INV_X1 U399 ( .A(n378), .ZN(n334) );
  NAND2_X1 U400 ( .A1(n335), .A2(n334), .ZN(n338) );
  NAND2_X1 U401 ( .A1(n336), .A2(n378), .ZN(n337) );
  NAND2_X1 U402 ( .A1(n338), .A2(n337), .ZN(n344) );
  XOR2_X1 U403 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n340) );
  XNOR2_X1 U404 ( .A(G120GAT), .B(KEYINPUT77), .ZN(n339) );
  XOR2_X1 U405 ( .A(n340), .B(n339), .Z(n342) );
  AND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U407 ( .A(G176GAT), .B(G64GAT), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n345), .B(KEYINPUT75), .ZN(n391) );
  XOR2_X1 U409 ( .A(G78GAT), .B(KEYINPUT69), .Z(n347) );
  XNOR2_X1 U410 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U412 ( .A(G71GAT), .B(n348), .Z(n442) );
  XOR2_X1 U413 ( .A(n391), .B(n442), .Z(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n582) );
  NOR2_X1 U415 ( .A1(n569), .A2(n582), .ZN(n491) );
  XOR2_X1 U416 ( .A(KEYINPUT88), .B(KEYINPUT1), .Z(n352) );
  XNOR2_X1 U417 ( .A(G1GAT), .B(KEYINPUT87), .ZN(n351) );
  XNOR2_X1 U418 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U419 ( .A(KEYINPUT4), .B(KEYINPUT89), .Z(n354) );
  XNOR2_X1 U420 ( .A(KEYINPUT90), .B(KEYINPUT5), .ZN(n353) );
  XNOR2_X1 U421 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U423 ( .A(G57GAT), .B(G148GAT), .Z(n358) );
  XNOR2_X1 U424 ( .A(G127GAT), .B(G162GAT), .ZN(n357) );
  XNOR2_X1 U425 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U427 ( .A(n361), .B(G155GAT), .Z(n364) );
  XNOR2_X1 U428 ( .A(n362), .B(KEYINPUT6), .ZN(n363) );
  XNOR2_X1 U429 ( .A(n364), .B(n363), .ZN(n371) );
  XOR2_X1 U430 ( .A(KEYINPUT85), .B(KEYINPUT3), .Z(n366) );
  XNOR2_X1 U431 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n365) );
  XNOR2_X1 U432 ( .A(n366), .B(n365), .ZN(n383) );
  XOR2_X1 U433 ( .A(G85GAT), .B(n383), .Z(n368) );
  NAND2_X1 U434 ( .A1(G225GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U435 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U436 ( .A(G29GAT), .B(n369), .Z(n370) );
  XOR2_X1 U437 ( .A(n371), .B(n370), .Z(n410) );
  XOR2_X1 U438 ( .A(KEYINPUT24), .B(KEYINPUT86), .Z(n373) );
  XNOR2_X1 U439 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U441 ( .A(n436), .B(G78GAT), .Z(n375) );
  XOR2_X1 U442 ( .A(G197GAT), .B(KEYINPUT21), .Z(n395) );
  XNOR2_X1 U443 ( .A(G211GAT), .B(n395), .ZN(n374) );
  XNOR2_X1 U444 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U445 ( .A(n377), .B(n376), .Z(n380) );
  XOR2_X1 U446 ( .A(KEYINPUT78), .B(G218GAT), .Z(n382) );
  XNOR2_X1 U447 ( .A(G50GAT), .B(G162GAT), .ZN(n381) );
  XNOR2_X1 U448 ( .A(n382), .B(n381), .ZN(n424) );
  XNOR2_X1 U449 ( .A(n383), .B(n424), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n385), .B(n384), .ZN(n474) );
  XNOR2_X1 U451 ( .A(G36GAT), .B(G190GAT), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n386), .B(KEYINPUT80), .ZN(n416) );
  XNOR2_X1 U453 ( .A(G8GAT), .B(G183GAT), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n387), .B(G211GAT), .ZN(n433) );
  XNOR2_X1 U455 ( .A(n416), .B(n433), .ZN(n400) );
  XOR2_X1 U456 ( .A(G204GAT), .B(KEYINPUT91), .Z(n389) );
  NAND2_X1 U457 ( .A1(G226GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U458 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U459 ( .A(n390), .B(KEYINPUT92), .Z(n394) );
  XNOR2_X1 U460 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n394), .B(n393), .ZN(n396) );
  XOR2_X1 U462 ( .A(n396), .B(n395), .Z(n398) );
  XNOR2_X1 U463 ( .A(G218GAT), .B(G92GAT), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U465 ( .A(n400), .B(n399), .ZN(n526) );
  NOR2_X1 U466 ( .A1(n526), .A2(n539), .ZN(n401) );
  NOR2_X1 U467 ( .A1(n474), .A2(n401), .ZN(n402) );
  XOR2_X1 U468 ( .A(KEYINPUT25), .B(n402), .Z(n407) );
  XOR2_X1 U469 ( .A(n526), .B(KEYINPUT93), .Z(n403) );
  XNOR2_X1 U470 ( .A(KEYINPUT27), .B(n403), .ZN(n411) );
  NAND2_X1 U471 ( .A1(n539), .A2(n474), .ZN(n404) );
  XNOR2_X1 U472 ( .A(n404), .B(KEYINPUT26), .ZN(n405) );
  NOR2_X1 U473 ( .A1(n411), .A2(n574), .ZN(n406) );
  NOR2_X1 U474 ( .A1(n407), .A2(n406), .ZN(n408) );
  NOR2_X1 U475 ( .A1(n410), .A2(n408), .ZN(n409) );
  XNOR2_X1 U476 ( .A(n409), .B(KEYINPUT95), .ZN(n414) );
  AND2_X1 U477 ( .A1(n539), .A2(n537), .ZN(n412) );
  INV_X1 U478 ( .A(n410), .ZN(n523) );
  NOR2_X1 U479 ( .A1(n523), .A2(n411), .ZN(n534) );
  NAND2_X1 U480 ( .A1(n412), .A2(n534), .ZN(n413) );
  NAND2_X1 U481 ( .A1(n414), .A2(n413), .ZN(n489) );
  XOR2_X1 U482 ( .A(KEYINPUT65), .B(G106GAT), .Z(n415) );
  XOR2_X1 U483 ( .A(KEYINPUT79), .B(KEYINPUT10), .Z(n419) );
  NAND2_X1 U484 ( .A1(G232GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U485 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U486 ( .A(n421), .B(n420), .Z(n423) );
  XNOR2_X1 U487 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n422) );
  XNOR2_X1 U488 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U489 ( .A(n425), .B(n424), .Z(n429) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U491 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n435) );
  XOR2_X1 U492 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n431) );
  XNOR2_X1 U493 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n441) );
  XOR2_X1 U497 ( .A(n437), .B(n436), .Z(n439) );
  NAND2_X1 U498 ( .A1(G231GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U500 ( .A(n441), .B(n440), .Z(n445) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U502 ( .A(n445), .B(n444), .Z(n563) );
  INV_X1 U503 ( .A(n563), .ZN(n585) );
  NOR2_X1 U504 ( .A1(n447), .A2(n446), .ZN(n449) );
  XNOR2_X1 U505 ( .A(KEYINPUT103), .B(KEYINPUT37), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n522) );
  NAND2_X1 U507 ( .A1(n491), .A2(n522), .ZN(n450) );
  XNOR2_X1 U508 ( .A(n450), .B(KEYINPUT104), .ZN(n451) );
  NOR2_X1 U509 ( .A1(n539), .A2(n509), .ZN(n455) );
  XNOR2_X1 U510 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n453) );
  INV_X1 U511 ( .A(G43GAT), .ZN(n452) );
  XOR2_X1 U512 ( .A(KEYINPUT123), .B(KEYINPUT55), .Z(n476) );
  XNOR2_X1 U513 ( .A(n582), .B(KEYINPUT41), .ZN(n479) );
  NOR2_X1 U514 ( .A1(n479), .A2(n569), .ZN(n457) );
  INV_X1 U515 ( .A(KEYINPUT46), .ZN(n456) );
  XNOR2_X1 U516 ( .A(n457), .B(n456), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n563), .B(KEYINPUT113), .ZN(n572) );
  INV_X1 U518 ( .A(n566), .ZN(n458) );
  NOR2_X1 U519 ( .A1(n572), .A2(n458), .ZN(n459) );
  NAND2_X1 U520 ( .A1(n460), .A2(n459), .ZN(n462) );
  NAND2_X1 U521 ( .A1(n585), .A2(n587), .ZN(n464) );
  XOR2_X1 U522 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n463) );
  XNOR2_X1 U523 ( .A(n464), .B(n463), .ZN(n466) );
  INV_X1 U524 ( .A(n582), .ZN(n465) );
  NAND2_X1 U525 ( .A1(n466), .A2(n465), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n577), .A2(n467), .ZN(n468) );
  NOR2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n470), .B(KEYINPUT48), .ZN(n536) );
  NOR2_X1 U529 ( .A1(n536), .A2(n526), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT54), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n472), .A2(n523), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n473), .B(KEYINPUT64), .ZN(n575) );
  NOR2_X1 U533 ( .A1(n575), .A2(n474), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n476), .B(n475), .ZN(n477) );
  NOR2_X1 U535 ( .A1(n539), .A2(n477), .ZN(n478) );
  INV_X1 U536 ( .A(n478), .ZN(n571) );
  XNOR2_X1 U537 ( .A(n479), .B(KEYINPUT108), .ZN(n542) );
  NOR2_X1 U538 ( .A1(n571), .A2(n542), .ZN(n483) );
  XNOR2_X1 U539 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n481) );
  XNOR2_X1 U540 ( .A(KEYINPUT57), .B(KEYINPUT124), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(G1349GAT) );
  NOR2_X1 U543 ( .A1(n566), .A2(n571), .ZN(n486) );
  INV_X1 U544 ( .A(G190GAT), .ZN(n484) );
  NAND2_X1 U545 ( .A1(n566), .A2(n585), .ZN(n487) );
  XOR2_X1 U546 ( .A(KEYINPUT16), .B(n487), .Z(n488) );
  NAND2_X1 U547 ( .A1(n489), .A2(n488), .ZN(n490) );
  XOR2_X1 U548 ( .A(KEYINPUT96), .B(n490), .Z(n512) );
  NAND2_X1 U549 ( .A1(n491), .A2(n512), .ZN(n501) );
  NOR2_X1 U550 ( .A1(n523), .A2(n501), .ZN(n493) );
  XNOR2_X1 U551 ( .A(KEYINPUT97), .B(KEYINPUT34), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U553 ( .A(G1GAT), .B(n494), .ZN(G1324GAT) );
  NOR2_X1 U554 ( .A1(n526), .A2(n501), .ZN(n495) );
  XOR2_X1 U555 ( .A(G8GAT), .B(n495), .Z(G1325GAT) );
  NOR2_X1 U556 ( .A1(n539), .A2(n501), .ZN(n500) );
  XOR2_X1 U557 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n497) );
  XNOR2_X1 U558 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U560 ( .A(KEYINPUT98), .B(n498), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1326GAT) );
  NOR2_X1 U562 ( .A1(n537), .A2(n501), .ZN(n503) );
  XNOR2_X1 U563 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U565 ( .A(G22GAT), .B(n504), .ZN(G1327GAT) );
  NOR2_X1 U566 ( .A1(n523), .A2(n509), .ZN(n506) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(G1328GAT) );
  NOR2_X1 U569 ( .A1(n526), .A2(n509), .ZN(n508) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n508), .B(n507), .ZN(G1329GAT) );
  NOR2_X1 U572 ( .A1(n537), .A2(n509), .ZN(n511) );
  XNOR2_X1 U573 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(G1331GAT) );
  NOR2_X1 U575 ( .A1(n577), .A2(n542), .ZN(n521) );
  NAND2_X1 U576 ( .A1(n521), .A2(n512), .ZN(n518) );
  NOR2_X1 U577 ( .A1(n523), .A2(n518), .ZN(n513) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n513), .Z(n514) );
  XNOR2_X1 U579 ( .A(KEYINPUT42), .B(n514), .ZN(G1332GAT) );
  NOR2_X1 U580 ( .A1(n526), .A2(n518), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(G1333GAT) );
  NOR2_X1 U583 ( .A1(n539), .A2(n518), .ZN(n517) );
  XOR2_X1 U584 ( .A(G71GAT), .B(n517), .Z(G1334GAT) );
  NOR2_X1 U585 ( .A1(n537), .A2(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NAND2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n530) );
  NOR2_X1 U589 ( .A1(n523), .A2(n530), .ZN(n524) );
  XOR2_X1 U590 ( .A(G85GAT), .B(n524), .Z(n525) );
  XNOR2_X1 U591 ( .A(KEYINPUT110), .B(n525), .ZN(G1336GAT) );
  NOR2_X1 U592 ( .A1(n526), .A2(n530), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(G1337GAT) );
  NOR2_X1 U595 ( .A1(n539), .A2(n530), .ZN(n529) );
  XOR2_X1 U596 ( .A(G99GAT), .B(n529), .Z(G1338GAT) );
  NOR2_X1 U597 ( .A1(n537), .A2(n530), .ZN(n532) );
  XNOR2_X1 U598 ( .A(KEYINPUT112), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U600 ( .A(G106GAT), .B(n533), .Z(G1339GAT) );
  XOR2_X1 U601 ( .A(G113GAT), .B(KEYINPUT115), .Z(n541) );
  INV_X1 U602 ( .A(n534), .ZN(n535) );
  NOR2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n554) );
  NAND2_X1 U604 ( .A1(n537), .A2(n554), .ZN(n538) );
  NOR2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n546) );
  NAND2_X1 U606 ( .A1(n546), .A2(n577), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1340GAT) );
  INV_X1 U608 ( .A(n546), .ZN(n550) );
  NOR2_X1 U609 ( .A1(n542), .A2(n550), .ZN(n544) );
  XNOR2_X1 U610 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(G120GAT), .B(n545), .ZN(G1341GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n548) );
  NAND2_X1 U614 ( .A1(n546), .A2(n572), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  NOR2_X1 U617 ( .A1(n566), .A2(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G134GAT), .B(n553), .ZN(G1343GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n565) );
  NOR2_X1 U622 ( .A1(n569), .A2(n565), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  NOR2_X1 U625 ( .A1(n479), .A2(n565), .ZN(n562) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n559) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n558) );
  XNOR2_X1 U628 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U629 ( .A(KEYINPUT120), .B(n560), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(G1345GAT) );
  NOR2_X1 U631 ( .A1(n563), .A2(n565), .ZN(n564) );
  XOR2_X1 U632 ( .A(G155GAT), .B(n564), .Z(G1346GAT) );
  NOR2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT122), .B(n567), .Z(n568) );
  XNOR2_X1 U635 ( .A(G162GAT), .B(n568), .ZN(G1347GAT) );
  NOR2_X1 U636 ( .A1(n569), .A2(n571), .ZN(n570) );
  XOR2_X1 U637 ( .A(G169GAT), .B(n570), .Z(G1348GAT) );
  NAND2_X1 U638 ( .A1(n478), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(KEYINPUT125), .B(n576), .Z(n588) );
  NAND2_X1 U642 ( .A1(n577), .A2(n588), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  NAND2_X1 U648 ( .A1(n588), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n588), .A2(n585), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n590) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

