

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777;

  NOR2_X1 U374 ( .A1(n420), .A2(n422), .ZN(n425) );
  XNOR2_X1 U375 ( .A(n388), .B(n497), .ZN(n448) );
  NOR2_X1 U376 ( .A1(n635), .A2(n634), .ZN(n647) );
  NOR2_X1 U377 ( .A1(n622), .A2(n650), .ZN(n726) );
  NOR2_X1 U378 ( .A1(n631), .A2(n638), .ZN(n430) );
  NOR2_X1 U379 ( .A1(n617), .A2(n628), .ZN(n618) );
  NOR2_X1 U380 ( .A1(G900), .A2(n614), .ZN(n616) );
  XNOR2_X1 U381 ( .A(n546), .B(n462), .ZN(n461) );
  XNOR2_X1 U382 ( .A(n556), .B(KEYINPUT95), .ZN(n613) );
  XNOR2_X1 U383 ( .A(n522), .B(n501), .ZN(n763) );
  XNOR2_X1 U384 ( .A(n502), .B(G125), .ZN(n522) );
  XNOR2_X2 U385 ( .A(n661), .B(KEYINPUT86), .ZN(n493) );
  XNOR2_X2 U386 ( .A(n474), .B(n473), .ZN(n376) );
  NAND2_X1 U387 ( .A1(n353), .A2(n363), .ZN(n392) );
  INV_X1 U388 ( .A(n448), .ZN(n353) );
  XOR2_X2 U389 ( .A(G116), .B(G107), .Z(n586) );
  XNOR2_X2 U390 ( .A(n354), .B(n515), .ZN(n550) );
  XNOR2_X2 U391 ( .A(n413), .B(n412), .ZN(n354) );
  NOR2_X1 U392 ( .A1(n742), .A2(G902), .ZN(n540) );
  NAND2_X1 U393 ( .A1(n621), .A2(n489), .ZN(n396) );
  XOR2_X1 U394 ( .A(n428), .B(KEYINPUT74), .Z(n355) );
  AND2_X2 U395 ( .A1(n440), .A2(n435), .ZN(n434) );
  XNOR2_X2 U396 ( .A(n648), .B(KEYINPUT40), .ZN(n776) );
  XNOR2_X1 U397 ( .A(n544), .B(KEYINPUT97), .ZN(n761) );
  AND2_X2 U398 ( .A1(n407), .A2(n355), .ZN(n665) );
  INV_X2 U399 ( .A(n506), .ZN(n508) );
  XNOR2_X2 U400 ( .A(G101), .B(KEYINPUT3), .ZN(n506) );
  XNOR2_X1 U401 ( .A(KEYINPUT38), .B(n646), .ZN(n688) );
  INV_X1 U402 ( .A(n678), .ZN(n631) );
  INV_X2 U403 ( .A(G953), .ZN(n764) );
  INV_X1 U404 ( .A(G146), .ZN(n502) );
  AND2_X1 U405 ( .A1(n647), .A2(n688), .ZN(n479) );
  XNOR2_X1 U406 ( .A(n527), .B(n526), .ZN(n751) );
  XNOR2_X1 U407 ( .A(n763), .B(n525), .ZN(n526) );
  XNOR2_X1 U408 ( .A(n534), .B(n533), .ZN(n544) );
  XNOR2_X1 U409 ( .A(n374), .B(n373), .ZN(n774) );
  XNOR2_X1 U410 ( .A(n479), .B(n478), .ZN(n654) );
  NAND2_X1 U411 ( .A1(n647), .A2(n463), .ZN(n391) );
  NOR2_X1 U412 ( .A1(n381), .A2(n378), .ZN(n630) );
  NOR2_X1 U413 ( .A1(n691), .A2(n693), .ZN(n649) );
  NAND2_X1 U414 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U415 ( .A1(n380), .A2(n379), .ZN(n378) );
  INV_X1 U416 ( .A(n396), .ZN(n395) );
  NAND2_X1 U417 ( .A1(n619), .A2(KEYINPUT110), .ZN(n382) );
  XNOR2_X1 U418 ( .A(KEYINPUT99), .B(n674), .ZN(n598) );
  XNOR2_X1 U419 ( .A(n385), .B(n384), .ZN(n527) );
  XNOR2_X1 U420 ( .A(n588), .B(KEYINPUT4), .ZN(n534) );
  XNOR2_X1 U421 ( .A(n570), .B(n509), .ZN(n462) );
  XNOR2_X1 U422 ( .A(n387), .B(G110), .ZN(n520) );
  XNOR2_X1 U423 ( .A(n519), .B(n521), .ZN(n384) );
  BUF_X1 U424 ( .A(n777), .Z(n356) );
  XNOR2_X1 U425 ( .A(n652), .B(n651), .ZN(n777) );
  NAND2_X1 U426 ( .A1(n563), .A2(n562), .ZN(n357) );
  NAND2_X1 U427 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U428 ( .A(n439), .B(KEYINPUT22), .ZN(n416) );
  XNOR2_X1 U429 ( .A(n621), .B(KEYINPUT1), .ZN(n680) );
  XNOR2_X1 U430 ( .A(n391), .B(n390), .ZN(n389) );
  INV_X1 U431 ( .A(KEYINPUT83), .ZN(n390) );
  AND2_X1 U432 ( .A1(n486), .A2(KEYINPUT44), .ZN(n442) );
  INV_X1 U433 ( .A(KEYINPUT48), .ZN(n473) );
  XNOR2_X1 U434 ( .A(n549), .B(n548), .ZN(n678) );
  XNOR2_X1 U435 ( .A(n593), .B(n457), .ZN(n603) );
  XNOR2_X1 U436 ( .A(G478), .B(KEYINPUT105), .ZN(n457) );
  INV_X1 U437 ( .A(n735), .ZN(n423) );
  INV_X1 U438 ( .A(KEYINPUT81), .ZN(n497) );
  NAND2_X1 U439 ( .A1(n498), .A2(n389), .ZN(n388) );
  OR2_X1 U440 ( .A1(G902), .A2(G237), .ZN(n552) );
  AND2_X1 U441 ( .A1(n774), .A2(n485), .ZN(n484) );
  XOR2_X1 U442 ( .A(KEYINPUT69), .B(KEYINPUT73), .Z(n536) );
  INV_X1 U443 ( .A(n534), .ZN(n412) );
  XOR2_X1 U444 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n511) );
  AND2_X1 U445 ( .A1(n680), .A2(n681), .ZN(n402) );
  XNOR2_X1 U446 ( .A(n582), .B(n581), .ZN(n602) );
  XNOR2_X1 U447 ( .A(KEYINPUT10), .B(G140), .ZN(n501) );
  XNOR2_X1 U448 ( .A(n761), .B(n465), .ZN(n742) );
  XNOR2_X1 U449 ( .A(n467), .B(n466), .ZN(n465) );
  XNOR2_X1 U450 ( .A(n361), .B(n535), .ZN(n466) );
  XNOR2_X1 U451 ( .A(n538), .B(n468), .ZN(n467) );
  INV_X1 U452 ( .A(n671), .ZN(n426) );
  XNOR2_X1 U453 ( .A(n403), .B(KEYINPUT34), .ZN(n375) );
  NOR2_X1 U454 ( .A1(n706), .A2(n404), .ZN(n403) );
  NAND2_X1 U455 ( .A1(n398), .A2(n595), .ZN(n439) );
  NOR2_X1 U456 ( .A1(n598), .A2(n691), .ZN(n595) );
  XNOR2_X1 U457 ( .A(n564), .B(n399), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n678), .B(KEYINPUT6), .ZN(n639) );
  XNOR2_X1 U459 ( .A(n591), .B(n592), .ZN(n748) );
  XNOR2_X1 U460 ( .A(n503), .B(n590), .ZN(n591) );
  XOR2_X1 U461 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n585) );
  NAND2_X1 U462 ( .A1(n376), .A2(n365), .ZN(n661) );
  NOR2_X1 U463 ( .A1(n423), .A2(n424), .ZN(n421) );
  AND2_X1 U464 ( .A1(n637), .A2(KEYINPUT72), .ZN(n424) );
  AND2_X1 U465 ( .A1(n448), .A2(KEYINPUT72), .ZN(n422) );
  INV_X1 U466 ( .A(KEYINPUT46), .ZN(n476) );
  NAND2_X1 U467 ( .A1(n441), .A2(n432), .ZN(n431) );
  NOR2_X1 U468 ( .A1(n433), .A2(n486), .ZN(n432) );
  NOR2_X1 U469 ( .A1(G953), .A2(G237), .ZN(n572) );
  NAND2_X1 U470 ( .A1(G237), .A2(G234), .ZN(n554) );
  XOR2_X1 U471 ( .A(KEYINPUT14), .B(KEYINPUT93), .Z(n555) );
  NAND2_X1 U472 ( .A1(n362), .A2(n395), .ZN(n383) );
  XNOR2_X1 U473 ( .A(G902), .B(KEYINPUT15), .ZN(n663) );
  XNOR2_X1 U474 ( .A(G134), .B(G137), .ZN(n532) );
  XOR2_X1 U475 ( .A(KEYINPUT5), .B(G119), .Z(n542) );
  XNOR2_X1 U476 ( .A(G116), .B(G146), .ZN(n541) );
  XOR2_X1 U477 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n574) );
  XNOR2_X1 U478 ( .A(G143), .B(G113), .ZN(n567) );
  XOR2_X1 U479 ( .A(G131), .B(KEYINPUT12), .Z(n568) );
  XNOR2_X1 U480 ( .A(G110), .B(G101), .ZN(n537) );
  INV_X1 U481 ( .A(n536), .ZN(n468) );
  XNOR2_X1 U482 ( .A(n360), .B(n366), .ZN(n706) );
  INV_X1 U483 ( .A(n639), .ZN(n400) );
  XNOR2_X1 U484 ( .A(KEYINPUT92), .B(n553), .ZN(n689) );
  INV_X1 U485 ( .A(KEYINPUT0), .ZN(n399) );
  INV_X1 U486 ( .A(KEYINPUT16), .ZN(n509) );
  INV_X1 U487 ( .A(G119), .ZN(n387) );
  XNOR2_X1 U488 ( .A(KEYINPUT23), .B(KEYINPUT84), .ZN(n521) );
  XNOR2_X1 U489 ( .A(G128), .B(G137), .ZN(n519) );
  XNOR2_X1 U490 ( .A(n520), .B(n386), .ZN(n385) );
  XNOR2_X1 U491 ( .A(KEYINPUT24), .B(KEYINPUT98), .ZN(n386) );
  XNOR2_X1 U492 ( .A(KEYINPUT71), .B(KEYINPUT39), .ZN(n478) );
  INV_X1 U493 ( .A(n767), .ZN(n427) );
  NOR2_X1 U494 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U495 ( .A(n470), .B(KEYINPUT35), .ZN(n373) );
  NAND2_X1 U496 ( .A1(n375), .A2(n599), .ZN(n374) );
  XNOR2_X1 U497 ( .A(n415), .B(n414), .ZN(n733) );
  XNOR2_X1 U498 ( .A(KEYINPUT31), .B(KEYINPUT100), .ZN(n414) );
  NOR2_X1 U499 ( .A1(n636), .A2(n464), .ZN(n463) );
  NAND2_X1 U500 ( .A1(n481), .A2(n631), .ZN(n418) );
  NOR2_X1 U501 ( .A1(n680), .A2(n675), .ZN(n481) );
  NAND2_X1 U502 ( .A1(n600), .A2(n639), .ZN(n438) );
  INV_X1 U503 ( .A(n751), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n747), .B(n748), .ZN(n446) );
  INV_X1 U505 ( .A(KEYINPUT60), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n740), .B(n451), .ZN(n445) );
  XNOR2_X1 U507 ( .A(n743), .B(n741), .ZN(n451) );
  XNOR2_X1 U508 ( .A(n411), .B(G110), .ZN(G12) );
  XOR2_X1 U509 ( .A(n586), .B(n520), .Z(n358) );
  AND2_X1 U510 ( .A1(n402), .A2(n401), .ZN(n359) );
  AND2_X1 U511 ( .A1(n400), .A2(n402), .ZN(n360) );
  INV_X1 U512 ( .A(n619), .ZN(n488) );
  XOR2_X1 U513 ( .A(G104), .B(G140), .Z(n361) );
  AND2_X1 U514 ( .A1(n488), .A2(n394), .ZN(n362) );
  NOR2_X1 U515 ( .A1(n637), .A2(KEYINPUT72), .ZN(n363) );
  AND2_X1 U516 ( .A1(n428), .A2(n426), .ZN(n364) );
  INV_X1 U517 ( .A(n631), .ZN(n401) );
  AND2_X1 U518 ( .A1(n660), .A2(KEYINPUT2), .ZN(n365) );
  XNOR2_X1 U519 ( .A(KEYINPUT33), .B(KEYINPUT70), .ZN(n366) );
  XOR2_X1 U520 ( .A(n714), .B(KEYINPUT62), .Z(n367) );
  XNOR2_X1 U521 ( .A(n744), .B(KEYINPUT59), .ZN(n368) );
  XNOR2_X1 U522 ( .A(n550), .B(n518), .ZN(n369) );
  INV_X1 U523 ( .A(KEYINPUT88), .ZN(n486) );
  INV_X1 U524 ( .A(KEYINPUT44), .ZN(n485) );
  XNOR2_X1 U525 ( .A(KEYINPUT63), .B(KEYINPUT112), .ZN(n370) );
  XOR2_X1 U526 ( .A(n713), .B(KEYINPUT53), .Z(n371) );
  XOR2_X1 U527 ( .A(n669), .B(KEYINPUT87), .Z(n372) );
  XNOR2_X2 U528 ( .A(n540), .B(n539), .ZN(n621) );
  NAND2_X1 U529 ( .A1(n376), .A2(n660), .ZN(n428) );
  NAND2_X2 U530 ( .A1(n377), .A2(n664), .ZN(n667) );
  NAND2_X1 U531 ( .A1(n377), .A2(n670), .ZN(n673) );
  NAND2_X2 U532 ( .A1(n490), .A2(n492), .ZN(n377) );
  INV_X1 U533 ( .A(n628), .ZN(n379) );
  NAND2_X1 U534 ( .A1(n396), .A2(KEYINPUT110), .ZN(n380) );
  INV_X1 U535 ( .A(n391), .ZN(n724) );
  NAND2_X1 U536 ( .A1(n392), .A2(n421), .ZN(n420) );
  NAND2_X1 U537 ( .A1(n395), .A2(n488), .ZN(n627) );
  INV_X1 U538 ( .A(KEYINPUT110), .ZN(n394) );
  NOR2_X2 U539 ( .A1(n410), .A2(n397), .ZN(n480) );
  INV_X1 U540 ( .A(n411), .ZN(n397) );
  XNOR2_X1 U541 ( .A(n405), .B(KEYINPUT32), .ZN(n410) );
  XNOR2_X1 U542 ( .A(n357), .B(KEYINPUT0), .ZN(n404) );
  XNOR2_X2 U543 ( .A(n551), .B(n504), .ZN(n658) );
  NOR2_X1 U544 ( .A1(n416), .A2(n419), .ZN(n405) );
  INV_X1 U545 ( .A(n646), .ZN(n406) );
  XNOR2_X1 U546 ( .A(n482), .B(KEYINPUT45), .ZN(n407) );
  XNOR2_X1 U547 ( .A(n482), .B(KEYINPUT45), .ZN(n408) );
  XNOR2_X1 U548 ( .A(n482), .B(KEYINPUT45), .ZN(n417) );
  NAND2_X1 U549 ( .A1(n746), .A2(G472), .ZN(n496) );
  NAND2_X1 U550 ( .A1(n495), .A2(n458), .ZN(n494) );
  XNOR2_X1 U551 ( .A(n496), .B(n367), .ZN(n495) );
  INV_X1 U552 ( .A(n752), .ZN(n458) );
  NAND2_X1 U553 ( .A1(n409), .A2(n774), .ZN(n469) );
  XNOR2_X2 U554 ( .A(n480), .B(KEYINPUT90), .ZN(n409) );
  XNOR2_X1 U555 ( .A(n409), .B(n611), .ZN(n612) );
  XNOR2_X1 U556 ( .A(n410), .B(n775), .ZN(G21) );
  OR2_X1 U557 ( .A1(n416), .A2(n418), .ZN(n411) );
  XNOR2_X1 U558 ( .A(n413), .B(KEYINPUT73), .ZN(n757) );
  XNOR2_X2 U559 ( .A(n461), .B(n358), .ZN(n413) );
  NAND2_X1 U560 ( .A1(n606), .A2(n359), .ZN(n415) );
  INV_X1 U561 ( .A(n404), .ZN(n606) );
  OR2_X1 U562 ( .A1(n416), .A2(n438), .ZN(n601) );
  NAND2_X1 U563 ( .A1(n417), .A2(n471), .ZN(n491) );
  NAND2_X1 U564 ( .A1(n472), .A2(n408), .ZN(n492) );
  OR2_X1 U565 ( .A1(n407), .A2(n671), .ZN(n670) );
  NAND2_X1 U566 ( .A1(n407), .A2(n764), .ZN(n756) );
  NAND2_X1 U567 ( .A1(n597), .A2(n639), .ZN(n419) );
  NAND2_X2 U568 ( .A1(n444), .A2(n483), .ZN(n482) );
  NAND2_X1 U569 ( .A1(n475), .A2(n425), .ZN(n474) );
  XNOR2_X1 U570 ( .A(n428), .B(n427), .ZN(n765) );
  NAND2_X1 U571 ( .A1(n429), .A2(n621), .ZN(n650) );
  XNOR2_X1 U572 ( .A(n430), .B(KEYINPUT28), .ZN(n429) );
  NAND2_X1 U573 ( .A1(n434), .A2(n431), .ZN(n444) );
  INV_X1 U574 ( .A(n610), .ZN(n433) );
  NAND2_X1 U575 ( .A1(n437), .A2(n436), .ZN(n435) );
  NAND2_X1 U576 ( .A1(n610), .A2(n443), .ZN(n436) );
  NAND2_X1 U577 ( .A1(n433), .A2(KEYINPUT88), .ZN(n437) );
  NAND2_X1 U578 ( .A1(n469), .A2(n442), .ZN(n440) );
  INV_X1 U579 ( .A(n469), .ZN(n441) );
  NAND2_X1 U580 ( .A1(KEYINPUT88), .A2(n485), .ZN(n443) );
  NOR2_X1 U581 ( .A1(n445), .A2(n752), .ZN(G54) );
  XNOR2_X1 U582 ( .A(n477), .B(n476), .ZN(n475) );
  NOR2_X1 U583 ( .A1(n446), .A2(n752), .ZN(G63) );
  NOR2_X2 U584 ( .A1(KEYINPUT2), .A2(n665), .ZN(n666) );
  XNOR2_X1 U585 ( .A(n447), .B(n371), .ZN(G75) );
  NAND2_X1 U586 ( .A1(n456), .A2(n764), .ZN(n447) );
  AND2_X1 U587 ( .A1(n449), .A2(n458), .ZN(G66) );
  XNOR2_X1 U588 ( .A(n750), .B(n450), .ZN(n449) );
  BUF_X2 U589 ( .A(n746), .Z(n749) );
  XNOR2_X1 U590 ( .A(n452), .B(n372), .ZN(G51) );
  NAND2_X1 U591 ( .A1(n460), .A2(n458), .ZN(n452) );
  XNOR2_X1 U592 ( .A(n454), .B(n453), .ZN(G60) );
  NAND2_X1 U593 ( .A1(n459), .A2(n458), .ZN(n454) );
  XNOR2_X2 U594 ( .A(G113), .B(KEYINPUT68), .ZN(n507) );
  XNOR2_X2 U595 ( .A(n508), .B(n507), .ZN(n546) );
  XNOR2_X1 U596 ( .A(n712), .B(KEYINPUT122), .ZN(n456) );
  INV_X1 U597 ( .A(n624), .ZN(n623) );
  XNOR2_X1 U598 ( .A(n692), .B(KEYINPUT82), .ZN(n624) );
  XNOR2_X1 U599 ( .A(n745), .B(n368), .ZN(n459) );
  XNOR2_X1 U600 ( .A(n668), .B(n369), .ZN(n460) );
  INV_X1 U601 ( .A(n493), .ZN(n471) );
  INV_X1 U602 ( .A(n406), .ZN(n464) );
  INV_X1 U603 ( .A(KEYINPUT78), .ZN(n470) );
  NOR2_X1 U604 ( .A1(n493), .A2(n662), .ZN(n472) );
  NAND2_X1 U605 ( .A1(n776), .A2(n777), .ZN(n477) );
  NAND2_X1 U606 ( .A1(n654), .A2(n729), .ZN(n648) );
  NAND2_X1 U607 ( .A1(n612), .A2(n484), .ZN(n483) );
  INV_X1 U608 ( .A(n563), .ZN(n622) );
  XNOR2_X2 U609 ( .A(n487), .B(KEYINPUT19), .ZN(n563) );
  NAND2_X1 U610 ( .A1(n658), .A2(n689), .ZN(n487) );
  XNOR2_X2 U611 ( .A(n531), .B(n530), .ZN(n619) );
  NOR2_X1 U612 ( .A1(n619), .A2(n598), .ZN(n681) );
  INV_X1 U613 ( .A(n598), .ZN(n489) );
  NAND2_X1 U614 ( .A1(n491), .A2(n662), .ZN(n490) );
  XNOR2_X2 U615 ( .A(G143), .B(G128), .ZN(n588) );
  XNOR2_X1 U616 ( .A(n494), .B(n370), .ZN(G57) );
  NAND2_X1 U617 ( .A1(n499), .A2(KEYINPUT47), .ZN(n498) );
  NAND2_X1 U618 ( .A1(n726), .A2(n692), .ZN(n499) );
  NOR2_X1 U619 ( .A1(n714), .A2(G902), .ZN(n548) );
  XNOR2_X1 U620 ( .A(n544), .B(n500), .ZN(n714) );
  XNOR2_X1 U621 ( .A(n547), .B(n543), .ZN(n500) );
  XNOR2_X1 U622 ( .A(n630), .B(n629), .ZN(n635) );
  NOR2_X2 U623 ( .A1(G902), .A2(n751), .ZN(n531) );
  XOR2_X1 U624 ( .A(n586), .B(n587), .Z(n503) );
  AND2_X1 U625 ( .A1(G210), .A2(n552), .ZN(n504) );
  AND2_X1 U626 ( .A1(G227), .A2(n764), .ZN(n505) );
  INV_X1 U627 ( .A(KEYINPUT89), .ZN(n611) );
  XNOR2_X1 U628 ( .A(n532), .B(G131), .ZN(n533) );
  INV_X1 U629 ( .A(KEYINPUT76), .ZN(n629) );
  INV_X1 U630 ( .A(G475), .ZN(n579) );
  XNOR2_X1 U631 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U632 ( .A(n505), .B(n537), .ZN(n538) );
  XNOR2_X1 U633 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U634 ( .A(n580), .B(n579), .ZN(n581) );
  NOR2_X1 U635 ( .A1(G952), .A2(n764), .ZN(n752) );
  XNOR2_X2 U636 ( .A(G122), .B(G104), .ZN(n570) );
  NAND2_X1 U637 ( .A1(G224), .A2(n764), .ZN(n510) );
  XNOR2_X1 U638 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U639 ( .A(n512), .B(KEYINPUT77), .Z(n514) );
  XNOR2_X1 U640 ( .A(n522), .B(n536), .ZN(n513) );
  XOR2_X1 U641 ( .A(KEYINPUT91), .B(KEYINPUT79), .Z(n517) );
  XNOR2_X1 U642 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n516) );
  XNOR2_X1 U643 ( .A(n517), .B(n516), .ZN(n518) );
  NAND2_X1 U644 ( .A1(n764), .A2(G234), .ZN(n524) );
  XNOR2_X1 U645 ( .A(KEYINPUT65), .B(KEYINPUT8), .ZN(n523) );
  XNOR2_X1 U646 ( .A(n524), .B(n523), .ZN(n583) );
  NAND2_X1 U647 ( .A1(G221), .A2(n583), .ZN(n525) );
  NAND2_X1 U648 ( .A1(G234), .A2(n663), .ZN(n528) );
  XNOR2_X1 U649 ( .A(KEYINPUT20), .B(n528), .ZN(n565) );
  NAND2_X1 U650 ( .A1(n565), .A2(G217), .ZN(n529) );
  XOR2_X1 U651 ( .A(KEYINPUT25), .B(n529), .Z(n530) );
  INV_X1 U652 ( .A(n619), .ZN(n675) );
  XNOR2_X1 U653 ( .A(G107), .B(G146), .ZN(n535) );
  XNOR2_X1 U654 ( .A(KEYINPUT67), .B(G469), .ZN(n539) );
  INV_X1 U655 ( .A(n680), .ZN(n600) );
  INV_X1 U656 ( .A(G472), .ZN(n549) );
  XNOR2_X1 U657 ( .A(n542), .B(n541), .ZN(n543) );
  NAND2_X1 U658 ( .A1(G210), .A2(n572), .ZN(n545) );
  NAND2_X1 U659 ( .A1(n550), .A2(n663), .ZN(n551) );
  NAND2_X1 U660 ( .A1(G214), .A2(n552), .ZN(n553) );
  XNOR2_X1 U661 ( .A(n555), .B(n554), .ZN(n558) );
  NAND2_X1 U662 ( .A1(n558), .A2(G902), .ZN(n556) );
  NOR2_X1 U663 ( .A1(G898), .A2(n764), .ZN(n758) );
  NAND2_X1 U664 ( .A1(n613), .A2(n758), .ZN(n557) );
  XNOR2_X1 U665 ( .A(KEYINPUT96), .B(n557), .ZN(n561) );
  NAND2_X1 U666 ( .A1(n558), .A2(G952), .ZN(n704) );
  NOR2_X1 U667 ( .A1(G953), .A2(n704), .ZN(n559) );
  XNOR2_X1 U668 ( .A(KEYINPUT94), .B(n559), .ZN(n615) );
  INV_X1 U669 ( .A(n615), .ZN(n560) );
  NAND2_X1 U670 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U671 ( .A1(n565), .A2(G221), .ZN(n566) );
  XNOR2_X1 U672 ( .A(n566), .B(KEYINPUT21), .ZN(n617) );
  INV_X1 U673 ( .A(n617), .ZN(n674) );
  XNOR2_X1 U674 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U675 ( .A(n763), .B(n569), .ZN(n578) );
  INV_X1 U676 ( .A(n570), .ZN(n571) );
  XNOR2_X1 U677 ( .A(n571), .B(KEYINPUT11), .ZN(n576) );
  NAND2_X1 U678 ( .A1(n572), .A2(G214), .ZN(n573) );
  XNOR2_X1 U679 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U680 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U681 ( .A(n578), .B(n577), .ZN(n744) );
  NOR2_X1 U682 ( .A1(G902), .A2(n744), .ZN(n582) );
  XNOR2_X1 U683 ( .A(KEYINPUT13), .B(KEYINPUT103), .ZN(n580) );
  NAND2_X1 U684 ( .A1(G217), .A2(n583), .ZN(n584) );
  XNOR2_X1 U685 ( .A(n585), .B(n584), .ZN(n592) );
  XNOR2_X1 U686 ( .A(KEYINPUT104), .B(G122), .ZN(n587) );
  INV_X1 U687 ( .A(n588), .ZN(n589) );
  XNOR2_X1 U688 ( .A(G134), .B(n589), .ZN(n590) );
  NOR2_X1 U689 ( .A1(G902), .A2(n748), .ZN(n593) );
  NOR2_X1 U690 ( .A1(n602), .A2(n603), .ZN(n594) );
  XNOR2_X1 U691 ( .A(n594), .B(KEYINPUT107), .ZN(n691) );
  NOR2_X1 U692 ( .A1(n600), .A2(n675), .ZN(n596) );
  XNOR2_X1 U693 ( .A(KEYINPUT108), .B(n596), .ZN(n597) );
  NAND2_X1 U694 ( .A1(n603), .A2(n602), .ZN(n636) );
  INV_X1 U695 ( .A(n636), .ZN(n599) );
  NOR2_X1 U696 ( .A1(n619), .A2(n601), .ZN(n715) );
  INV_X1 U697 ( .A(n602), .ZN(n604) );
  NAND2_X1 U698 ( .A1(n603), .A2(n604), .ZN(n653) );
  NOR2_X2 U699 ( .A1(n604), .A2(n603), .ZN(n729) );
  INV_X1 U700 ( .A(n729), .ZN(n642) );
  NAND2_X1 U701 ( .A1(n653), .A2(n642), .ZN(n605) );
  XNOR2_X1 U702 ( .A(n605), .B(KEYINPUT106), .ZN(n692) );
  NAND2_X1 U703 ( .A1(n606), .A2(n631), .ZN(n607) );
  NOR2_X1 U704 ( .A1(n627), .A2(n607), .ZN(n717) );
  NOR2_X1 U705 ( .A1(n733), .A2(n717), .ZN(n608) );
  NOR2_X1 U706 ( .A1(n623), .A2(n608), .ZN(n609) );
  NOR2_X1 U707 ( .A1(n715), .A2(n609), .ZN(n610) );
  NAND2_X1 U708 ( .A1(G953), .A2(n613), .ZN(n614) );
  NOR2_X1 U709 ( .A1(n616), .A2(n615), .ZN(n628) );
  XNOR2_X1 U710 ( .A(KEYINPUT66), .B(n618), .ZN(n620) );
  NAND2_X1 U711 ( .A1(n620), .A2(n619), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n726), .A2(n624), .ZN(n626) );
  XNOR2_X1 U713 ( .A(KEYINPUT47), .B(KEYINPUT64), .ZN(n625) );
  NOR2_X1 U714 ( .A1(n626), .A2(n625), .ZN(n637) );
  INV_X1 U715 ( .A(n689), .ZN(n632) );
  NOR2_X1 U716 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U717 ( .A(KEYINPUT30), .B(n633), .Z(n634) );
  INV_X1 U718 ( .A(n658), .ZN(n646) );
  NOR2_X1 U719 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U720 ( .A(n640), .B(KEYINPUT109), .ZN(n641) );
  NOR2_X1 U721 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n689), .A2(n643), .ZN(n655) );
  NOR2_X1 U723 ( .A1(n646), .A2(n655), .ZN(n644) );
  XNOR2_X1 U724 ( .A(n644), .B(KEYINPUT36), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n645), .A2(n680), .ZN(n735) );
  NAND2_X1 U726 ( .A1(n689), .A2(n688), .ZN(n693) );
  XNOR2_X1 U727 ( .A(KEYINPUT41), .B(n649), .ZN(n705) );
  NOR2_X1 U728 ( .A1(n705), .A2(n650), .ZN(n652) );
  XNOR2_X1 U729 ( .A(KEYINPUT42), .B(KEYINPUT111), .ZN(n651) );
  INV_X1 U730 ( .A(n653), .ZN(n732) );
  NAND2_X1 U731 ( .A1(n732), .A2(n654), .ZN(n738) );
  NOR2_X1 U732 ( .A1(n680), .A2(n655), .ZN(n656) );
  XNOR2_X1 U733 ( .A(n656), .B(KEYINPUT43), .ZN(n657) );
  NOR2_X1 U734 ( .A1(n406), .A2(n657), .ZN(n739) );
  INV_X1 U735 ( .A(n739), .ZN(n659) );
  AND2_X1 U736 ( .A1(n738), .A2(n659), .ZN(n660) );
  INV_X1 U737 ( .A(KEYINPUT75), .ZN(n662) );
  INV_X1 U738 ( .A(n663), .ZN(n664) );
  NOR2_X4 U739 ( .A1(n667), .A2(n666), .ZN(n746) );
  NAND2_X1 U740 ( .A1(n746), .A2(G210), .ZN(n668) );
  INV_X1 U741 ( .A(KEYINPUT56), .ZN(n669) );
  XNOR2_X1 U742 ( .A(KEYINPUT2), .B(KEYINPUT80), .ZN(n671) );
  XOR2_X1 U743 ( .A(KEYINPUT85), .B(n364), .Z(n672) );
  NOR2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n711) );
  NOR2_X1 U745 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U746 ( .A(KEYINPUT49), .B(n676), .Z(n677) );
  NOR2_X1 U747 ( .A1(n401), .A2(n677), .ZN(n679) );
  XOR2_X1 U748 ( .A(KEYINPUT118), .B(n679), .Z(n684) );
  NOR2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U750 ( .A(KEYINPUT50), .B(n682), .ZN(n683) );
  NOR2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U752 ( .A1(n359), .A2(n685), .ZN(n686) );
  XOR2_X1 U753 ( .A(KEYINPUT51), .B(n686), .Z(n687) );
  NOR2_X1 U754 ( .A1(n705), .A2(n687), .ZN(n700) );
  NOR2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n697) );
  INV_X1 U757 ( .A(n692), .ZN(n694) );
  NOR2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U759 ( .A(KEYINPUT119), .B(n695), .Z(n696) );
  NOR2_X1 U760 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U761 ( .A1(n706), .A2(n698), .ZN(n699) );
  NOR2_X1 U762 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U763 ( .A(n701), .B(KEYINPUT52), .ZN(n702) );
  XNOR2_X1 U764 ( .A(KEYINPUT120), .B(n702), .ZN(n703) );
  NOR2_X1 U765 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U766 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U767 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U768 ( .A(n709), .B(KEYINPUT121), .ZN(n710) );
  INV_X1 U769 ( .A(KEYINPUT123), .ZN(n713) );
  XOR2_X1 U770 ( .A(G101), .B(n715), .Z(G3) );
  NAND2_X1 U771 ( .A1(n717), .A2(n729), .ZN(n716) );
  XNOR2_X1 U772 ( .A(n716), .B(G104), .ZN(G6) );
  XOR2_X1 U773 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n719) );
  NAND2_X1 U774 ( .A1(n717), .A2(n732), .ZN(n718) );
  XNOR2_X1 U775 ( .A(n719), .B(n718), .ZN(n721) );
  XOR2_X1 U776 ( .A(G107), .B(KEYINPUT27), .Z(n720) );
  XNOR2_X1 U777 ( .A(n721), .B(n720), .ZN(G9) );
  XOR2_X1 U778 ( .A(G128), .B(KEYINPUT29), .Z(n723) );
  NAND2_X1 U779 ( .A1(n726), .A2(n732), .ZN(n722) );
  XNOR2_X1 U780 ( .A(n723), .B(n722), .ZN(G30) );
  XOR2_X1 U781 ( .A(n724), .B(G143), .Z(n725) );
  XNOR2_X1 U782 ( .A(KEYINPUT114), .B(n725), .ZN(G45) );
  XOR2_X1 U783 ( .A(G146), .B(KEYINPUT115), .Z(n728) );
  NAND2_X1 U784 ( .A1(n726), .A2(n729), .ZN(n727) );
  XNOR2_X1 U785 ( .A(n728), .B(n727), .ZN(G48) );
  NAND2_X1 U786 ( .A1(n733), .A2(n729), .ZN(n730) );
  XNOR2_X1 U787 ( .A(n730), .B(KEYINPUT116), .ZN(n731) );
  XNOR2_X1 U788 ( .A(G113), .B(n731), .ZN(G15) );
  NAND2_X1 U789 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U790 ( .A(n734), .B(G116), .ZN(G18) );
  XNOR2_X1 U791 ( .A(KEYINPUT117), .B(KEYINPUT37), .ZN(n736) );
  XNOR2_X1 U792 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U793 ( .A(G125), .B(n737), .ZN(G27) );
  XNOR2_X1 U794 ( .A(G134), .B(n738), .ZN(G36) );
  XOR2_X1 U795 ( .A(G140), .B(n739), .Z(G42) );
  XOR2_X1 U796 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n741) );
  NAND2_X1 U797 ( .A1(n749), .A2(G469), .ZN(n740) );
  BUF_X1 U798 ( .A(n742), .Z(n743) );
  NAND2_X1 U799 ( .A1(n746), .A2(G475), .ZN(n745) );
  NAND2_X1 U800 ( .A1(G478), .A2(n749), .ZN(n747) );
  NAND2_X1 U801 ( .A1(G217), .A2(n749), .ZN(n750) );
  NAND2_X1 U802 ( .A1(G953), .A2(G224), .ZN(n753) );
  XNOR2_X1 U803 ( .A(KEYINPUT61), .B(n753), .ZN(n754) );
  NAND2_X1 U804 ( .A1(n754), .A2(G898), .ZN(n755) );
  NAND2_X1 U805 ( .A1(n756), .A2(n755), .ZN(n760) );
  NOR2_X1 U806 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U807 ( .A(n760), .B(n759), .ZN(G69) );
  BUF_X1 U808 ( .A(n761), .Z(n762) );
  XNOR2_X1 U809 ( .A(n763), .B(n762), .ZN(n767) );
  NAND2_X1 U810 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U811 ( .A(KEYINPUT124), .B(n766), .ZN(n773) );
  XNOR2_X1 U812 ( .A(n767), .B(G227), .ZN(n768) );
  XNOR2_X1 U813 ( .A(n768), .B(KEYINPUT125), .ZN(n769) );
  NAND2_X1 U814 ( .A1(n769), .A2(G900), .ZN(n770) );
  NAND2_X1 U815 ( .A1(G953), .A2(n770), .ZN(n771) );
  XNOR2_X1 U816 ( .A(KEYINPUT126), .B(n771), .ZN(n772) );
  NAND2_X1 U817 ( .A1(n773), .A2(n772), .ZN(G72) );
  XNOR2_X1 U818 ( .A(G122), .B(n774), .ZN(G24) );
  XNOR2_X1 U819 ( .A(G119), .B(KEYINPUT127), .ZN(n775) );
  XNOR2_X1 U820 ( .A(G131), .B(n776), .ZN(G33) );
  XNOR2_X1 U821 ( .A(G137), .B(n356), .ZN(G39) );
endmodule

