//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954;
  INV_X1    g000(.A(G113gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G120gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT70), .B(G120gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(new_n202), .ZN(new_n205));
  AND2_X1   g004(.A1(G127gat), .A2(G134gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(G127gat), .A2(G134gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT71), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G127gat), .ZN(new_n209));
  INV_X1    g008(.A(G134gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT71), .ZN(new_n212));
  NAND2_X1  g011(.A1(G127gat), .A2(G134gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n208), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G120gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(G113gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n202), .A2(G120gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT69), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(G113gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT69), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n203), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n215), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n206), .A2(new_n207), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n205), .A2(new_n216), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(G169gat), .A3(G176gat), .ZN(new_n230));
  INV_X1    g029(.A(G169gat), .ZN(new_n231));
  INV_X1    g030(.A(G176gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n228), .A2(new_n230), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT23), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n241), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n235), .A2(new_n240), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n247), .B1(new_n246), .B2(new_n248), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n240), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n242), .A2(KEYINPUT25), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n249), .A2(new_n250), .A3(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n228), .A2(new_n230), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT26), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G183gat), .ZN(new_n260));
  INV_X1    g059(.A(G190gat), .ZN(new_n261));
  OAI22_X1  g060(.A1(new_n255), .A2(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n260), .A2(KEYINPUT27), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT27), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G183gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n261), .B1(KEYINPUT67), .B2(KEYINPUT28), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT68), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n268), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT27), .B(G183gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n262), .B1(new_n263), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n269), .A2(new_n273), .A3(KEYINPUT67), .A4(KEYINPUT28), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n226), .B1(new_n254), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G227gat), .ZN(new_n279));
  INV_X1    g078(.A(G233gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n246), .A2(new_n248), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT66), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n284));
  INV_X1    g083(.A(new_n253), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G113gat), .B(G120gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n215), .B1(new_n287), .B2(new_n222), .ZN(new_n288));
  INV_X1    g087(.A(new_n223), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n225), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n205), .A2(new_n215), .A3(new_n214), .A4(new_n208), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n276), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n286), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n281), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT33), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G15gat), .B(G43gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(G71gat), .B(G99gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n296), .B1(new_n302), .B2(KEYINPUT33), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n295), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n304), .B1(new_n295), .B2(new_n305), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT34), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n278), .A2(new_n294), .ZN(new_n310));
  INV_X1    g109(.A(new_n281), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI211_X1 g111(.A(KEYINPUT34), .B(new_n281), .C1(new_n278), .C2(new_n294), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n308), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n314), .B(new_n303), .C1(new_n307), .C2(new_n306), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT73), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT36), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n301), .B1(new_n295), .B2(new_n297), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n295), .A2(new_n305), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT72), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n295), .A2(new_n304), .A3(new_n305), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(new_n314), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n318), .A2(new_n319), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT36), .ZN(new_n328));
  XOR2_X1   g127(.A(G1gat), .B(G29gat), .Z(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G57gat), .B(G85gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G141gat), .B(G148gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT2), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(G155gat), .B2(G162gat), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n337), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G141gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G148gat), .ZN(new_n343));
  INV_X1    g142(.A(G148gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G141gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G155gat), .B(G162gat), .ZN(new_n347));
  INV_X1    g146(.A(G155gat), .ZN(new_n348));
  INV_X1    g147(.A(G162gat), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT2), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n341), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n225), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n203), .A2(new_n221), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT1), .B1(new_n354), .B2(KEYINPUT69), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n353), .B1(new_n355), .B2(new_n223), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n208), .A2(new_n214), .A3(new_n215), .ZN(new_n357));
  AND2_X1   g156(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n218), .B1(new_n360), .B2(G113gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n352), .B1(new_n356), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n341), .A2(new_n351), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(new_n290), .A3(new_n291), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(KEYINPUT78), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n292), .A2(new_n369), .A3(new_n352), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n366), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n372));
  AND4_X1   g171(.A1(new_n372), .A2(new_n364), .A3(new_n290), .A4(new_n291), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n372), .B1(new_n226), .B2(new_n364), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n341), .A2(new_n351), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n352), .A2(KEYINPUT3), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n292), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n373), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  OAI211_X1 g178(.A(KEYINPUT5), .B(new_n371), .C1(new_n379), .C2(new_n368), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n376), .ZN(new_n381));
  OAI211_X1 g180(.A(KEYINPUT4), .B(new_n365), .C1(new_n381), .C2(new_n226), .ZN(new_n382));
  INV_X1    g181(.A(new_n373), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n368), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT5), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n334), .B1(new_n380), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT6), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n380), .A2(new_n386), .A3(new_n334), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n391), .A2(new_n392), .A3(new_n387), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n380), .A2(new_n386), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n333), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n333), .B1(new_n384), .B2(new_n385), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT6), .B1(new_n396), .B2(new_n380), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT80), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n388), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT76), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT29), .B1(new_n286), .B2(new_n293), .ZN(new_n401));
  NAND2_X1  g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n400), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(G211gat), .A2(G218gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(G211gat), .A2(G218gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(KEYINPUT75), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT75), .ZN(new_n409));
  INV_X1    g208(.A(new_n407), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(new_n405), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT74), .ZN(new_n412));
  INV_X1    g211(.A(G197gat), .ZN(new_n413));
  INV_X1    g212(.A(G204gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G197gat), .A2(G204gat), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT22), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n415), .A2(new_n416), .B1(new_n417), .B2(new_n407), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n416), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n420), .B1(KEYINPUT22), .B2(new_n410), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n421), .A2(KEYINPUT74), .A3(new_n411), .A4(new_n408), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n286), .A2(new_n293), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(new_n403), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n253), .B1(new_n282), .B2(KEYINPUT66), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n427), .A2(new_n284), .B1(new_n276), .B2(new_n275), .ZN(new_n428));
  OAI211_X1 g227(.A(KEYINPUT76), .B(new_n402), .C1(new_n428), .C2(KEYINPUT29), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n404), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT29), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n403), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n428), .A2(new_n402), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n424), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  XOR2_X1   g233(.A(G8gat), .B(G36gat), .Z(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(KEYINPUT77), .ZN(new_n436));
  XNOR2_X1  g235(.A(G64gat), .B(G92gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n430), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT30), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n430), .A2(new_n434), .A3(KEYINPUT30), .A4(new_n439), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n430), .A2(new_n434), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n438), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n399), .A2(new_n446), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n376), .A2(new_n431), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n448), .A2(new_n423), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT29), .B1(new_n419), .B2(new_n422), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n352), .B1(new_n450), .B2(KEYINPUT3), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G228gat), .A2(G233gat), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n448), .A2(new_n423), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n408), .A2(new_n411), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n421), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n418), .A2(new_n408), .A3(new_n411), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n431), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n364), .B1(new_n460), .B2(new_n375), .ZN(new_n461));
  OR3_X1    g260(.A1(new_n456), .A2(new_n461), .A3(new_n454), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT31), .B(G50gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n455), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n453), .B1(new_n449), .B2(new_n451), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n456), .A2(new_n461), .A3(new_n454), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G78gat), .B(G106gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(G22gat), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n465), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n470), .B1(new_n465), .B2(new_n468), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n327), .A2(new_n328), .B1(new_n447), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT81), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n442), .A2(new_n445), .A3(KEYINPUT81), .A4(new_n443), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n379), .A2(new_n368), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(KEYINPUT39), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(new_n333), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n366), .A2(new_n370), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n480), .B(KEYINPUT39), .C1(new_n368), .C2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n482), .A2(KEYINPUT40), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT40), .B1(new_n482), .B2(new_n484), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n485), .A2(new_n486), .A3(new_n387), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n478), .A2(new_n479), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n438), .B1(new_n444), .B2(KEYINPUT37), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT37), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n430), .B2(new_n434), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT38), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n395), .A2(new_n397), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n493), .A2(new_n388), .A3(new_n440), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n432), .A2(new_n433), .A3(new_n424), .ZN(new_n495));
  INV_X1    g294(.A(new_n433), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n404), .A2(new_n496), .A3(new_n429), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n424), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT82), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(KEYINPUT82), .A3(new_n424), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n490), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT38), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n503), .B(new_n438), .C1(new_n444), .C2(KEYINPUT37), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n492), .B(new_n494), .C1(new_n502), .C2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n505), .A3(new_n473), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n475), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n388), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n392), .B1(new_n391), .B2(new_n387), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n395), .A2(new_n397), .A3(KEYINPUT80), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(new_n476), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n473), .B1(new_n324), .B2(new_n314), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n308), .A2(new_n315), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT83), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT83), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n316), .A2(new_n317), .A3(new_n516), .A4(new_n473), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n512), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n318), .A2(new_n326), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n493), .A2(new_n388), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT35), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(new_n473), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n478), .B2(new_n479), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n518), .A2(KEYINPUT35), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n507), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT16), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(G1gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(G1gat), .B2(new_n526), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n529), .B(G8gat), .Z(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NOR3_X1   g331(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT87), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(KEYINPUT87), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT88), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n533), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(KEYINPUT88), .A3(new_n537), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n540), .A2(new_n541), .B1(G29gat), .B2(G36gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(G43gat), .B(G50gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT15), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n533), .B(KEYINPUT90), .Z(new_n545));
  AND2_X1   g344(.A1(new_n545), .A2(new_n538), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n547));
  XOR2_X1   g346(.A(KEYINPUT89), .B(G50gat), .Z(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(new_n548), .B2(G43gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(G29gat), .A2(G36gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(new_n544), .A3(new_n550), .ZN(new_n551));
  OAI221_X1 g350(.A(new_n532), .B1(new_n542), .B2(new_n544), .C1(new_n546), .C2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n542), .A2(new_n544), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n551), .B1(new_n538), .B2(new_n545), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT17), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n531), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n553), .A2(new_n554), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(new_n530), .ZN(new_n558));
  NAND2_X1  g357(.A1(G229gat), .A2(G233gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n556), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n557), .B(new_n530), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n559), .B(KEYINPUT13), .Z(new_n566));
  AOI22_X1  g365(.A1(new_n561), .A2(KEYINPUT18), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G169gat), .B(G197gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT85), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G113gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT86), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G141gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n570), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT12), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n564), .B(new_n567), .C1(KEYINPUT92), .C2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n555), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT17), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n530), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n558), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n579), .A2(KEYINPUT18), .A3(new_n580), .A4(new_n559), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n581), .B(new_n582), .C1(new_n561), .C2(new_n563), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(KEYINPUT92), .A3(new_n582), .ZN(new_n584));
  INV_X1    g383(.A(new_n575), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n576), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n525), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT93), .ZN(new_n591));
  NAND2_X1  g390(.A1(G71gat), .A2(G78gat), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G57gat), .B(G64gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n591), .A2(KEYINPUT9), .ZN(new_n595));
  OAI221_X1 g394(.A(new_n593), .B1(new_n591), .B2(new_n592), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G64gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(G57gat), .ZN(new_n598));
  XOR2_X1   g397(.A(KEYINPUT94), .B(G57gat), .Z(new_n599));
  OAI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(new_n597), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n590), .A2(KEYINPUT9), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n592), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n600), .A2(KEYINPUT95), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT95), .B1(new_n600), .B2(new_n602), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n596), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n607));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  AOI21_X1  g408(.A(new_n531), .B1(new_n606), .B2(KEYINPUT21), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT97), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT96), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n613), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n611), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G190gat), .B(G218gat), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G85gat), .A2(G92gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT7), .ZN(new_n624));
  NAND2_X1  g423(.A1(G99gat), .A2(G106gat), .ZN(new_n625));
  INV_X1    g424(.A(G85gat), .ZN(new_n626));
  INV_X1    g425(.A(G92gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(KEYINPUT8), .A2(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G99gat), .B(G106gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n632), .B1(new_n577), .B2(new_n578), .ZN(new_n633));
  INV_X1    g432(.A(new_n557), .ZN(new_n634));
  AND2_X1   g433(.A1(G232gat), .A2(G233gat), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n634), .A2(new_n631), .B1(KEYINPUT41), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n622), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G134gat), .B(G162gat), .Z(new_n639));
  NOR2_X1   g438(.A1(new_n635), .A2(KEYINPUT41), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(KEYINPUT98), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n633), .A2(new_n636), .A3(new_n622), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n638), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n641), .B(KEYINPUT98), .Z(new_n645));
  INV_X1    g444(.A(new_n643), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n645), .B1(new_n646), .B2(new_n637), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n620), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n605), .A2(new_n632), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n631), .B(new_n596), .C1(new_n604), .C2(new_n603), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n631), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G230gat), .A2(G233gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n657), .B1(new_n651), .B2(new_n652), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n664), .B(new_n665), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n666), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n658), .A2(new_n660), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n667), .A2(KEYINPUT101), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT101), .B1(new_n667), .B2(new_n669), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n650), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n589), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n399), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT102), .B(G1gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1324gat));
  INV_X1    g478(.A(new_n676), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n478), .A2(new_n479), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT16), .B(G8gat), .Z(new_n683));
  NAND4_X1  g482(.A1(new_n680), .A2(KEYINPUT42), .A3(new_n682), .A4(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT104), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n680), .A2(new_n682), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n683), .B2(KEYINPUT103), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(KEYINPUT103), .B2(new_n683), .ZN(new_n689));
  OAI22_X1  g488(.A1(new_n686), .A2(new_n689), .B1(new_n687), .B2(G8gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n685), .A2(new_n690), .ZN(G1325gat));
  INV_X1    g490(.A(new_n519), .ZN(new_n692));
  OR3_X1    g491(.A1(new_n676), .A2(G15gat), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n327), .A2(new_n328), .ZN(new_n694));
  OAI21_X1  g493(.A(G15gat), .B1(new_n676), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(G1326gat));
  NOR2_X1   g495(.A1(new_n676), .A2(new_n473), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT43), .B(G22gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(new_n673), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n619), .A2(new_n700), .A3(new_n648), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT105), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n589), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n703), .A2(G29gat), .A3(new_n399), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT45), .Z(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n474), .B1(new_n511), .B2(new_n476), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT107), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n474), .B(new_n709), .C1(new_n511), .C2(new_n476), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n708), .A2(new_n710), .B1(new_n327), .B2(new_n328), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n518), .A2(KEYINPUT35), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n523), .A2(new_n519), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n711), .A2(new_n506), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n706), .B1(new_n714), .B2(new_n648), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n648), .A2(new_n706), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n507), .B2(new_n524), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n673), .B(KEYINPUT106), .Z(new_n718));
  NOR3_X1   g517(.A1(new_n718), .A2(new_n588), .A3(new_n619), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n715), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G29gat), .B1(new_n720), .B2(new_n399), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n721), .ZN(G1328gat));
  NOR3_X1   g521(.A1(new_n703), .A2(G36gat), .A3(new_n681), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT46), .ZN(new_n724));
  OAI21_X1  g523(.A(G36gat), .B1(new_n720), .B2(new_n681), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1329gat));
  NOR2_X1   g525(.A1(new_n703), .A2(new_n692), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n327), .A2(G43gat), .A3(new_n328), .ZN(new_n728));
  OAI22_X1  g527(.A1(new_n727), .A2(G43gat), .B1(new_n720), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g529(.A1(new_n703), .A2(new_n473), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n474), .A2(new_n548), .ZN(new_n732));
  OAI22_X1  g531(.A1(new_n731), .A2(new_n548), .B1(new_n720), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g533(.A(new_n709), .B1(new_n447), .B2(new_n474), .ZN(new_n735));
  INV_X1    g534(.A(new_n710), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n506), .B(new_n694), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n712), .A2(new_n713), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n718), .A2(new_n588), .A3(new_n650), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n511), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(new_n599), .ZN(G1332gat));
  NOR2_X1   g543(.A1(new_n741), .A2(new_n681), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  AND2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n745), .B2(new_n746), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT108), .ZN(G1333gat));
  OR3_X1    g549(.A1(new_n741), .A2(G71gat), .A3(new_n692), .ZN(new_n751));
  OAI21_X1  g550(.A(G71gat), .B1(new_n741), .B2(new_n694), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n742), .A2(new_n474), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  OAI21_X1  g556(.A(KEYINPUT112), .B1(new_n714), .B2(new_n648), .ZN(new_n758));
  OR3_X1    g557(.A1(new_n619), .A2(KEYINPUT110), .A3(new_n587), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT110), .B1(new_n619), .B2(new_n587), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n739), .A2(new_n762), .A3(new_n649), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n758), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n758), .A2(new_n763), .A3(KEYINPUT51), .A4(new_n761), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n768), .A2(new_n626), .A3(new_n511), .A4(new_n700), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n673), .B1(new_n759), .B2(new_n760), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n648), .B1(new_n737), .B2(new_n738), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n717), .B(new_n770), .C1(new_n771), .C2(KEYINPUT44), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n715), .A2(new_n774), .A3(new_n717), .A4(new_n770), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776), .B2(new_n399), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n769), .A2(new_n777), .ZN(G1336gat));
  INV_X1    g577(.A(new_n718), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n682), .A2(new_n627), .ZN(new_n780));
  AOI211_X1 g579(.A(new_n779), .B(new_n780), .C1(new_n766), .C2(new_n767), .ZN(new_n781));
  INV_X1    g580(.A(new_n772), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n627), .B1(new_n782), .B2(new_n682), .ZN(new_n783));
  OR3_X1    g582(.A1(new_n781), .A2(KEYINPUT52), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n773), .A2(new_n682), .A3(new_n775), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n785), .A2(new_n786), .A3(G92gat), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(new_n785), .B2(G92gat), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n787), .A2(new_n781), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n784), .B1(new_n789), .B2(new_n790), .ZN(G1337gat));
  NOR3_X1   g590(.A1(new_n692), .A2(new_n673), .A3(G99gat), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n768), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G99gat), .B1(new_n776), .B2(new_n694), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(G1338gat));
  AOI21_X1  g594(.A(new_n779), .B1(new_n766), .B2(new_n767), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n473), .A2(G106gat), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n474), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT53), .B1(new_n799), .B2(G106gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n773), .A2(new_n474), .A3(new_n775), .ZN(new_n802));
  AOI22_X1  g601(.A1(new_n796), .A2(new_n797), .B1(G106gat), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(G1339gat));
  XNOR2_X1  g604(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n666), .B1(new_n658), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n656), .B2(new_n657), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n654), .A2(G230gat), .A3(G233gat), .A4(new_n655), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n812), .B1(new_n811), .B2(new_n813), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n809), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n809), .B(KEYINPUT55), .C1(new_n814), .C2(new_n815), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n587), .A2(new_n818), .A3(new_n669), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n559), .B1(new_n579), .B2(new_n580), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n565), .A2(new_n566), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n574), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n564), .A2(new_n567), .A3(new_n575), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n823), .B(new_n824), .C1(new_n671), .C2(new_n672), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n649), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n818), .A2(new_n669), .A3(new_n819), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n824), .A2(new_n644), .A3(new_n647), .A4(new_n823), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n620), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n650), .A2(new_n588), .A3(new_n673), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n682), .A2(new_n399), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n832), .A2(new_n473), .A3(new_n519), .A4(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G113gat), .B1(new_n834), .B2(new_n588), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n833), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n515), .A2(new_n517), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n587), .A2(new_n202), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT116), .Z(G1340gat));
  OAI21_X1  g641(.A(G120gat), .B1(new_n834), .B2(new_n779), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n700), .A2(new_n360), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n839), .B2(new_n844), .ZN(G1341gat));
  OAI21_X1  g644(.A(G127gat), .B1(new_n834), .B2(new_n620), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n619), .A2(new_n209), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n839), .B2(new_n847), .ZN(G1342gat));
  NOR3_X1   g647(.A1(new_n839), .A2(G134gat), .A3(new_n648), .ZN(new_n849));
  XOR2_X1   g648(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n850));
  OR2_X1    g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  OAI21_X1  g651(.A(G134gat), .B1(new_n834), .B2(new_n648), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  AND4_X1   g653(.A1(new_n474), .A2(new_n832), .A3(new_n694), .A4(new_n833), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n342), .A3(new_n587), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(KEYINPUT118), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n833), .A2(new_n694), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n832), .A2(new_n474), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(KEYINPUT57), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n832), .A2(KEYINPUT57), .A3(new_n474), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n587), .B(new_n860), .C1(new_n863), .C2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n858), .B1(new_n866), .B2(G141gat), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n857), .A2(KEYINPUT118), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n867), .B(new_n868), .ZN(G1344gat));
  NAND3_X1  g668(.A1(new_n855), .A2(new_n344), .A3(new_n700), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n863), .A2(new_n865), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n700), .A3(new_n860), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n872), .A2(new_n873), .A3(G148gat), .ZN(new_n874));
  OR3_X1    g673(.A1(new_n826), .A2(KEYINPUT119), .A3(new_n829), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT119), .B1(new_n826), .B2(new_n829), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n876), .A3(new_n620), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n473), .B1(new_n877), .B2(new_n831), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n864), .B1(new_n878), .B2(KEYINPUT57), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n700), .A3(new_n860), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n873), .B1(new_n880), .B2(G148gat), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n870), .B1(new_n874), .B2(new_n881), .ZN(G1345gat));
  NAND3_X1  g681(.A1(new_n855), .A2(new_n348), .A3(new_n619), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n871), .A2(new_n619), .A3(new_n860), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n883), .B1(new_n885), .B2(new_n348), .ZN(G1346gat));
  OAI211_X1 g685(.A(new_n649), .B(new_n860), .C1(new_n863), .C2(new_n865), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n349), .B1(new_n887), .B2(KEYINPUT120), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(KEYINPUT120), .B2(new_n887), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n855), .A2(new_n349), .A3(new_n649), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1347gat));
  NOR2_X1   g690(.A1(new_n681), .A2(new_n511), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n832), .A2(new_n838), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n231), .A3(new_n587), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n894), .B(KEYINPUT121), .Z(new_n895));
  NOR3_X1   g694(.A1(new_n692), .A2(new_n511), .A3(new_n681), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n832), .A2(new_n473), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G169gat), .B1(new_n898), .B2(new_n588), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n895), .A2(new_n899), .ZN(G1348gat));
  OAI21_X1  g699(.A(G176gat), .B1(new_n898), .B2(new_n779), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n893), .A2(new_n232), .A3(new_n700), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1349gat));
  OAI21_X1  g702(.A(G183gat), .B1(new_n898), .B2(new_n620), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n893), .A2(new_n271), .A3(new_n619), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g706(.A(new_n261), .B1(new_n897), .B2(new_n649), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n910), .A2(KEYINPUT123), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  OR3_X1    g711(.A1(new_n908), .A2(new_n912), .A3(new_n909), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n908), .B2(new_n909), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n910), .A2(KEYINPUT123), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n911), .A2(new_n913), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n893), .A2(new_n261), .A3(new_n649), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1351gat));
  NAND2_X1  g717(.A1(new_n892), .A2(new_n694), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n861), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(G197gat), .B1(new_n920), .B2(new_n587), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n876), .A2(new_n620), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n826), .A2(KEYINPUT119), .A3(new_n829), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n831), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n474), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n865), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n919), .B(KEYINPUT124), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n588), .A2(new_n413), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n921), .B1(new_n929), .B2(new_n930), .ZN(G1352gat));
  NAND3_X1  g730(.A1(new_n920), .A2(new_n414), .A3(new_n700), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT62), .Z(new_n933));
  NOR3_X1   g732(.A1(new_n927), .A2(new_n779), .A3(new_n928), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n414), .B2(new_n934), .ZN(G1353gat));
  NOR2_X1   g734(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n919), .A2(new_n620), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT57), .B1(new_n924), .B2(new_n474), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n937), .B(new_n938), .C1(new_n939), .C2(new_n865), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G211gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n937), .B1(new_n879), .B2(new_n938), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n944));
  INV_X1    g743(.A(new_n938), .ZN(new_n945));
  OAI21_X1  g744(.A(KEYINPUT125), .B1(new_n927), .B2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n936), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n946), .A2(G211gat), .A3(new_n947), .A4(new_n940), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n943), .A2(new_n944), .A3(new_n948), .ZN(new_n949));
  OR3_X1    g748(.A1(new_n861), .A2(G211gat), .A3(new_n945), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1354gat));
  AOI21_X1  g750(.A(G218gat), .B1(new_n920), .B2(new_n649), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n649), .A2(G218gat), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT127), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n952), .B1(new_n929), .B2(new_n954), .ZN(G1355gat));
endmodule


