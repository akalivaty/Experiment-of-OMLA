

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593;

  XNOR2_X1 U326 ( .A(n363), .B(n362), .ZN(n566) );
  NOR2_X1 U327 ( .A1(n378), .A2(n584), .ZN(n380) );
  XNOR2_X1 U328 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U329 ( .A(n361), .B(n360), .ZN(n362) );
  AND2_X1 U330 ( .A1(G227GAT), .A2(G233GAT), .ZN(n294) );
  INV_X1 U331 ( .A(KEYINPUT118), .ZN(n379) );
  XNOR2_X1 U332 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U333 ( .A(G15GAT), .B(G127GAT), .Z(n330) );
  XOR2_X1 U334 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n349) );
  XNOR2_X1 U335 ( .A(n299), .B(n294), .ZN(n300) );
  XNOR2_X1 U336 ( .A(n351), .B(n350), .ZN(n352) );
  INV_X1 U337 ( .A(KEYINPUT37), .ZN(n481) );
  XNOR2_X1 U338 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U339 ( .A(n566), .B(KEYINPUT77), .ZN(n455) );
  XNOR2_X1 U340 ( .A(n484), .B(n483), .ZN(n527) );
  INV_X1 U341 ( .A(G43GAT), .ZN(n487) );
  XNOR2_X1 U342 ( .A(n310), .B(n404), .ZN(n541) );
  XNOR2_X1 U343 ( .A(n456), .B(KEYINPUT58), .ZN(n457) );
  XNOR2_X1 U344 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U345 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n490), .B(n489), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(G99GAT), .B(n330), .Z(n296) );
  XOR2_X1 U348 ( .A(G190GAT), .B(G134GAT), .Z(n354) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(n354), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n301) );
  XOR2_X1 U351 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n298) );
  XNOR2_X1 U352 ( .A(G113GAT), .B(G71GAT), .ZN(n297) );
  XNOR2_X1 U353 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U354 ( .A(n302), .B(G176GAT), .Z(n305) );
  XNOR2_X1 U355 ( .A(G120GAT), .B(KEYINPUT83), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n303), .B(KEYINPUT0), .ZN(n445) );
  XNOR2_X1 U357 ( .A(n445), .B(KEYINPUT20), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n310) );
  XOR2_X1 U359 ( .A(KEYINPUT86), .B(G183GAT), .Z(n307) );
  XNOR2_X1 U360 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n309) );
  XOR2_X1 U362 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n404) );
  XNOR2_X1 U364 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n311), .B(G29GAT), .ZN(n312) );
  XOR2_X1 U366 ( .A(n312), .B(KEYINPUT7), .Z(n314) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(G50GAT), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n357) );
  XNOR2_X1 U369 ( .A(G141GAT), .B(G113GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n315), .B(G1GAT), .ZN(n440) );
  XOR2_X1 U371 ( .A(G197GAT), .B(n440), .Z(n317) );
  NAND2_X1 U372 ( .A1(G229GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U374 ( .A(n318), .B(G22GAT), .Z(n326) );
  XOR2_X1 U375 ( .A(KEYINPUT29), .B(G8GAT), .Z(n320) );
  XNOR2_X1 U376 ( .A(G169GAT), .B(G15GAT), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U378 ( .A(KEYINPUT70), .B(KEYINPUT68), .Z(n322) );
  XNOR2_X1 U379 ( .A(KEYINPUT30), .B(KEYINPUT69), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U383 ( .A(n357), .B(n327), .Z(n580) );
  INV_X1 U384 ( .A(n580), .ZN(n515) );
  XNOR2_X1 U385 ( .A(KEYINPUT71), .B(n515), .ZN(n568) );
  XOR2_X1 U386 ( .A(KEYINPUT12), .B(KEYINPUT81), .Z(n329) );
  XNOR2_X1 U387 ( .A(KEYINPUT82), .B(KEYINPUT79), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n334) );
  XOR2_X1 U389 ( .A(G22GAT), .B(G155GAT), .Z(n414) );
  XOR2_X1 U390 ( .A(n414), .B(n330), .Z(n332) );
  XNOR2_X1 U391 ( .A(G1GAT), .B(G183GAT), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U393 ( .A(n334), .B(n333), .Z(n336) );
  NAND2_X1 U394 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U396 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n338) );
  XNOR2_X1 U397 ( .A(G64GAT), .B(KEYINPUT80), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U399 ( .A(n340), .B(n339), .Z(n345) );
  XNOR2_X1 U400 ( .A(G8GAT), .B(G211GAT), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n341), .B(KEYINPUT78), .ZN(n394) );
  XOR2_X1 U402 ( .A(KEYINPUT13), .B(G57GAT), .Z(n343) );
  XNOR2_X1 U403 ( .A(G71GAT), .B(G78GAT), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n370) );
  XNOR2_X1 U405 ( .A(n394), .B(n370), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n493) );
  XOR2_X1 U407 ( .A(G92GAT), .B(G85GAT), .Z(n347) );
  XNOR2_X1 U408 ( .A(G99GAT), .B(G106GAT), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n347), .B(n346), .ZN(n371) );
  XNOR2_X1 U410 ( .A(KEYINPUT67), .B(n371), .ZN(n353) );
  XNOR2_X1 U411 ( .A(KEYINPUT9), .B(KEYINPUT64), .ZN(n348) );
  XOR2_X1 U412 ( .A(n349), .B(n348), .Z(n351) );
  AND2_X1 U413 ( .A1(G232GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n356) );
  XOR2_X1 U415 ( .A(G218GAT), .B(G162GAT), .Z(n418) );
  XNOR2_X1 U416 ( .A(n354), .B(n418), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n363) );
  INV_X1 U418 ( .A(n357), .ZN(n361) );
  XOR2_X1 U419 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n359) );
  XNOR2_X1 U420 ( .A(KEYINPUT76), .B(KEYINPUT11), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U422 ( .A(KEYINPUT36), .B(n455), .ZN(n479) );
  NOR2_X1 U423 ( .A1(n493), .A2(n479), .ZN(n364) );
  XOR2_X1 U424 ( .A(KEYINPUT45), .B(n364), .Z(n378) );
  XOR2_X1 U425 ( .A(KEYINPUT73), .B(KEYINPUT33), .Z(n366) );
  XNOR2_X1 U426 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n377) );
  XOR2_X1 U428 ( .A(G204GAT), .B(G148GAT), .Z(n413) );
  XOR2_X1 U429 ( .A(G176GAT), .B(G64GAT), .Z(n395) );
  XNOR2_X1 U430 ( .A(n413), .B(n395), .ZN(n375) );
  XOR2_X1 U431 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n368) );
  NAND2_X1 U432 ( .A1(G230GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U434 ( .A(n369), .B(KEYINPUT72), .Z(n373) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n584) );
  NOR2_X1 U439 ( .A1(n568), .A2(n381), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n382), .B(KEYINPUT119), .ZN(n389) );
  XOR2_X1 U441 ( .A(KEYINPUT117), .B(KEYINPUT46), .Z(n384) );
  INV_X1 U442 ( .A(n584), .ZN(n485) );
  XNOR2_X1 U443 ( .A(KEYINPUT41), .B(n485), .ZN(n571) );
  NAND2_X1 U444 ( .A1(n580), .A2(n571), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U446 ( .A(KEYINPUT116), .B(n493), .ZN(n550) );
  NAND2_X1 U447 ( .A1(n385), .A2(n550), .ZN(n386) );
  NOR2_X1 U448 ( .A1(n566), .A2(n386), .ZN(n387) );
  XNOR2_X1 U449 ( .A(KEYINPUT47), .B(n387), .ZN(n388) );
  NAND2_X1 U450 ( .A1(n389), .A2(n388), .ZN(n391) );
  INV_X1 U451 ( .A(KEYINPUT48), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n391), .B(n390), .ZN(n538) );
  XOR2_X1 U453 ( .A(G92GAT), .B(G218GAT), .Z(n393) );
  XNOR2_X1 U454 ( .A(G36GAT), .B(G190GAT), .ZN(n392) );
  XNOR2_X1 U455 ( .A(n393), .B(n392), .ZN(n403) );
  XOR2_X1 U456 ( .A(n395), .B(n394), .Z(n397) );
  NAND2_X1 U457 ( .A1(G226GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U458 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U459 ( .A(n398), .B(KEYINPUT97), .Z(n401) );
  XNOR2_X1 U460 ( .A(G197GAT), .B(KEYINPUT90), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n399), .B(KEYINPUT21), .ZN(n426) );
  XNOR2_X1 U462 ( .A(n426), .B(G204GAT), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n529) );
  NOR2_X1 U466 ( .A1(n538), .A2(n529), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n406), .B(KEYINPUT54), .ZN(n576) );
  XOR2_X1 U468 ( .A(KEYINPUT22), .B(G78GAT), .Z(n408) );
  XNOR2_X1 U469 ( .A(G50GAT), .B(G106GAT), .ZN(n407) );
  XNOR2_X1 U470 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U471 ( .A(G211GAT), .B(KEYINPUT88), .Z(n410) );
  XNOR2_X1 U472 ( .A(G141GAT), .B(KEYINPUT89), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U474 ( .A(n412), .B(n411), .Z(n420) );
  XOR2_X1 U475 ( .A(n414), .B(n413), .Z(n416) );
  NAND2_X1 U476 ( .A1(G228GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U477 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U480 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n422) );
  XNOR2_X1 U481 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U483 ( .A(n424), .B(n423), .Z(n428) );
  XNOR2_X1 U484 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n425) );
  XNOR2_X1 U485 ( .A(n425), .B(KEYINPUT91), .ZN(n443) );
  XNOR2_X1 U486 ( .A(n443), .B(n426), .ZN(n427) );
  XNOR2_X1 U487 ( .A(n428), .B(n427), .ZN(n472) );
  XOR2_X1 U488 ( .A(KEYINPUT6), .B(G155GAT), .Z(n430) );
  XNOR2_X1 U489 ( .A(G127GAT), .B(G148GAT), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U491 ( .A(KEYINPUT96), .B(KEYINPUT4), .Z(n432) );
  XNOR2_X1 U492 ( .A(KEYINPUT94), .B(KEYINPUT1), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U494 ( .A(n434), .B(n433), .Z(n439) );
  XOR2_X1 U495 ( .A(G57GAT), .B(KEYINPUT5), .Z(n436) );
  NAND2_X1 U496 ( .A1(G225GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U497 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U498 ( .A(KEYINPUT95), .B(n437), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n449) );
  XOR2_X1 U500 ( .A(G85GAT), .B(G162GAT), .Z(n442) );
  XNOR2_X1 U501 ( .A(n440), .B(G134GAT), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U503 ( .A(n444), .B(n443), .Z(n447) );
  XNOR2_X1 U504 ( .A(G29GAT), .B(n445), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n577) );
  INV_X1 U507 ( .A(n577), .ZN(n450) );
  NOR2_X1 U508 ( .A1(n472), .A2(n450), .ZN(n451) );
  AND2_X1 U509 ( .A1(n576), .A2(n451), .ZN(n452) );
  XNOR2_X1 U510 ( .A(n452), .B(KEYINPUT55), .ZN(n453) );
  NOR2_X1 U511 ( .A1(n541), .A2(n453), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n454), .B(KEYINPUT124), .ZN(n572) );
  INV_X1 U513 ( .A(n572), .ZN(n459) );
  BUF_X1 U514 ( .A(n455), .Z(n554) );
  NOR2_X1 U515 ( .A1(n459), .A2(n554), .ZN(n458) );
  INV_X1 U516 ( .A(G190GAT), .ZN(n456) );
  NOR2_X1 U517 ( .A1(n459), .A2(n550), .ZN(n462) );
  INV_X1 U518 ( .A(KEYINPUT126), .ZN(n460) );
  XNOR2_X1 U519 ( .A(n460), .B(G183GAT), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n462), .B(n461), .ZN(G1350GAT) );
  NAND2_X1 U521 ( .A1(n472), .A2(n541), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n463), .B(KEYINPUT26), .ZN(n579) );
  INV_X1 U523 ( .A(n579), .ZN(n465) );
  XOR2_X1 U524 ( .A(KEYINPUT27), .B(KEYINPUT98), .Z(n464) );
  XNOR2_X1 U525 ( .A(n529), .B(n464), .ZN(n540) );
  NAND2_X1 U526 ( .A1(n465), .A2(n540), .ZN(n466) );
  NAND2_X1 U527 ( .A1(n466), .A2(n577), .ZN(n471) );
  NOR2_X1 U528 ( .A1(n541), .A2(n529), .ZN(n467) );
  NOR2_X1 U529 ( .A1(n472), .A2(n467), .ZN(n468) );
  XNOR2_X1 U530 ( .A(KEYINPUT25), .B(n468), .ZN(n469) );
  XNOR2_X1 U531 ( .A(KEYINPUT99), .B(n469), .ZN(n470) );
  NOR2_X1 U532 ( .A1(n471), .A2(n470), .ZN(n477) );
  XOR2_X1 U533 ( .A(n472), .B(KEYINPUT28), .Z(n542) );
  NAND2_X1 U534 ( .A1(n540), .A2(n542), .ZN(n474) );
  XNOR2_X1 U535 ( .A(KEYINPUT87), .B(n541), .ZN(n473) );
  NOR2_X1 U536 ( .A1(n474), .A2(n473), .ZN(n475) );
  NOR2_X1 U537 ( .A1(n475), .A2(n577), .ZN(n476) );
  NOR2_X1 U538 ( .A1(n477), .A2(n476), .ZN(n478) );
  XOR2_X1 U539 ( .A(KEYINPUT100), .B(n478), .Z(n496) );
  NOR2_X1 U540 ( .A1(n496), .A2(n479), .ZN(n480) );
  NAND2_X1 U541 ( .A1(n480), .A2(n493), .ZN(n484) );
  XOR2_X1 U542 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n482) );
  NAND2_X1 U543 ( .A1(n568), .A2(n485), .ZN(n498) );
  NOR2_X1 U544 ( .A1(n527), .A2(n498), .ZN(n486) );
  XOR2_X1 U545 ( .A(KEYINPUT38), .B(n486), .Z(n513) );
  NOR2_X1 U546 ( .A1(n541), .A2(n513), .ZN(n490) );
  XNOR2_X1 U547 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n488) );
  XOR2_X1 U548 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n492) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(n501) );
  INV_X1 U551 ( .A(n493), .ZN(n588) );
  NAND2_X1 U552 ( .A1(n554), .A2(n588), .ZN(n494) );
  XNOR2_X1 U553 ( .A(KEYINPUT16), .B(n494), .ZN(n495) );
  NOR2_X1 U554 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U555 ( .A(n497), .B(KEYINPUT101), .ZN(n516) );
  NOR2_X1 U556 ( .A1(n516), .A2(n498), .ZN(n499) );
  XOR2_X1 U557 ( .A(KEYINPUT102), .B(n499), .Z(n506) );
  NOR2_X1 U558 ( .A1(n506), .A2(n577), .ZN(n500) );
  XOR2_X1 U559 ( .A(n501), .B(n500), .Z(G1324GAT) );
  NOR2_X1 U560 ( .A1(n506), .A2(n529), .ZN(n502) );
  XOR2_X1 U561 ( .A(G8GAT), .B(n502), .Z(G1325GAT) );
  XNOR2_X1 U562 ( .A(KEYINPUT35), .B(KEYINPUT105), .ZN(n504) );
  NOR2_X1 U563 ( .A1(n541), .A2(n506), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U565 ( .A(G15GAT), .B(n505), .Z(G1326GAT) );
  NOR2_X1 U566 ( .A1(n542), .A2(n506), .ZN(n507) );
  XOR2_X1 U567 ( .A(G22GAT), .B(n507), .Z(G1327GAT) );
  NOR2_X1 U568 ( .A1(n513), .A2(n577), .ZN(n509) );
  XNOR2_X1 U569 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U571 ( .A(G29GAT), .B(n510), .ZN(G1328GAT) );
  NOR2_X1 U572 ( .A1(n513), .A2(n529), .ZN(n512) );
  XNOR2_X1 U573 ( .A(G36GAT), .B(KEYINPUT109), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n512), .B(n511), .ZN(G1329GAT) );
  NOR2_X1 U575 ( .A1(n542), .A2(n513), .ZN(n514) );
  XOR2_X1 U576 ( .A(G50GAT), .B(n514), .Z(G1331GAT) );
  XNOR2_X1 U577 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n520) );
  NAND2_X1 U578 ( .A1(n515), .A2(n571), .ZN(n526) );
  OR2_X1 U579 ( .A1(n516), .A2(n526), .ZN(n523) );
  NOR2_X1 U580 ( .A1(n577), .A2(n523), .ZN(n518) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(KEYINPUT112), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(G1332GAT) );
  NOR2_X1 U584 ( .A1(n529), .A2(n523), .ZN(n521) );
  XOR2_X1 U585 ( .A(G64GAT), .B(n521), .Z(G1333GAT) );
  NOR2_X1 U586 ( .A1(n541), .A2(n523), .ZN(n522) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n522), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n542), .A2(n523), .ZN(n525) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  OR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n534) );
  NOR2_X1 U592 ( .A1(n577), .A2(n534), .ZN(n528) );
  XOR2_X1 U593 ( .A(G85GAT), .B(n528), .Z(G1336GAT) );
  NOR2_X1 U594 ( .A1(n529), .A2(n534), .ZN(n531) );
  XNOR2_X1 U595 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n532), .B(G92GAT), .ZN(G1337GAT) );
  NOR2_X1 U598 ( .A1(n541), .A2(n534), .ZN(n533) );
  XOR2_X1 U599 ( .A(G99GAT), .B(n533), .Z(G1338GAT) );
  NOR2_X1 U600 ( .A1(n542), .A2(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(KEYINPUT44), .B(KEYINPUT115), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U603 ( .A(G106GAT), .B(n537), .ZN(G1339GAT) );
  NOR2_X1 U604 ( .A1(n577), .A2(n538), .ZN(n539) );
  NAND2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n558) );
  NOR2_X1 U606 ( .A1(n541), .A2(n558), .ZN(n543) );
  NAND2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U608 ( .A(KEYINPUT120), .B(n544), .Z(n549) );
  NAND2_X1 U609 ( .A1(n549), .A2(n568), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n545), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT121), .B(KEYINPUT49), .Z(n547) );
  NAND2_X1 U612 ( .A1(n549), .A2(n571), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U614 ( .A(G120GAT), .B(n548), .Z(G1341GAT) );
  INV_X1 U615 ( .A(n549), .ZN(n553) );
  NOR2_X1 U616 ( .A1(n553), .A2(n550), .ZN(n551) );
  XOR2_X1 U617 ( .A(KEYINPUT50), .B(n551), .Z(n552) );
  XNOR2_X1 U618 ( .A(G127GAT), .B(n552), .ZN(G1342GAT) );
  XNOR2_X1 U619 ( .A(KEYINPUT122), .B(KEYINPUT51), .ZN(n556) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G134GAT), .B(n557), .ZN(G1343GAT) );
  XOR2_X1 U623 ( .A(G141GAT), .B(KEYINPUT123), .Z(n560) );
  NOR2_X1 U624 ( .A1(n579), .A2(n558), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n565), .A2(n580), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1344GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n562) );
  NAND2_X1 U628 ( .A1(n565), .A2(n571), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(n563), .ZN(G1345GAT) );
  NAND2_X1 U631 ( .A1(n588), .A2(n565), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U635 ( .A(G169GAT), .B(KEYINPUT125), .Z(n570) );
  NAND2_X1 U636 ( .A1(n568), .A2(n572), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1348GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n574) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G176GAT), .B(n575), .ZN(G1349GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n582) );
  NAND2_X1 U643 ( .A1(n576), .A2(n577), .ZN(n578) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n590) );
  NAND2_X1 U645 ( .A1(n590), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U649 ( .A1(n590), .A2(n584), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(G204GAT), .B(n587), .Z(G1353GAT) );
  NAND2_X1 U652 ( .A1(n590), .A2(n588), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G211GAT), .B(n589), .ZN(G1354GAT) );
  INV_X1 U654 ( .A(n590), .ZN(n591) );
  NOR2_X1 U655 ( .A1(n479), .A2(n591), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(n592), .Z(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

