

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738;

  INV_X2 U367 ( .A(G953), .ZN(n728) );
  XNOR2_X1 U368 ( .A(G128), .B(G110), .ZN(n443) );
  XNOR2_X1 U369 ( .A(KEYINPUT67), .B(G131), .ZN(n426) );
  XNOR2_X1 U370 ( .A(n488), .B(n487), .ZN(n512) );
  INV_X1 U371 ( .A(n598), .ZN(n486) );
  XNOR2_X1 U372 ( .A(n531), .B(n530), .ZN(n672) );
  AND2_X2 U373 ( .A1(n356), .A2(n355), .ZN(n354) );
  NOR2_X2 U374 ( .A1(n517), .A2(n589), .ZN(n519) );
  NAND2_X2 U375 ( .A1(n354), .A2(n351), .ZN(n583) );
  AND2_X4 U376 ( .A1(n644), .A2(n643), .ZN(n716) );
  AND2_X1 U377 ( .A1(n563), .A2(n562), .ZN(n565) );
  NOR2_X1 U378 ( .A1(n562), .A2(n561), .ZN(n546) );
  NOR2_X1 U379 ( .A1(n719), .A2(G902), .ZN(n347) );
  XNOR2_X1 U380 ( .A(n367), .B(n366), .ZN(n562) );
  XNOR2_X1 U381 ( .A(n726), .B(G146), .ZN(n470) );
  XNOR2_X1 U382 ( .A(n428), .B(n427), .ZN(n726) );
  XNOR2_X1 U383 ( .A(n409), .B(n382), .ZN(n427) );
  XNOR2_X2 U384 ( .A(n347), .B(n348), .ZN(n545) );
  XOR2_X1 U385 ( .A(n472), .B(n471), .Z(n348) );
  INV_X1 U386 ( .A(n507), .ZN(n353) );
  INV_X1 U387 ( .A(G472), .ZN(n435) );
  XNOR2_X1 U388 ( .A(n601), .B(n600), .ZN(n614) );
  XNOR2_X1 U389 ( .A(n573), .B(n572), .ZN(n575) );
  INV_X1 U390 ( .A(KEYINPUT30), .ZN(n572) );
  NAND2_X1 U391 ( .A1(n353), .A2(n352), .ZN(n351) );
  NOR2_X1 U392 ( .A1(n506), .A2(KEYINPUT19), .ZN(n352) );
  XNOR2_X1 U393 ( .A(n567), .B(n361), .ZN(n585) );
  INV_X1 U394 ( .A(KEYINPUT22), .ZN(n369) );
  XNOR2_X1 U395 ( .A(n456), .B(n459), .ZN(n366) );
  NOR2_X1 U396 ( .A1(n673), .A2(G902), .ZN(n367) );
  INV_X1 U397 ( .A(KEYINPUT72), .ZN(n364) );
  XNOR2_X1 U398 ( .A(n376), .B(n375), .ZN(n509) );
  XNOR2_X1 U399 ( .A(KEYINPUT14), .B(KEYINPUT86), .ZN(n376) );
  XNOR2_X1 U400 ( .A(G143), .B(G113), .ZN(n392) );
  XNOR2_X1 U401 ( .A(KEYINPUT4), .B(G137), .ZN(n425) );
  XNOR2_X1 U402 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n408) );
  XNOR2_X1 U403 ( .A(G146), .B(G125), .ZN(n412) );
  OR2_X1 U404 ( .A1(n516), .A2(n515), .ZN(n520) );
  NOR2_X1 U405 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U406 ( .A(G137), .B(G119), .ZN(n446) );
  INV_X1 U407 ( .A(KEYINPUT9), .ZN(n378) );
  XNOR2_X1 U408 ( .A(G110), .B(G101), .ZN(n464) );
  NOR2_X1 U409 ( .A1(n651), .A2(n727), .ZN(n623) );
  XNOR2_X1 U410 ( .A(n614), .B(n602), .ZN(n604) );
  XNOR2_X1 U411 ( .A(n438), .B(n437), .ZN(n571) );
  XNOR2_X1 U412 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U413 ( .A(n433), .B(n403), .ZN(n357) );
  AND2_X1 U414 ( .A1(n647), .A2(G953), .ZN(n723) );
  INV_X1 U415 ( .A(n585), .ZN(n360) );
  NOR2_X1 U416 ( .A1(n585), .A2(n584), .ZN(n704) );
  INV_X1 U417 ( .A(KEYINPUT53), .ZN(n362) );
  NOR2_X1 U418 ( .A1(n632), .A2(n631), .ZN(n633) );
  AND2_X1 U419 ( .A1(n649), .A2(n648), .ZN(n349) );
  AND2_X1 U420 ( .A1(n363), .A2(n712), .ZN(n350) );
  XNOR2_X1 U421 ( .A(n452), .B(n724), .ZN(n673) );
  XNOR2_X1 U422 ( .A(n357), .B(n406), .ZN(n658) );
  NAND2_X1 U423 ( .A1(n353), .A2(n611), .ZN(n603) );
  NAND2_X1 U424 ( .A1(n506), .A2(KEYINPUT19), .ZN(n355) );
  NAND2_X1 U425 ( .A1(n507), .A2(KEYINPUT19), .ZN(n356) );
  XNOR2_X2 U426 ( .A(n359), .B(n358), .ZN(n433) );
  XNOR2_X2 U427 ( .A(KEYINPUT3), .B(G119), .ZN(n358) );
  XNOR2_X2 U428 ( .A(G101), .B(G113), .ZN(n359) );
  NAND2_X1 U429 ( .A1(n360), .A2(n545), .ZN(n568) );
  INV_X1 U430 ( .A(KEYINPUT28), .ZN(n361) );
  XNOR2_X1 U431 ( .A(n634), .B(n362), .ZN(G75) );
  NAND2_X1 U432 ( .A1(n608), .A2(n350), .ZN(n610) );
  XNOR2_X1 U433 ( .A(n365), .B(n364), .ZN(n363) );
  NAND2_X1 U434 ( .A1(n596), .A2(n595), .ZN(n365) );
  XNOR2_X2 U435 ( .A(n368), .B(n369), .ZN(n527) );
  NOR2_X2 U436 ( .A1(n541), .A2(n523), .ZN(n368) );
  XNOR2_X2 U437 ( .A(n370), .B(KEYINPUT0), .ZN(n541) );
  NAND2_X1 U438 ( .A1(n583), .A2(n511), .ZN(n370) );
  XNOR2_X1 U439 ( .A(n646), .B(n645), .ZN(n649) );
  NAND2_X1 U440 ( .A1(n716), .A2(G478), .ZN(n646) );
  NOR2_X2 U441 ( .A1(n699), .A2(n672), .ZN(n533) );
  BUF_X1 U442 ( .A(n635), .Z(n626) );
  XNOR2_X2 U443 ( .A(n421), .B(n420), .ZN(n507) );
  AND2_X1 U444 ( .A1(n735), .A2(n551), .ZN(n371) );
  XOR2_X1 U445 ( .A(n485), .B(KEYINPUT102), .Z(n372) );
  AND2_X1 U446 ( .A1(n575), .A2(n574), .ZN(n373) );
  INV_X1 U447 ( .A(KEYINPUT83), .ZN(n532) );
  XNOR2_X1 U448 ( .A(n533), .B(n532), .ZN(n534) );
  INV_X1 U449 ( .A(KEYINPUT44), .ZN(n535) );
  XNOR2_X1 U450 ( .A(n446), .B(n445), .ZN(n447) );
  INV_X1 U451 ( .A(KEYINPUT68), .ZN(n564) );
  XNOR2_X1 U452 ( .A(n379), .B(n378), .ZN(n380) );
  INV_X1 U453 ( .A(KEYINPUT109), .ZN(n602) );
  XNOR2_X1 U454 ( .A(n381), .B(n380), .ZN(n386) );
  INV_X1 U455 ( .A(KEYINPUT105), .ZN(n600) );
  INV_X1 U456 ( .A(KEYINPUT34), .ZN(n513) );
  BUF_X1 U457 ( .A(n637), .Z(n727) );
  INV_X1 U458 ( .A(KEYINPUT32), .ZN(n530) );
  XNOR2_X1 U459 ( .A(n580), .B(n579), .ZN(n736) );
  NAND2_X1 U460 ( .A1(G237), .A2(G234), .ZN(n375) );
  NAND2_X1 U461 ( .A1(G952), .A2(n509), .ZN(n508) );
  NAND2_X1 U462 ( .A1(G234), .A2(n728), .ZN(n377) );
  XOR2_X1 U463 ( .A(KEYINPUT8), .B(n377), .Z(n449) );
  NAND2_X1 U464 ( .A1(G217), .A2(n449), .ZN(n381) );
  XOR2_X1 U465 ( .A(KEYINPUT99), .B(KEYINPUT7), .Z(n379) );
  XNOR2_X2 U466 ( .A(G143), .B(G128), .ZN(n409) );
  INV_X1 U467 ( .A(G134), .ZN(n382) );
  XNOR2_X1 U468 ( .A(G107), .B(G116), .ZN(n403) );
  INV_X1 U469 ( .A(G122), .ZN(n383) );
  XNOR2_X1 U470 ( .A(n403), .B(n383), .ZN(n384) );
  XNOR2_X1 U471 ( .A(n427), .B(n384), .ZN(n385) );
  XNOR2_X1 U472 ( .A(n386), .B(n385), .ZN(n645) );
  INV_X1 U473 ( .A(G902), .ZN(n419) );
  NAND2_X1 U474 ( .A1(n645), .A2(n419), .ZN(n387) );
  XNOR2_X1 U475 ( .A(n387), .B(G478), .ZN(n516) );
  XOR2_X1 U476 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n389) );
  XNOR2_X1 U477 ( .A(KEYINPUT97), .B(KEYINPUT95), .ZN(n388) );
  XNOR2_X1 U478 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U479 ( .A(G104), .B(G122), .ZN(n405) );
  XNOR2_X1 U480 ( .A(n390), .B(n405), .ZN(n396) );
  NOR2_X1 U481 ( .A1(G953), .A2(G237), .ZN(n429) );
  NAND2_X1 U482 ( .A1(G214), .A2(n429), .ZN(n391) );
  XNOR2_X1 U483 ( .A(n391), .B(n426), .ZN(n394) );
  XNOR2_X1 U484 ( .A(n392), .B(KEYINPUT96), .ZN(n393) );
  XNOR2_X1 U485 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U486 ( .A(n396), .B(n395), .ZN(n400) );
  INV_X1 U487 ( .A(G140), .ZN(n397) );
  XNOR2_X1 U488 ( .A(n412), .B(n397), .ZN(n399) );
  XOR2_X1 U489 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n398) );
  XNOR2_X1 U490 ( .A(n399), .B(n398), .ZN(n724) );
  XNOR2_X1 U491 ( .A(n400), .B(n724), .ZN(n679) );
  NAND2_X1 U492 ( .A1(n679), .A2(n419), .ZN(n402) );
  XOR2_X1 U493 ( .A(KEYINPUT13), .B(G475), .Z(n401) );
  XNOR2_X1 U494 ( .A(n402), .B(n401), .ZN(n515) );
  XNOR2_X1 U495 ( .A(G110), .B(KEYINPUT16), .ZN(n404) );
  XNOR2_X1 U496 ( .A(n405), .B(n404), .ZN(n406) );
  NAND2_X1 U497 ( .A1(n728), .A2(G224), .ZN(n407) );
  XNOR2_X1 U498 ( .A(n408), .B(n407), .ZN(n410) );
  XNOR2_X1 U499 ( .A(n410), .B(n409), .ZN(n414) );
  XNOR2_X1 U500 ( .A(KEYINPUT4), .B(KEYINPUT76), .ZN(n411) );
  XNOR2_X1 U501 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U502 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U503 ( .A(n658), .B(n415), .ZN(n685) );
  XNOR2_X1 U504 ( .A(G902), .B(KEYINPUT85), .ZN(n417) );
  INV_X1 U505 ( .A(KEYINPUT15), .ZN(n416) );
  XNOR2_X1 U506 ( .A(n417), .B(n416), .ZN(n453) );
  INV_X1 U507 ( .A(n453), .ZN(n640) );
  OR2_X2 U508 ( .A1(n685), .A2(n640), .ZN(n421) );
  INV_X1 U509 ( .A(G237), .ZN(n418) );
  NAND2_X1 U510 ( .A1(n419), .A2(n418), .ZN(n422) );
  NAND2_X1 U511 ( .A1(n422), .A2(G210), .ZN(n420) );
  BUF_X1 U512 ( .A(n507), .Z(n617) );
  XOR2_X1 U513 ( .A(KEYINPUT38), .B(n617), .Z(n576) );
  INV_X1 U514 ( .A(n576), .ZN(n489) );
  NAND2_X1 U515 ( .A1(n422), .A2(G214), .ZN(n611) );
  NAND2_X1 U516 ( .A1(n489), .A2(n611), .ZN(n492) );
  NOR2_X1 U517 ( .A1(n520), .A2(n492), .ZN(n424) );
  XNOR2_X1 U518 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n423) );
  XNOR2_X1 U519 ( .A(n424), .B(n423), .ZN(n569) );
  XNOR2_X1 U520 ( .A(n426), .B(n425), .ZN(n428) );
  NAND2_X1 U521 ( .A1(n429), .A2(G210), .ZN(n431) );
  XNOR2_X1 U522 ( .A(G116), .B(KEYINPUT5), .ZN(n430) );
  XNOR2_X1 U523 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U524 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U525 ( .A(n470), .B(n434), .ZN(n666) );
  NOR2_X1 U526 ( .A1(G902), .A2(n666), .ZN(n438) );
  INV_X1 U527 ( .A(KEYINPUT71), .ZN(n436) );
  INV_X1 U528 ( .A(n571), .ZN(n566) );
  INV_X1 U529 ( .A(KEYINPUT23), .ZN(n439) );
  NAND2_X1 U530 ( .A1(KEYINPUT24), .A2(n439), .ZN(n442) );
  INV_X1 U531 ( .A(KEYINPUT24), .ZN(n440) );
  NAND2_X1 U532 ( .A1(n440), .A2(KEYINPUT23), .ZN(n441) );
  NAND2_X1 U533 ( .A1(n442), .A2(n441), .ZN(n444) );
  XNOR2_X1 U534 ( .A(n444), .B(n443), .ZN(n448) );
  INV_X1 U535 ( .A(KEYINPUT88), .ZN(n445) );
  XNOR2_X1 U536 ( .A(n448), .B(n447), .ZN(n451) );
  NAND2_X1 U537 ( .A1(n449), .A2(G221), .ZN(n450) );
  XNOR2_X1 U538 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U539 ( .A(KEYINPUT89), .B(KEYINPUT20), .Z(n455) );
  NAND2_X1 U540 ( .A1(G234), .A2(n453), .ZN(n454) );
  XNOR2_X1 U541 ( .A(n455), .B(n454), .ZN(n460) );
  NAND2_X1 U542 ( .A1(G217), .A2(n460), .ZN(n456) );
  XOR2_X1 U543 ( .A(KEYINPUT91), .B(KEYINPUT75), .Z(n458) );
  XNOR2_X1 U544 ( .A(KEYINPUT90), .B(KEYINPUT25), .ZN(n457) );
  XNOR2_X1 U545 ( .A(n458), .B(n457), .ZN(n459) );
  AND2_X1 U546 ( .A1(n460), .A2(G221), .ZN(n462) );
  INV_X1 U547 ( .A(KEYINPUT21), .ZN(n461) );
  XNOR2_X1 U548 ( .A(n462), .B(n461), .ZN(n561) );
  XNOR2_X1 U549 ( .A(G107), .B(KEYINPUT87), .ZN(n463) );
  XNOR2_X1 U550 ( .A(n464), .B(n463), .ZN(n468) );
  XNOR2_X1 U551 ( .A(G104), .B(G140), .ZN(n466) );
  NAND2_X1 U552 ( .A1(n728), .A2(G227), .ZN(n465) );
  XNOR2_X1 U553 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U554 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U555 ( .A(n470), .B(n469), .ZN(n719) );
  XNOR2_X1 U556 ( .A(KEYINPUT70), .B(G469), .ZN(n472) );
  INV_X1 U557 ( .A(KEYINPUT69), .ZN(n471) );
  XNOR2_X1 U558 ( .A(n545), .B(KEYINPUT1), .ZN(n474) );
  NAND2_X1 U559 ( .A1(n546), .A2(n474), .ZN(n485) );
  NOR2_X1 U560 ( .A1(n566), .A2(n485), .ZN(n473) );
  XOR2_X1 U561 ( .A(KEYINPUT93), .B(n473), .Z(n542) );
  INV_X1 U562 ( .A(n474), .ZN(n612) );
  INV_X1 U563 ( .A(n612), .ZN(n606) );
  NOR2_X1 U564 ( .A1(n546), .A2(n606), .ZN(n475) );
  XOR2_X1 U565 ( .A(KEYINPUT50), .B(n475), .Z(n479) );
  NAND2_X1 U566 ( .A1(n562), .A2(n561), .ZN(n476) );
  XNOR2_X1 U567 ( .A(n476), .B(KEYINPUT115), .ZN(n477) );
  XNOR2_X1 U568 ( .A(KEYINPUT49), .B(n477), .ZN(n478) );
  NAND2_X1 U569 ( .A1(n479), .A2(n478), .ZN(n480) );
  NOR2_X1 U570 ( .A1(n571), .A2(n480), .ZN(n481) );
  XNOR2_X1 U571 ( .A(n481), .B(KEYINPUT116), .ZN(n482) );
  NOR2_X1 U572 ( .A1(n542), .A2(n482), .ZN(n483) );
  XOR2_X1 U573 ( .A(KEYINPUT51), .B(n483), .Z(n484) );
  NOR2_X1 U574 ( .A1(n569), .A2(n484), .ZN(n499) );
  XNOR2_X1 U575 ( .A(n571), .B(KEYINPUT6), .ZN(n598) );
  NAND2_X1 U576 ( .A1(n372), .A2(n486), .ZN(n488) );
  XNOR2_X1 U577 ( .A(KEYINPUT103), .B(KEYINPUT33), .ZN(n487) );
  NOR2_X1 U578 ( .A1(n489), .A2(n611), .ZN(n490) );
  NOR2_X1 U579 ( .A1(n520), .A2(n490), .ZN(n495) );
  XOR2_X1 U580 ( .A(n515), .B(KEYINPUT98), .Z(n491) );
  NOR2_X1 U581 ( .A1(n491), .A2(n516), .ZN(n703) );
  INV_X1 U582 ( .A(n703), .ZN(n706) );
  AND2_X1 U583 ( .A1(n491), .A2(n516), .ZN(n700) );
  INV_X1 U584 ( .A(n700), .ZN(n708) );
  NAND2_X1 U585 ( .A1(n706), .A2(n708), .ZN(n586) );
  INV_X1 U586 ( .A(n586), .ZN(n493) );
  NOR2_X1 U587 ( .A1(n493), .A2(n492), .ZN(n494) );
  NOR2_X1 U588 ( .A1(n495), .A2(n494), .ZN(n496) );
  XOR2_X1 U589 ( .A(KEYINPUT117), .B(n496), .Z(n497) );
  NOR2_X1 U590 ( .A1(n512), .A2(n497), .ZN(n498) );
  NOR2_X1 U591 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U592 ( .A(n500), .B(KEYINPUT52), .ZN(n501) );
  NOR2_X1 U593 ( .A1(n508), .A2(n501), .ZN(n502) );
  XNOR2_X1 U594 ( .A(n502), .B(KEYINPUT118), .ZN(n504) );
  NOR2_X1 U595 ( .A1(n512), .A2(n569), .ZN(n503) );
  NOR2_X1 U596 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U597 ( .A(KEYINPUT119), .B(n505), .ZN(n632) );
  INV_X1 U598 ( .A(n611), .ZN(n506) );
  NOR2_X1 U599 ( .A1(n508), .A2(G953), .ZN(n558) );
  NAND2_X1 U600 ( .A1(G902), .A2(n509), .ZN(n554) );
  INV_X1 U601 ( .A(G898), .ZN(n655) );
  NAND2_X1 U602 ( .A1(G953), .A2(n655), .ZN(n659) );
  NOR2_X1 U603 ( .A1(n554), .A2(n659), .ZN(n510) );
  OR2_X1 U604 ( .A1(n558), .A2(n510), .ZN(n511) );
  NOR2_X1 U605 ( .A1(n512), .A2(n541), .ZN(n514) );
  XNOR2_X1 U606 ( .A(n514), .B(n513), .ZN(n517) );
  NAND2_X1 U607 ( .A1(n516), .A2(n515), .ZN(n589) );
  XOR2_X1 U608 ( .A(KEYINPUT77), .B(KEYINPUT35), .Z(n518) );
  XNOR2_X1 U609 ( .A(n519), .B(n518), .ZN(n650) );
  INV_X1 U610 ( .A(n520), .ZN(n522) );
  INV_X1 U611 ( .A(n561), .ZN(n521) );
  NAND2_X1 U612 ( .A1(n522), .A2(n521), .ZN(n523) );
  NAND2_X1 U613 ( .A1(n566), .A2(n612), .ZN(n524) );
  OR2_X2 U614 ( .A1(n527), .A2(n524), .ZN(n525) );
  XNOR2_X1 U615 ( .A(n525), .B(KEYINPUT65), .ZN(n526) );
  AND2_X2 U616 ( .A1(n526), .A2(n562), .ZN(n699) );
  NOR2_X2 U617 ( .A1(n486), .A2(n527), .ZN(n537) );
  NAND2_X1 U618 ( .A1(n606), .A2(n562), .ZN(n528) );
  XNOR2_X1 U619 ( .A(n528), .B(KEYINPUT101), .ZN(n529) );
  NAND2_X1 U620 ( .A1(n537), .A2(n529), .ZN(n531) );
  NAND2_X1 U621 ( .A1(n650), .A2(n534), .ZN(n536) );
  XNOR2_X1 U622 ( .A(n536), .B(n535), .ZN(n552) );
  XNOR2_X1 U623 ( .A(n537), .B(KEYINPUT82), .ZN(n539) );
  NOR2_X1 U624 ( .A1(n606), .A2(n562), .ZN(n538) );
  NAND2_X1 U625 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U626 ( .A(n540), .B(KEYINPUT100), .ZN(n735) );
  INV_X1 U627 ( .A(n541), .ZN(n548) );
  NAND2_X1 U628 ( .A1(n542), .A2(n548), .ZN(n544) );
  XOR2_X1 U629 ( .A(KEYINPUT31), .B(KEYINPUT94), .Z(n543) );
  XNOR2_X1 U630 ( .A(n544), .B(n543), .ZN(n709) );
  NAND2_X1 U631 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U632 ( .A(n547), .B(KEYINPUT92), .ZN(n591) );
  NOR2_X1 U633 ( .A1(n591), .A2(n571), .ZN(n549) );
  NAND2_X1 U634 ( .A1(n549), .A2(n548), .ZN(n694) );
  NAND2_X1 U635 ( .A1(n709), .A2(n694), .ZN(n550) );
  NAND2_X1 U636 ( .A1(n550), .A2(n586), .ZN(n551) );
  NAND2_X1 U637 ( .A1(n552), .A2(n371), .ZN(n553) );
  XNOR2_X1 U638 ( .A(n553), .B(KEYINPUT45), .ZN(n635) );
  INV_X1 U639 ( .A(n626), .ZN(n651) );
  XOR2_X1 U640 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n582) );
  NOR2_X1 U641 ( .A1(G900), .A2(n554), .ZN(n555) );
  NAND2_X1 U642 ( .A1(G953), .A2(n555), .ZN(n556) );
  XOR2_X1 U643 ( .A(KEYINPUT104), .B(n556), .Z(n557) );
  XOR2_X1 U644 ( .A(KEYINPUT78), .B(n559), .Z(n574) );
  INV_X1 U645 ( .A(n574), .ZN(n560) );
  NOR2_X1 U646 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U647 ( .A(n565), .B(n564), .ZN(n597) );
  NOR2_X1 U648 ( .A1(n597), .A2(n566), .ZN(n567) );
  NOR2_X1 U649 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U650 ( .A(KEYINPUT42), .B(n570), .Z(n738) );
  NAND2_X1 U651 ( .A1(n571), .A2(n611), .ZN(n573) );
  NOR2_X1 U652 ( .A1(n591), .A2(n576), .ZN(n577) );
  NAND2_X1 U653 ( .A1(n373), .A2(n577), .ZN(n578) );
  XNOR2_X1 U654 ( .A(KEYINPUT39), .B(n578), .ZN(n619) );
  NAND2_X1 U655 ( .A1(n619), .A2(n703), .ZN(n580) );
  XOR2_X1 U656 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n579) );
  NAND2_X1 U657 ( .A1(n738), .A2(n736), .ZN(n581) );
  XNOR2_X1 U658 ( .A(n582), .B(n581), .ZN(n608) );
  NAND2_X1 U659 ( .A1(n583), .A2(n545), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n704), .A2(n586), .ZN(n588) );
  NOR2_X1 U661 ( .A1(KEYINPUT73), .A2(KEYINPUT47), .ZN(n587) );
  XNOR2_X1 U662 ( .A(n588), .B(n587), .ZN(n596) );
  NAND2_X1 U663 ( .A1(KEYINPUT73), .A2(KEYINPUT47), .ZN(n594) );
  OR2_X1 U664 ( .A1(n589), .A2(n617), .ZN(n590) );
  NOR2_X1 U665 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n373), .A2(n592), .ZN(n593) );
  XNOR2_X1 U667 ( .A(KEYINPUT106), .B(n593), .ZN(n737) );
  AND2_X1 U668 ( .A1(n594), .A2(n737), .ZN(n595) );
  NOR2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n703), .A2(n599), .ZN(n601) );
  NOR2_X1 U671 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U672 ( .A(n605), .B(KEYINPUT36), .ZN(n607) );
  NAND2_X1 U673 ( .A1(n607), .A2(n606), .ZN(n712) );
  INV_X1 U674 ( .A(KEYINPUT48), .ZN(n609) );
  XNOR2_X1 U675 ( .A(n610), .B(n609), .ZN(n622) );
  NAND2_X1 U676 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U677 ( .A1(n614), .A2(n613), .ZN(n616) );
  INV_X1 U678 ( .A(KEYINPUT43), .ZN(n615) );
  XNOR2_X1 U679 ( .A(n616), .B(n615), .ZN(n618) );
  NAND2_X1 U680 ( .A1(n618), .A2(n617), .ZN(n664) );
  AND2_X1 U681 ( .A1(n700), .A2(n619), .ZN(n714) );
  INV_X1 U682 ( .A(n714), .ZN(n620) );
  AND2_X1 U683 ( .A1(n664), .A2(n620), .ZN(n621) );
  NAND2_X1 U684 ( .A1(n622), .A2(n621), .ZN(n637) );
  NOR2_X1 U685 ( .A1(n623), .A2(KEYINPUT2), .ZN(n629) );
  INV_X1 U686 ( .A(n637), .ZN(n624) );
  NAND2_X1 U687 ( .A1(n624), .A2(KEYINPUT2), .ZN(n625) );
  XNOR2_X1 U688 ( .A(n625), .B(KEYINPUT81), .ZN(n627) );
  NAND2_X1 U689 ( .A1(n627), .A2(n626), .ZN(n643) );
  INV_X1 U690 ( .A(n643), .ZN(n628) );
  NOR2_X1 U691 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U692 ( .A(KEYINPUT80), .B(n630), .ZN(n631) );
  NAND2_X1 U693 ( .A1(n633), .A2(n728), .ZN(n634) );
  NAND2_X1 U694 ( .A1(n635), .A2(n640), .ZN(n636) );
  XNOR2_X1 U695 ( .A(n636), .B(KEYINPUT79), .ZN(n639) );
  XOR2_X1 U696 ( .A(KEYINPUT74), .B(n637), .Z(n638) );
  NAND2_X1 U697 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U698 ( .A1(n640), .A2(KEYINPUT2), .ZN(n641) );
  NAND2_X1 U699 ( .A1(n642), .A2(n641), .ZN(n644) );
  INV_X1 U700 ( .A(G952), .ZN(n647) );
  INV_X1 U701 ( .A(n723), .ZN(n648) );
  XNOR2_X1 U702 ( .A(n349), .B(KEYINPUT124), .ZN(G63) );
  XNOR2_X1 U703 ( .A(n650), .B(G122), .ZN(G24) );
  NOR2_X1 U704 ( .A1(n651), .A2(G953), .ZN(n657) );
  NAND2_X1 U705 ( .A1(G224), .A2(G953), .ZN(n652) );
  XNOR2_X1 U706 ( .A(n652), .B(KEYINPUT61), .ZN(n653) );
  XNOR2_X1 U707 ( .A(n653), .B(KEYINPUT127), .ZN(n654) );
  NOR2_X1 U708 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U709 ( .A1(n657), .A2(n656), .ZN(n662) );
  INV_X1 U710 ( .A(n658), .ZN(n660) );
  NAND2_X1 U711 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U712 ( .A(n662), .B(n661), .ZN(G69) );
  XNOR2_X1 U713 ( .A(G140), .B(KEYINPUT114), .ZN(n663) );
  XNOR2_X1 U714 ( .A(n664), .B(n663), .ZN(G42) );
  INV_X1 U715 ( .A(KEYINPUT63), .ZN(n671) );
  NAND2_X1 U716 ( .A1(n716), .A2(G472), .ZN(n668) );
  XNOR2_X1 U717 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n665) );
  XNOR2_X1 U718 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U719 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X2 U720 ( .A1(n669), .A2(n723), .ZN(n670) );
  XNOR2_X1 U721 ( .A(n671), .B(n670), .ZN(G57) );
  XOR2_X1 U722 ( .A(n672), .B(G119), .Z(G21) );
  NAND2_X1 U723 ( .A1(n716), .A2(G217), .ZN(n675) );
  XOR2_X1 U724 ( .A(KEYINPUT125), .B(n673), .Z(n674) );
  XNOR2_X1 U725 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X2 U726 ( .A1(n676), .A2(n723), .ZN(n677) );
  XNOR2_X1 U727 ( .A(n677), .B(KEYINPUT126), .ZN(G66) );
  NAND2_X1 U728 ( .A1(n716), .A2(G475), .ZN(n681) );
  XNOR2_X1 U729 ( .A(KEYINPUT122), .B(KEYINPUT59), .ZN(n678) );
  XNOR2_X1 U730 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U731 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X2 U732 ( .A1(n682), .A2(n723), .ZN(n684) );
  XOR2_X1 U733 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n683) );
  XNOR2_X1 U734 ( .A(n684), .B(n683), .ZN(G60) );
  NAND2_X1 U735 ( .A1(n716), .A2(G210), .ZN(n689) );
  XOR2_X1 U736 ( .A(KEYINPUT84), .B(KEYINPUT54), .Z(n686) );
  XNOR2_X1 U737 ( .A(n686), .B(KEYINPUT55), .ZN(n687) );
  XNOR2_X1 U738 ( .A(n685), .B(n687), .ZN(n688) );
  XNOR2_X1 U739 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X2 U740 ( .A1(n690), .A2(n723), .ZN(n692) );
  XNOR2_X1 U741 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n691) );
  XNOR2_X1 U742 ( .A(n692), .B(n691), .ZN(G51) );
  NOR2_X1 U743 ( .A1(n706), .A2(n694), .ZN(n693) );
  XOR2_X1 U744 ( .A(G104), .B(n693), .Z(G6) );
  NOR2_X1 U745 ( .A1(n694), .A2(n708), .ZN(n698) );
  XOR2_X1 U746 ( .A(KEYINPUT26), .B(KEYINPUT111), .Z(n696) );
  XNOR2_X1 U747 ( .A(G107), .B(KEYINPUT27), .ZN(n695) );
  XNOR2_X1 U748 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U749 ( .A(n698), .B(n697), .ZN(G9) );
  XOR2_X1 U750 ( .A(n699), .B(G110), .Z(G12) );
  XOR2_X1 U751 ( .A(G128), .B(KEYINPUT29), .Z(n702) );
  NAND2_X1 U752 ( .A1(n704), .A2(n700), .ZN(n701) );
  XNOR2_X1 U753 ( .A(n702), .B(n701), .ZN(G30) );
  NAND2_X1 U754 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U755 ( .A(n705), .B(G146), .ZN(G48) );
  NOR2_X1 U756 ( .A1(n709), .A2(n706), .ZN(n707) );
  XOR2_X1 U757 ( .A(G113), .B(n707), .Z(G15) );
  NOR2_X1 U758 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U759 ( .A(KEYINPUT112), .B(n710), .Z(n711) );
  XNOR2_X1 U760 ( .A(G116), .B(n711), .ZN(G18) );
  XOR2_X1 U761 ( .A(n712), .B(G125), .Z(n713) );
  XNOR2_X1 U762 ( .A(n713), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U763 ( .A(G134), .B(n714), .ZN(n715) );
  XNOR2_X1 U764 ( .A(n715), .B(KEYINPUT113), .ZN(G36) );
  NAND2_X1 U765 ( .A1(n716), .A2(G469), .ZN(n721) );
  XOR2_X1 U766 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n717) );
  XOR2_X1 U767 ( .A(n717), .B(KEYINPUT121), .Z(n718) );
  XNOR2_X1 U768 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U769 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U770 ( .A1(n723), .A2(n722), .ZN(G54) );
  XNOR2_X1 U771 ( .A(n724), .B(KEYINPUT87), .ZN(n725) );
  XNOR2_X1 U772 ( .A(n726), .B(n725), .ZN(n730) );
  XNOR2_X1 U773 ( .A(n730), .B(n727), .ZN(n729) );
  NAND2_X1 U774 ( .A1(n729), .A2(n728), .ZN(n734) );
  XNOR2_X1 U775 ( .A(G227), .B(n730), .ZN(n731) );
  NAND2_X1 U776 ( .A1(n731), .A2(G900), .ZN(n732) );
  NAND2_X1 U777 ( .A1(G953), .A2(n732), .ZN(n733) );
  NAND2_X1 U778 ( .A1(n734), .A2(n733), .ZN(G72) );
  XNOR2_X1 U779 ( .A(G101), .B(n735), .ZN(G3) );
  XNOR2_X1 U780 ( .A(G131), .B(n736), .ZN(G33) );
  XNOR2_X1 U781 ( .A(G143), .B(n737), .ZN(G45) );
  XNOR2_X1 U782 ( .A(G137), .B(n738), .ZN(G39) );
endmodule

