

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814;

  BUF_X1 U368 ( .A(n636), .Z(n643) );
  XNOR2_X1 U369 ( .A(n432), .B(n386), .ZN(n461) );
  NOR2_X1 U370 ( .A1(n754), .A2(n753), .ZN(n638) );
  XNOR2_X1 U371 ( .A(n600), .B(n599), .ZN(n697) );
  XNOR2_X1 U372 ( .A(n368), .B(n506), .ZN(n458) );
  AND2_X1 U373 ( .A1(n453), .A2(n684), .ZN(n452) );
  XNOR2_X1 U374 ( .A(n551), .B(n362), .ZN(n636) );
  NOR2_X1 U375 ( .A1(n660), .A2(n659), .ZN(n423) );
  NOR2_X1 U376 ( .A1(n666), .A2(n753), .ZN(n390) );
  AND2_X1 U377 ( .A1(n378), .A2(n778), .ZN(n348) );
  NOR2_X1 U378 ( .A1(n458), .A2(n528), .ZN(n457) );
  NOR2_X1 U379 ( .A1(n439), .A2(n813), .ZN(n370) );
  AND2_X1 U380 ( .A1(n488), .A2(n485), .ZN(n484) );
  AND2_X1 U381 ( .A1(n487), .A2(n674), .ZN(n485) );
  NAND2_X1 U382 ( .A1(n490), .A2(n489), .ZN(n486) );
  NAND2_X1 U383 ( .A1(n636), .A2(n581), .ZN(n410) );
  XNOR2_X1 U384 ( .A(n635), .B(n634), .ZN(n773) );
  XNOR2_X1 U385 ( .A(n423), .B(KEYINPUT81), .ZN(n394) );
  XNOR2_X1 U386 ( .A(n621), .B(KEYINPUT38), .ZN(n661) );
  XNOR2_X1 U387 ( .A(n657), .B(KEYINPUT6), .ZN(n630) );
  AND2_X1 U388 ( .A1(n500), .A2(n499), .ZN(n498) );
  OR2_X1 U389 ( .A1(n733), .A2(n497), .ZN(n496) );
  XOR2_X1 U390 ( .A(G137), .B(KEYINPUT4), .Z(n583) );
  XNOR2_X1 U391 ( .A(G143), .B(G128), .ZN(n569) );
  XNOR2_X1 U392 ( .A(KEYINPUT101), .B(KEYINPUT82), .ZN(n416) );
  BUF_X1 U393 ( .A(n620), .Z(n621) );
  NOR2_X1 U394 ( .A1(n663), .A2(n662), .ZN(n665) );
  AND2_X1 U395 ( .A1(n347), .A2(n348), .ZN(n377) );
  NAND2_X1 U396 ( .A1(n509), .A2(n379), .ZN(n347) );
  NOR2_X2 U397 ( .A1(n451), .A2(n457), .ZN(n739) );
  NAND2_X1 U398 ( .A1(n455), .A2(n452), .ZN(n451) );
  NOR2_X1 U399 ( .A1(n739), .A2(KEYINPUT2), .ZN(n740) );
  XNOR2_X2 U400 ( .A(n656), .B(n350), .ZN(n349) );
  INV_X1 U401 ( .A(n349), .ZN(n738) );
  XOR2_X1 U402 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n350) );
  AND2_X2 U403 ( .A1(n731), .A2(G217), .ZN(n690) );
  XNOR2_X2 U404 ( .A(n465), .B(n363), .ZN(n450) );
  INV_X1 U405 ( .A(G104), .ZN(n537) );
  XNOR2_X1 U406 ( .A(KEYINPUT80), .B(G110), .ZN(n538) );
  NAND2_X1 U407 ( .A1(n661), .A2(n525), .ZN(n523) );
  NAND2_X1 U408 ( .A1(n394), .A2(n525), .ZN(n513) );
  XNOR2_X1 U409 ( .A(n391), .B(n531), .ZN(n407) );
  NAND2_X1 U410 ( .A1(n446), .A2(n532), .ZN(n391) );
  NAND2_X1 U411 ( .A1(G469), .A2(n426), .ZN(n497) );
  NAND2_X1 U412 ( .A1(n590), .A2(G902), .ZN(n499) );
  XNOR2_X1 U413 ( .A(n437), .B(n536), .ZN(n805) );
  XNOR2_X1 U414 ( .A(n596), .B(KEYINPUT16), .ZN(n437) );
  XNOR2_X1 U415 ( .A(n539), .B(n803), .ZN(n588) );
  NAND2_X1 U416 ( .A1(n790), .A2(n524), .ZN(n521) );
  XNOR2_X1 U417 ( .A(n628), .B(KEYINPUT98), .ZN(n650) );
  AND2_X1 U418 ( .A1(n527), .A2(n528), .ZN(n456) );
  XOR2_X1 U419 ( .A(G104), .B(G122), .Z(n554) );
  XNOR2_X1 U420 ( .A(G113), .B(G143), .ZN(n553) );
  XOR2_X1 U421 ( .A(KEYINPUT105), .B(KEYINPUT107), .Z(n556) );
  NAND2_X1 U422 ( .A1(n686), .A2(KEYINPUT2), .ZN(n529) );
  NAND2_X1 U423 ( .A1(n689), .A2(n426), .ZN(n507) );
  NOR2_X1 U424 ( .A1(n747), .A2(n402), .ZN(n401) );
  NOR2_X1 U425 ( .A1(n745), .A2(KEYINPUT41), .ZN(n400) );
  INV_X1 U426 ( .A(n521), .ZN(n517) );
  OR2_X2 U427 ( .A1(n428), .A2(n424), .ZN(n657) );
  NAND2_X1 U428 ( .A1(n430), .A2(n429), .ZN(n428) );
  NAND2_X1 U429 ( .A1(G902), .A2(G472), .ZN(n429) );
  XNOR2_X1 U430 ( .A(n568), .B(n567), .ZN(n606) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n568) );
  INV_X1 U432 ( .A(KEYINPUT88), .ZN(n373) );
  INV_X1 U433 ( .A(G107), .ZN(n534) );
  XNOR2_X1 U434 ( .A(G122), .B(G116), .ZN(n535) );
  XNOR2_X1 U435 ( .A(n564), .B(n563), .ZN(n431) );
  INV_X1 U436 ( .A(n588), .ZN(n414) );
  OR2_X1 U437 ( .A1(n505), .A2(n508), .ZN(n378) );
  INV_X1 U438 ( .A(KEYINPUT86), .ZN(n510) );
  AND2_X1 U439 ( .A1(n473), .A2(n744), .ZN(n406) );
  NOR2_X1 U440 ( .A1(n678), .A2(n361), .ZN(n473) );
  NAND2_X1 U441 ( .A1(n494), .A2(n492), .ZN(n754) );
  NAND2_X1 U442 ( .A1(n357), .A2(n498), .ZN(n494) );
  NAND2_X1 U443 ( .A1(n493), .A2(KEYINPUT1), .ZN(n492) );
  XNOR2_X1 U444 ( .A(n372), .B(G478), .ZN(n436) );
  NAND2_X1 U445 ( .A1(n695), .A2(n426), .ZN(n372) );
  INV_X1 U446 ( .A(n436), .ZN(n645) );
  NAND2_X1 U447 ( .A1(n521), .A2(KEYINPUT40), .ZN(n516) );
  NAND2_X1 U448 ( .A1(n682), .A2(n790), .ZN(n672) );
  NAND2_X1 U449 ( .A1(n650), .A2(KEYINPUT44), .ZN(n383) );
  INV_X1 U450 ( .A(KEYINPUT96), .ZN(n481) );
  INV_X1 U451 ( .A(n672), .ZN(n749) );
  NAND2_X1 U452 ( .A1(n454), .A2(KEYINPUT92), .ZN(n453) );
  INV_X1 U453 ( .A(KEYINPUT48), .ZN(n506) );
  INV_X1 U454 ( .A(G237), .ZN(n541) );
  NAND2_X1 U455 ( .A1(n427), .A2(n426), .ZN(n425) );
  INV_X1 U456 ( .A(G472), .ZN(n427) );
  XOR2_X1 U457 ( .A(G116), .B(KEYINPUT104), .Z(n593) );
  XNOR2_X1 U458 ( .A(n502), .B(n501), .ZN(n596) );
  XNOR2_X1 U459 ( .A(G119), .B(G113), .ZN(n502) );
  XNOR2_X1 U460 ( .A(KEYINPUT75), .B(KEYINPUT3), .ZN(n501) );
  XNOR2_X1 U461 ( .A(KEYINPUT8), .B(KEYINPUT70), .ZN(n374) );
  NOR2_X1 U462 ( .A1(G953), .A2(G237), .ZN(n591) );
  XNOR2_X1 U463 ( .A(KEYINPUT11), .B(KEYINPUT106), .ZN(n555) );
  NOR2_X1 U464 ( .A1(n687), .A2(n503), .ZN(n476) );
  INV_X1 U465 ( .A(n529), .ZN(n503) );
  NAND2_X1 U466 ( .A1(n529), .A2(KEYINPUT90), .ZN(n504) );
  AND2_X1 U467 ( .A1(n739), .A2(n448), .ZN(n478) );
  NOR2_X1 U468 ( .A1(n685), .A2(n449), .ZN(n448) );
  INV_X1 U469 ( .A(KEYINPUT90), .ZN(n449) );
  XNOR2_X1 U470 ( .A(n417), .B(n416), .ZN(n415) );
  XNOR2_X1 U471 ( .A(KEYINPUT17), .B(KEYINPUT4), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n420), .B(n569), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n633), .B(n632), .ZN(n634) );
  NAND2_X1 U474 ( .A1(n468), .A2(n467), .ZN(n466) );
  AND2_X1 U475 ( .A1(n757), .A2(n358), .ZN(n467) );
  INV_X1 U476 ( .A(KEYINPUT126), .ZN(n433) );
  INV_X1 U477 ( .A(G953), .ZN(n797) );
  XNOR2_X1 U478 ( .A(n604), .B(n603), .ZN(n605) );
  INV_X1 U479 ( .A(KEYINPUT102), .ZN(n603) );
  XNOR2_X1 U480 ( .A(n405), .B(n404), .ZN(n403) );
  INV_X1 U481 ( .A(KEYINPUT43), .ZN(n404) );
  NAND2_X1 U482 ( .A1(n399), .A2(n397), .ZN(n772) );
  NOR2_X1 U483 ( .A1(n400), .A2(n356), .ZN(n399) );
  XNOR2_X1 U484 ( .A(n793), .B(n434), .ZN(n682) );
  INV_X1 U485 ( .A(KEYINPUT111), .ZN(n434) );
  AND2_X1 U486 ( .A1(n441), .A2(n513), .ZN(n440) );
  NOR2_X1 U487 ( .A1(n517), .A2(n514), .ZN(n441) );
  INV_X1 U488 ( .A(n523), .ZN(n514) );
  AND2_X1 U489 ( .A1(n754), .A2(n630), .ZN(n408) );
  XOR2_X1 U490 ( .A(KEYINPUT62), .B(n697), .Z(n698) );
  XNOR2_X1 U491 ( .A(n576), .B(n575), .ZN(n695) );
  XNOR2_X1 U492 ( .A(n431), .B(n703), .ZN(n704) );
  XOR2_X1 U493 ( .A(G107), .B(G140), .Z(n585) );
  XNOR2_X1 U494 ( .A(n711), .B(n714), .ZN(n715) );
  INV_X1 U495 ( .A(G140), .ZN(n622) );
  NOR2_X2 U496 ( .A1(n470), .A2(n469), .ZN(n795) );
  NAND2_X1 U497 ( .A1(n472), .A2(n471), .ZN(n470) );
  NOR2_X1 U498 ( .A1(n680), .A2(n352), .ZN(n471) );
  XNOR2_X1 U499 ( .A(n675), .B(n393), .ZN(n392) );
  OR2_X1 U500 ( .A1(n394), .A2(n422), .ZN(n675) );
  NAND2_X1 U501 ( .A1(n674), .A2(n621), .ZN(n422) );
  INV_X1 U502 ( .A(G131), .ZN(n438) );
  XNOR2_X1 U503 ( .A(n392), .B(G143), .ZN(G45) );
  AND2_X1 U504 ( .A1(n513), .A2(n523), .ZN(n351) );
  AND2_X1 U505 ( .A1(n678), .A2(n361), .ZN(n352) );
  XOR2_X1 U506 ( .A(KEYINPUT78), .B(KEYINPUT34), .Z(n353) );
  NAND2_X1 U507 ( .A1(n403), .A2(n678), .ZN(n527) );
  INV_X1 U508 ( .A(n527), .ZN(n454) );
  XOR2_X1 U509 ( .A(n542), .B(KEYINPUT85), .Z(n354) );
  XNOR2_X1 U510 ( .A(KEYINPUT71), .B(KEYINPUT10), .ZN(n355) );
  NOR2_X1 U511 ( .A1(n401), .A2(KEYINPUT41), .ZN(n356) );
  AND2_X1 U512 ( .A1(n496), .A2(n495), .ZN(n357) );
  AND2_X1 U513 ( .A1(n743), .A2(n618), .ZN(n358) );
  NAND2_X1 U514 ( .A1(n644), .A2(n645), .ZN(n790) );
  INV_X1 U515 ( .A(n790), .ZN(n532) );
  AND2_X1 U516 ( .A1(n662), .A2(n390), .ZN(n359) );
  INV_X1 U517 ( .A(G902), .ZN(n426) );
  INV_X1 U518 ( .A(KEYINPUT1), .ZN(n495) );
  AND2_X1 U519 ( .A1(n532), .A2(KEYINPUT40), .ZN(n360) );
  XOR2_X1 U520 ( .A(KEYINPUT117), .B(KEYINPUT36), .Z(n361) );
  XOR2_X1 U521 ( .A(KEYINPUT67), .B(KEYINPUT0), .Z(n362) );
  XOR2_X1 U522 ( .A(KEYINPUT83), .B(KEYINPUT32), .Z(n363) );
  INV_X1 U523 ( .A(KEYINPUT113), .ZN(n533) );
  INV_X1 U524 ( .A(KEYINPUT40), .ZN(n524) );
  INV_X1 U525 ( .A(n353), .ZN(n491) );
  XNOR2_X1 U526 ( .A(G902), .B(KEYINPUT15), .ZN(n685) );
  INV_X1 U527 ( .A(KEYINPUT92), .ZN(n528) );
  INV_X1 U528 ( .A(KEYINPUT2), .ZN(n530) );
  NAND2_X1 U529 ( .A1(n484), .A2(n486), .ZN(n388) );
  NOR2_X1 U530 ( .A1(n679), .A2(n619), .ZN(n405) );
  AND2_X1 U531 ( .A1(n679), .A2(n361), .ZN(n469) );
  NAND2_X1 U532 ( .A1(n407), .A2(n744), .ZN(n679) );
  XNOR2_X1 U533 ( .A(n383), .B(KEYINPUT66), .ZN(n382) );
  XNOR2_X1 U534 ( .A(n507), .B(n610), .ZN(n364) );
  XNOR2_X1 U535 ( .A(n507), .B(n610), .ZN(n629) );
  NOR2_X1 U536 ( .A1(n630), .A2(n663), .ZN(n447) );
  XOR2_X1 U537 ( .A(KEYINPUT72), .B(G131), .Z(n365) );
  XNOR2_X1 U538 ( .A(n447), .B(n533), .ZN(n446) );
  INV_X1 U539 ( .A(n667), .ZN(n459) );
  AND2_X1 U540 ( .A1(n367), .A2(n366), .ZN(n371) );
  INV_X1 U541 ( .A(n795), .ZN(n366) );
  XNOR2_X1 U542 ( .A(n677), .B(KEYINPUT79), .ZN(n367) );
  NAND2_X1 U543 ( .A1(n371), .A2(n369), .ZN(n368) );
  XNOR2_X1 U544 ( .A(n370), .B(KEYINPUT46), .ZN(n369) );
  NAND2_X1 U545 ( .A1(n377), .A2(n375), .ZN(n380) );
  NAND2_X1 U546 ( .A1(n376), .A2(KEYINPUT91), .ZN(n375) );
  INV_X1 U547 ( .A(n509), .ZN(n376) );
  AND2_X1 U548 ( .A1(n505), .A2(n508), .ZN(n379) );
  XNOR2_X1 U549 ( .A(n380), .B(n779), .ZN(G75) );
  XNOR2_X1 U550 ( .A(n381), .B(KEYINPUT95), .ZN(n655) );
  NAND2_X1 U551 ( .A1(n384), .A2(n382), .ZN(n381) );
  XNOR2_X1 U552 ( .A(n385), .B(n481), .ZN(n384) );
  NAND2_X1 U553 ( .A1(n482), .A2(n387), .ZN(n385) );
  XNOR2_X1 U554 ( .A(n559), .B(n386), .ZN(n564) );
  XNOR2_X1 U555 ( .A(n386), .B(n433), .ZN(n722) );
  XNOR2_X2 U556 ( .A(n464), .B(n355), .ZN(n386) );
  NAND2_X1 U557 ( .A1(n811), .A2(KEYINPUT44), .ZN(n387) );
  XNOR2_X2 U558 ( .A(n388), .B(KEYINPUT35), .ZN(n811) );
  NAND2_X1 U559 ( .A1(n389), .A2(n491), .ZN(n487) );
  INV_X1 U560 ( .A(n643), .ZN(n389) );
  AND2_X1 U561 ( .A1(n643), .A2(n353), .ZN(n490) );
  NAND2_X1 U562 ( .A1(n390), .A2(n358), .ZN(n660) );
  NAND2_X1 U563 ( .A1(n676), .A2(n392), .ZN(n677) );
  INV_X1 U564 ( .A(KEYINPUT115), .ZN(n393) );
  OR2_X1 U565 ( .A1(n394), .A2(n522), .ZN(n518) );
  NOR2_X2 U566 ( .A1(n788), .A2(n749), .ZN(n673) );
  XNOR2_X2 U567 ( .A(n395), .B(KEYINPUT84), .ZN(n788) );
  OR2_X2 U568 ( .A1(n668), .A2(n396), .ZN(n395) );
  NAND2_X1 U569 ( .A1(n459), .A2(n671), .ZN(n396) );
  XNOR2_X1 U570 ( .A(n665), .B(n664), .ZN(n668) );
  NAND2_X1 U571 ( .A1(n745), .A2(n398), .ZN(n397) );
  AND2_X1 U572 ( .A1(n401), .A2(KEYINPUT41), .ZN(n398) );
  NAND2_X1 U573 ( .A1(n745), .A2(n744), .ZN(n748) );
  INV_X1 U574 ( .A(n744), .ZN(n402) );
  NOR2_X1 U575 ( .A1(n460), .A2(n772), .ZN(n669) );
  NAND2_X1 U576 ( .A1(n407), .A2(n406), .ZN(n472) );
  NAND2_X1 U577 ( .A1(n623), .A2(n408), .ZN(n443) );
  NAND2_X1 U578 ( .A1(n623), .A2(n409), .ZN(n465) );
  AND2_X1 U579 ( .A1(n626), .A2(n630), .ZN(n409) );
  XNOR2_X2 U580 ( .A(n410), .B(n582), .ZN(n623) );
  NOR2_X1 U581 ( .A1(n680), .A2(n756), .ZN(n626) );
  XNOR2_X1 U582 ( .A(n411), .B(n414), .ZN(n413) );
  XNOR2_X1 U583 ( .A(n421), .B(n419), .ZN(n411) );
  INV_X1 U584 ( .A(n627), .ZN(n474) );
  XNOR2_X2 U585 ( .A(n461), .B(n607), .ZN(n689) );
  INV_X2 U586 ( .A(KEYINPUT64), .ZN(n540) );
  XNOR2_X2 U587 ( .A(KEYINPUT68), .B(G101), .ZN(n595) );
  XNOR2_X1 U588 ( .A(n463), .B(n605), .ZN(n462) );
  XNOR2_X2 U589 ( .A(n412), .B(n354), .ZN(n620) );
  NOR2_X2 U590 ( .A1(n710), .A2(n686), .ZN(n412) );
  XNOR2_X1 U591 ( .A(n413), .B(n805), .ZN(n710) );
  XNOR2_X1 U592 ( .A(n418), .B(n415), .ZN(n421) );
  XNOR2_X1 U593 ( .A(n552), .B(KEYINPUT18), .ZN(n418) );
  NAND2_X1 U594 ( .A1(n724), .A2(G224), .ZN(n420) );
  XNOR2_X2 U595 ( .A(n540), .B(G953), .ZN(n724) );
  NAND2_X1 U596 ( .A1(n697), .A2(G472), .ZN(n430) );
  NAND2_X1 U597 ( .A1(n657), .A2(n744), .ZN(n658) );
  NOR2_X1 U598 ( .A1(n697), .A2(n425), .ZN(n424) );
  NAND2_X1 U599 ( .A1(n431), .A2(n426), .ZN(n566) );
  INV_X1 U600 ( .A(n462), .ZN(n432) );
  INV_X1 U601 ( .A(n637), .ZN(n644) );
  XNOR2_X2 U602 ( .A(n435), .B(KEYINPUT110), .ZN(n793) );
  NAND2_X1 U603 ( .A1(n436), .A2(n637), .ZN(n435) );
  XNOR2_X1 U604 ( .A(n439), .B(n438), .ZN(G33) );
  NAND2_X1 U605 ( .A1(n520), .A2(n519), .ZN(n439) );
  NAND2_X1 U606 ( .A1(n440), .A2(n518), .ZN(n512) );
  INV_X1 U607 ( .A(n483), .ZN(n648) );
  NAND2_X1 U608 ( .A1(n442), .A2(n756), .ZN(n483) );
  XNOR2_X1 U609 ( .A(n443), .B(n624), .ZN(n442) );
  XNOR2_X1 U610 ( .A(n444), .B(n583), .ZN(n445) );
  XNOR2_X1 U611 ( .A(n560), .B(n526), .ZN(n444) );
  XNOR2_X2 U612 ( .A(n721), .B(G146), .ZN(n600) );
  XNOR2_X2 U613 ( .A(n445), .B(n584), .ZN(n721) );
  NAND2_X1 U614 ( .A1(n450), .A2(n474), .ZN(n628) );
  XNOR2_X1 U615 ( .A(n450), .B(G119), .ZN(G21) );
  NAND2_X1 U616 ( .A1(n458), .A2(n456), .ZN(n455) );
  OR2_X1 U617 ( .A1(n668), .A2(n667), .ZN(n460) );
  XNOR2_X1 U618 ( .A(n602), .B(n601), .ZN(n463) );
  XNOR2_X1 U619 ( .A(n552), .B(n622), .ZN(n464) );
  XNOR2_X2 U620 ( .A(n466), .B(KEYINPUT74), .ZN(n663) );
  INV_X1 U621 ( .A(n629), .ZN(n468) );
  INV_X1 U622 ( .A(n657), .ZN(n662) );
  NAND2_X1 U623 ( .A1(n475), .A2(n504), .ZN(n479) );
  NAND2_X1 U624 ( .A1(n349), .A2(n476), .ZN(n475) );
  NAND2_X1 U625 ( .A1(n479), .A2(n477), .ZN(n480) );
  NAND2_X1 U626 ( .A1(n349), .A2(n478), .ZN(n477) );
  AND2_X2 U627 ( .A1(n480), .A2(n505), .ZN(n709) );
  AND2_X1 U628 ( .A1(n483), .A2(n647), .ZN(n482) );
  NAND2_X1 U629 ( .A1(n773), .A2(n491), .ZN(n488) );
  INV_X1 U630 ( .A(n773), .ZN(n489) );
  NAND2_X1 U631 ( .A1(n498), .A2(n496), .ZN(n493) );
  NAND2_X1 U632 ( .A1(n498), .A2(n496), .ZN(n666) );
  NAND2_X1 U633 ( .A1(n733), .A2(n590), .ZN(n500) );
  NAND2_X1 U634 ( .A1(n688), .A2(n349), .ZN(n505) );
  AND2_X2 U635 ( .A1(n731), .A2(G478), .ZN(n694) );
  INV_X1 U636 ( .A(KEYINPUT91), .ZN(n508) );
  XNOR2_X1 U637 ( .A(n511), .B(n510), .ZN(n509) );
  NAND2_X1 U638 ( .A1(n741), .A2(n742), .ZN(n511) );
  NAND2_X1 U639 ( .A1(n512), .A2(n516), .ZN(n520) );
  NAND2_X1 U640 ( .A1(n351), .A2(n518), .ZN(n681) );
  NAND2_X1 U641 ( .A1(n351), .A2(n515), .ZN(n519) );
  AND2_X1 U642 ( .A1(n518), .A2(n360), .ZN(n515) );
  OR2_X1 U643 ( .A1(n661), .A2(n525), .ZN(n522) );
  INV_X1 U644 ( .A(KEYINPUT39), .ZN(n525) );
  INV_X1 U645 ( .A(KEYINPUT73), .ZN(n526) );
  INV_X1 U646 ( .A(KEYINPUT114), .ZN(n531) );
  INV_X1 U647 ( .A(KEYINPUT33), .ZN(n632) );
  INV_X1 U648 ( .A(KEYINPUT28), .ZN(n664) );
  XNOR2_X1 U649 ( .A(n572), .B(n571), .ZN(n576) );
  XNOR2_X1 U650 ( .A(G110), .B(KEYINPUT120), .ZN(n614) );
  XNOR2_X1 U651 ( .A(n535), .B(n534), .ZN(n574) );
  INV_X1 U652 ( .A(n574), .ZN(n536) );
  XNOR2_X1 U653 ( .A(n538), .B(n537), .ZN(n803) );
  XNOR2_X1 U654 ( .A(n595), .B(KEYINPUT76), .ZN(n539) );
  XNOR2_X2 U655 ( .A(G146), .B(G125), .ZN(n552) );
  INV_X1 U656 ( .A(n685), .ZN(n686) );
  NAND2_X1 U657 ( .A1(n541), .A2(n426), .ZN(n543) );
  NAND2_X1 U658 ( .A1(n543), .A2(G210), .ZN(n542) );
  NAND2_X1 U659 ( .A1(n543), .A2(G214), .ZN(n744) );
  NAND2_X1 U660 ( .A1(n620), .A2(n744), .ZN(n545) );
  INV_X1 U661 ( .A(KEYINPUT19), .ZN(n544) );
  XNOR2_X1 U662 ( .A(n545), .B(n544), .ZN(n670) );
  NAND2_X1 U663 ( .A1(G237), .A2(G234), .ZN(n546) );
  XNOR2_X1 U664 ( .A(n546), .B(KEYINPUT14), .ZN(n743) );
  INV_X1 U665 ( .A(G898), .ZN(n806) );
  AND2_X1 U666 ( .A1(n806), .A2(G902), .ZN(n547) );
  NAND2_X1 U667 ( .A1(n547), .A2(G953), .ZN(n548) );
  NAND2_X1 U668 ( .A1(n797), .A2(G952), .ZN(n616) );
  NAND2_X1 U669 ( .A1(n548), .A2(n616), .ZN(n549) );
  NAND2_X1 U670 ( .A1(n743), .A2(n549), .ZN(n550) );
  NOR2_X2 U671 ( .A1(n670), .A2(n550), .ZN(n551) );
  XNOR2_X1 U672 ( .A(n554), .B(n553), .ZN(n558) );
  XNOR2_X1 U673 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U674 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X2 U675 ( .A(KEYINPUT72), .B(G131), .ZN(n560) );
  XOR2_X1 U676 ( .A(n365), .B(KEYINPUT12), .Z(n562) );
  NAND2_X1 U677 ( .A1(G214), .A2(n591), .ZN(n561) );
  XNOR2_X1 U678 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U679 ( .A(KEYINPUT13), .B(G475), .ZN(n565) );
  XNOR2_X1 U680 ( .A(n566), .B(n565), .ZN(n637) );
  NAND2_X1 U681 ( .A1(n724), .A2(G234), .ZN(n567) );
  NAND2_X1 U682 ( .A1(G217), .A2(n606), .ZN(n572) );
  XNOR2_X1 U683 ( .A(n569), .B(G134), .ZN(n584) );
  XNOR2_X1 U684 ( .A(KEYINPUT7), .B(KEYINPUT109), .ZN(n570) );
  XNOR2_X1 U685 ( .A(n584), .B(n570), .ZN(n571) );
  XOR2_X1 U686 ( .A(KEYINPUT108), .B(KEYINPUT9), .Z(n573) );
  XNOR2_X1 U687 ( .A(n574), .B(n573), .ZN(n575) );
  NAND2_X1 U688 ( .A1(n637), .A2(n645), .ZN(n747) );
  XOR2_X1 U689 ( .A(KEYINPUT103), .B(KEYINPUT20), .Z(n578) );
  NAND2_X1 U690 ( .A1(G234), .A2(n685), .ZN(n577) );
  XNOR2_X1 U691 ( .A(n578), .B(n577), .ZN(n608) );
  AND2_X1 U692 ( .A1(n608), .A2(G221), .ZN(n579) );
  XNOR2_X1 U693 ( .A(n579), .B(KEYINPUT21), .ZN(n757) );
  INV_X1 U694 ( .A(n757), .ZN(n580) );
  NOR2_X1 U695 ( .A1(n747), .A2(n580), .ZN(n581) );
  INV_X1 U696 ( .A(KEYINPUT22), .ZN(n582) );
  NAND2_X1 U697 ( .A1(n724), .A2(G227), .ZN(n586) );
  XNOR2_X1 U698 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U699 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U700 ( .A(n600), .B(n589), .ZN(n733) );
  INV_X1 U701 ( .A(G469), .ZN(n590) );
  NAND2_X1 U702 ( .A1(n591), .A2(G210), .ZN(n592) );
  XNOR2_X1 U703 ( .A(n593), .B(n592), .ZN(n594) );
  XOR2_X1 U704 ( .A(n594), .B(KEYINPUT5), .Z(n598) );
  XNOR2_X1 U705 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U706 ( .A(n598), .B(n597), .ZN(n599) );
  XOR2_X1 U707 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n602) );
  XNOR2_X1 U708 ( .A(G137), .B(G110), .ZN(n601) );
  XNOR2_X1 U709 ( .A(G119), .B(G128), .ZN(n604) );
  NAND2_X1 U710 ( .A1(n606), .A2(G221), .ZN(n607) );
  AND2_X1 U711 ( .A1(G217), .A2(n608), .ZN(n609) );
  XNOR2_X1 U712 ( .A(KEYINPUT25), .B(n609), .ZN(n610) );
  BUF_X1 U713 ( .A(n364), .Z(n756) );
  INV_X1 U714 ( .A(n756), .ZN(n611) );
  AND2_X1 U715 ( .A1(n662), .A2(n611), .ZN(n612) );
  AND2_X1 U716 ( .A1(n754), .A2(n612), .ZN(n613) );
  AND2_X1 U717 ( .A1(n623), .A2(n613), .ZN(n627) );
  XOR2_X1 U718 ( .A(n614), .B(n627), .Z(G12) );
  INV_X1 U719 ( .A(n754), .ZN(n619) );
  INV_X1 U720 ( .A(n724), .ZN(n692) );
  NOR2_X1 U721 ( .A1(n426), .A2(G900), .ZN(n615) );
  NAND2_X1 U722 ( .A1(n692), .A2(n615), .ZN(n617) );
  NAND2_X1 U723 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U724 ( .A(n454), .B(n622), .ZN(G42) );
  INV_X1 U725 ( .A(KEYINPUT94), .ZN(n624) );
  XOR2_X1 U726 ( .A(G101), .B(n648), .Z(G3) );
  INV_X1 U727 ( .A(KEYINPUT99), .ZN(n625) );
  XNOR2_X1 U728 ( .A(n754), .B(n625), .ZN(n680) );
  NAND2_X1 U729 ( .A1(n757), .A2(n364), .ZN(n753) );
  INV_X1 U730 ( .A(n630), .ZN(n631) );
  NAND2_X1 U731 ( .A1(n638), .A2(n631), .ZN(n635) );
  XOR2_X1 U732 ( .A(KEYINPUT77), .B(KEYINPUT112), .Z(n633) );
  NOR2_X1 U733 ( .A1(n637), .A2(n645), .ZN(n674) );
  INV_X1 U734 ( .A(n638), .ZN(n639) );
  OR2_X1 U735 ( .A1(n662), .A2(n639), .ZN(n763) );
  INV_X1 U736 ( .A(n763), .ZN(n640) );
  NAND2_X1 U737 ( .A1(n643), .A2(n640), .ZN(n642) );
  INV_X1 U738 ( .A(KEYINPUT31), .ZN(n641) );
  XNOR2_X1 U739 ( .A(n642), .B(n641), .ZN(n792) );
  BUF_X1 U740 ( .A(n657), .Z(n760) );
  NAND2_X1 U741 ( .A1(n643), .A2(n359), .ZN(n781) );
  NAND2_X1 U742 ( .A1(n792), .A2(n781), .ZN(n646) );
  NAND2_X1 U743 ( .A1(n646), .A2(n672), .ZN(n647) );
  OR2_X1 U744 ( .A1(n811), .A2(KEYINPUT44), .ZN(n649) );
  XNOR2_X1 U745 ( .A(n649), .B(KEYINPUT69), .ZN(n653) );
  BUF_X1 U746 ( .A(n650), .Z(n651) );
  XNOR2_X1 U747 ( .A(n651), .B(KEYINPUT97), .ZN(n652) );
  NAND2_X1 U748 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U749 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U750 ( .A(n658), .B(KEYINPUT30), .ZN(n659) );
  INV_X1 U751 ( .A(n661), .ZN(n745) );
  XNOR2_X1 U752 ( .A(n666), .B(KEYINPUT116), .ZN(n667) );
  XNOR2_X1 U753 ( .A(n669), .B(KEYINPUT42), .ZN(n813) );
  INV_X1 U754 ( .A(n670), .ZN(n671) );
  XNOR2_X1 U755 ( .A(n673), .B(KEYINPUT47), .ZN(n676) );
  INV_X1 U756 ( .A(n621), .ZN(n678) );
  NOR2_X1 U757 ( .A1(n681), .A2(n682), .ZN(n683) );
  XNOR2_X1 U758 ( .A(n683), .B(KEYINPUT118), .ZN(n814) );
  INV_X1 U759 ( .A(n814), .ZN(n684) );
  NAND2_X1 U760 ( .A1(n739), .A2(n686), .ZN(n687) );
  INV_X1 U761 ( .A(n739), .ZN(n723) );
  NOR2_X1 U762 ( .A1(n723), .A2(n530), .ZN(n688) );
  BUF_X2 U763 ( .A(n709), .Z(n731) );
  XNOR2_X1 U764 ( .A(n690), .B(n689), .ZN(n693) );
  INV_X1 U765 ( .A(G952), .ZN(n691) );
  NAND2_X1 U766 ( .A1(n692), .A2(n691), .ZN(n717) );
  INV_X1 U767 ( .A(n717), .ZN(n736) );
  NOR2_X1 U768 ( .A1(n693), .A2(n736), .ZN(G66) );
  XNOR2_X1 U769 ( .A(n694), .B(n695), .ZN(n696) );
  NOR2_X1 U770 ( .A1(n696), .A2(n736), .ZN(G63) );
  NAND2_X1 U771 ( .A1(n709), .A2(G472), .ZN(n699) );
  XNOR2_X1 U772 ( .A(n699), .B(n698), .ZN(n700) );
  NAND2_X1 U773 ( .A1(n700), .A2(n717), .ZN(n702) );
  XNOR2_X1 U774 ( .A(KEYINPUT100), .B(KEYINPUT63), .ZN(n701) );
  XNOR2_X1 U775 ( .A(n702), .B(n701), .ZN(G57) );
  NAND2_X1 U776 ( .A1(n709), .A2(G475), .ZN(n705) );
  XOR2_X1 U777 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n703) );
  XNOR2_X1 U778 ( .A(n705), .B(n704), .ZN(n706) );
  NAND2_X1 U779 ( .A1(n706), .A2(n717), .ZN(n708) );
  INV_X1 U780 ( .A(KEYINPUT60), .ZN(n707) );
  XNOR2_X1 U781 ( .A(n708), .B(n707), .ZN(G60) );
  NAND2_X1 U782 ( .A1(n709), .A2(G210), .ZN(n716) );
  BUF_X1 U783 ( .A(n710), .Z(n711) );
  XNOR2_X1 U784 ( .A(KEYINPUT123), .B(KEYINPUT54), .ZN(n713) );
  XNOR2_X1 U785 ( .A(KEYINPUT55), .B(KEYINPUT87), .ZN(n712) );
  XNOR2_X1 U786 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U787 ( .A(n716), .B(n715), .ZN(n718) );
  NAND2_X1 U788 ( .A1(n718), .A2(n717), .ZN(n720) );
  XNOR2_X1 U789 ( .A(KEYINPUT93), .B(KEYINPUT56), .ZN(n719) );
  XNOR2_X1 U790 ( .A(n720), .B(n719), .ZN(G51) );
  XOR2_X1 U791 ( .A(n722), .B(n721), .Z(n726) );
  XNOR2_X1 U792 ( .A(n723), .B(n726), .ZN(n725) );
  NAND2_X1 U793 ( .A1(n725), .A2(n724), .ZN(n730) );
  XNOR2_X1 U794 ( .A(G227), .B(n726), .ZN(n727) );
  NAND2_X1 U795 ( .A1(n727), .A2(G900), .ZN(n728) );
  NAND2_X1 U796 ( .A1(n728), .A2(G953), .ZN(n729) );
  NAND2_X1 U797 ( .A1(n730), .A2(n729), .ZN(G72) );
  NAND2_X1 U798 ( .A1(n731), .A2(G469), .ZN(n735) );
  XOR2_X1 U799 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n732) );
  XNOR2_X1 U800 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U801 ( .A(n735), .B(n734), .ZN(n737) );
  NOR2_X1 U802 ( .A1(n737), .A2(n736), .ZN(G54) );
  NAND2_X1 U803 ( .A1(n738), .A2(n530), .ZN(n742) );
  XNOR2_X1 U804 ( .A(n740), .B(KEYINPUT89), .ZN(n741) );
  NAND2_X1 U805 ( .A1(G952), .A2(n743), .ZN(n771) );
  NOR2_X1 U806 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U807 ( .A1(n747), .A2(n746), .ZN(n751) );
  NOR2_X1 U808 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U809 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U810 ( .A1(n773), .A2(n752), .ZN(n768) );
  NAND2_X1 U811 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U812 ( .A(n755), .B(KEYINPUT50), .ZN(n762) );
  NOR2_X1 U813 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U814 ( .A(KEYINPUT49), .B(n758), .Z(n759) );
  NOR2_X1 U815 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U816 ( .A1(n762), .A2(n761), .ZN(n764) );
  NAND2_X1 U817 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U818 ( .A(KEYINPUT51), .B(n765), .ZN(n766) );
  NOR2_X1 U819 ( .A1(n766), .A2(n772), .ZN(n767) );
  NOR2_X1 U820 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U821 ( .A(n769), .B(KEYINPUT52), .ZN(n770) );
  NOR2_X1 U822 ( .A1(n771), .A2(n770), .ZN(n775) );
  NOR2_X1 U823 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U824 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U825 ( .A(n776), .B(KEYINPUT121), .ZN(n777) );
  NOR2_X1 U826 ( .A1(n777), .A2(G953), .ZN(n778) );
  XOR2_X1 U827 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n779) );
  NOR2_X1 U828 ( .A1(n790), .A2(n781), .ZN(n780) );
  XOR2_X1 U829 ( .A(G104), .B(n780), .Z(G6) );
  NOR2_X1 U830 ( .A1(n781), .A2(n793), .ZN(n785) );
  XOR2_X1 U831 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n783) );
  XNOR2_X1 U832 ( .A(G107), .B(KEYINPUT119), .ZN(n782) );
  XNOR2_X1 U833 ( .A(n783), .B(n782), .ZN(n784) );
  XNOR2_X1 U834 ( .A(n785), .B(n784), .ZN(G9) );
  XNOR2_X1 U835 ( .A(G128), .B(KEYINPUT29), .ZN(n787) );
  NOR2_X1 U836 ( .A1(n793), .A2(n788), .ZN(n786) );
  XNOR2_X1 U837 ( .A(n787), .B(n786), .ZN(G30) );
  NOR2_X1 U838 ( .A1(n788), .A2(n790), .ZN(n789) );
  XOR2_X1 U839 ( .A(G146), .B(n789), .Z(G48) );
  NOR2_X1 U840 ( .A1(n790), .A2(n792), .ZN(n791) );
  XOR2_X1 U841 ( .A(G113), .B(n791), .Z(G15) );
  NOR2_X1 U842 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U843 ( .A(G116), .B(n794), .Z(G18) );
  XNOR2_X1 U844 ( .A(G125), .B(n795), .ZN(n796) );
  XNOR2_X1 U845 ( .A(n796), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U846 ( .A1(n349), .A2(n797), .ZN(n801) );
  NAND2_X1 U847 ( .A1(G953), .A2(G224), .ZN(n798) );
  XNOR2_X1 U848 ( .A(KEYINPUT61), .B(n798), .ZN(n799) );
  NAND2_X1 U849 ( .A1(n799), .A2(G898), .ZN(n800) );
  NAND2_X1 U850 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U851 ( .A(n802), .B(KEYINPUT125), .ZN(n810) );
  XOR2_X1 U852 ( .A(n803), .B(G101), .Z(n804) );
  XNOR2_X1 U853 ( .A(n805), .B(n804), .ZN(n808) );
  NAND2_X1 U854 ( .A1(n806), .A2(G953), .ZN(n807) );
  AND2_X1 U855 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U856 ( .A(n810), .B(n809), .Z(G69) );
  XNOR2_X1 U857 ( .A(G122), .B(n811), .ZN(n812) );
  XNOR2_X1 U858 ( .A(n812), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U859 ( .A(G137), .B(n813), .Z(G39) );
  XOR2_X1 U860 ( .A(G134), .B(n814), .Z(G36) );
endmodule

