//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1308, new_n1309, new_n1310;
  NOR4_X1   g0000(.A1(KEYINPUT64), .A2(G50), .A3(G58), .A4(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(G50), .ZN(new_n204));
  AOI21_X1  g0004(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NOR3_X1   g0005(.A1(new_n201), .A2(new_n205), .A3(G77), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G77), .A2(G244), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G68), .A2(G238), .ZN(new_n213));
  AND3_X1   g0013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n209), .A2(new_n210), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT1), .Z(new_n218));
  NOR2_X1   g0018(.A1(new_n216), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT0), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G20), .ZN(new_n224));
  INV_X1    g0024(.A(new_n203), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n218), .B(new_n221), .C1(new_n224), .C2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT66), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G264), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(G270), .Z(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  INV_X1    g0036(.A(G107), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(G97), .ZN(new_n238));
  INV_X1    g0038(.A(G97), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G107), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G87), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(G200), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G223), .A3(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(G222), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G77), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n260), .B(new_n262), .C1(new_n263), .C2(new_n259), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n223), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n254), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n266), .A2(new_n252), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G226), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n250), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n268), .A2(G190), .A3(new_n270), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT68), .ZN(new_n273));
  INV_X1    g0073(.A(G20), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G33), .ZN(new_n275));
  AND2_X1   g0075(.A1(KEYINPUT8), .A2(G58), .ZN(new_n276));
  NOR2_X1   g0076(.A1(KEYINPUT8), .A2(G58), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G150), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n273), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(G20), .B1(new_n201), .B2(new_n205), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  OAI211_X1 g0084(.A(KEYINPUT68), .B(new_n280), .C1(new_n284), .C2(new_n275), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(KEYINPUT67), .B1(new_n216), .B2(new_n256), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT67), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n288), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n287), .A2(new_n222), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G50), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n290), .B1(new_n251), .B2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G50), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n291), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT9), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n293), .B1(new_n286), .B2(new_n290), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(new_n300), .A3(new_n296), .ZN(new_n301));
  AOI211_X1 g0101(.A(new_n271), .B(new_n272), .C1(new_n298), .C2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  AOI21_X1  g0103(.A(KEYINPUT72), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n271), .B1(new_n298), .B2(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n264), .A2(new_n267), .ZN(new_n306));
  INV_X1    g0106(.A(new_n254), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n306), .A2(new_n307), .A3(new_n270), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G190), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n305), .A2(KEYINPUT72), .A3(new_n303), .A4(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n271), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n299), .A2(new_n300), .A3(new_n296), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n300), .B1(new_n299), .B2(new_n296), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n309), .B(new_n312), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT73), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT10), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n316), .B1(new_n315), .B2(KEYINPUT10), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n304), .A2(new_n311), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(KEYINPUT3), .A2(G33), .ZN(new_n321));
  OAI211_X1 g0121(.A(G226), .B(new_n261), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(G232), .B(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G33), .A2(G97), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n254), .B1(new_n325), .B2(new_n267), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n269), .A2(G238), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT13), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT13), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n326), .A2(new_n330), .A3(new_n327), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(G190), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n325), .A2(new_n267), .ZN(new_n333));
  AND4_X1   g0133(.A1(new_n330), .A2(new_n333), .A3(new_n327), .A4(new_n307), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n330), .B1(new_n326), .B2(new_n327), .ZN(new_n335));
  OAI21_X1  g0135(.A(G200), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n295), .A2(G68), .ZN(new_n337));
  INV_X1    g0137(.A(G68), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G20), .ZN(new_n339));
  INV_X1    g0139(.A(new_n279), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n339), .B1(new_n275), .B2(new_n263), .C1(new_n340), .C2(new_n204), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n290), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT11), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(KEYINPUT11), .A3(new_n290), .ZN(new_n345));
  INV_X1    g0145(.A(new_n292), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n338), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT12), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n337), .A2(new_n344), .A3(new_n345), .A4(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AND3_X1   g0150(.A1(new_n332), .A2(new_n336), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(G169), .B1(new_n334), .B2(new_n335), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT14), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n329), .A2(G179), .A3(new_n331), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT14), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n355), .B(G169), .C1(new_n334), .C2(new_n335), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n351), .B1(new_n357), .B2(new_n349), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n319), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT16), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G58), .A2(G68), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n274), .B1(new_n225), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n257), .A2(new_n274), .A3(new_n258), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT7), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n320), .A2(new_n321), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(KEYINPUT7), .A3(new_n274), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n362), .B1(new_n368), .B2(G68), .ZN(new_n369));
  INV_X1    g0169(.A(G159), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n340), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n360), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n338), .B1(new_n365), .B2(new_n367), .ZN(new_n374));
  NOR4_X1   g0174(.A1(new_n374), .A2(KEYINPUT16), .A3(new_n371), .A4(new_n362), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n290), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n276), .A2(new_n277), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(new_n292), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n251), .A2(G20), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  XOR2_X1   g0181(.A(new_n381), .B(KEYINPUT74), .Z(new_n382));
  NOR3_X1   g0182(.A1(new_n382), .A2(new_n290), .A3(new_n346), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n376), .A2(new_n379), .A3(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(G226), .B(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n386));
  OAI211_X1 g0186(.A(G223), .B(new_n261), .C1(new_n320), .C2(new_n321), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT75), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n256), .B2(new_n242), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n388), .A2(new_n256), .A3(new_n242), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n267), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n392), .A2(new_n307), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n269), .A2(G232), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G169), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G179), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(new_n398), .A3(new_n394), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n385), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT18), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n385), .A2(KEYINPUT18), .A3(new_n397), .A4(new_n399), .ZN(new_n403));
  INV_X1    g0203(.A(new_n290), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT7), .B1(new_n366), .B2(new_n274), .ZN(new_n405));
  NOR4_X1   g0205(.A1(new_n320), .A2(new_n321), .A3(new_n364), .A4(G20), .ZN(new_n406));
  OAI21_X1  g0206(.A(G68), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n362), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(new_n372), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT16), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n407), .A2(new_n360), .A3(new_n372), .A4(new_n408), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n404), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n412), .A2(new_n378), .A3(new_n383), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT17), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n395), .A2(G200), .ZN(new_n415));
  AND4_X1   g0215(.A1(G190), .A2(new_n392), .A3(new_n394), .A4(new_n307), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n413), .A2(new_n414), .A3(new_n415), .A4(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n376), .A2(new_n384), .A3(new_n379), .A4(new_n417), .ZN(new_n419));
  INV_X1    g0219(.A(new_n415), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT17), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n402), .A2(new_n403), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n377), .B(KEYINPUT70), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n279), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT15), .B(G87), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n425), .B(KEYINPUT71), .ZN(new_n426));
  OAI221_X1 g0226(.A(new_n424), .B1(new_n274), .B2(new_n263), .C1(new_n275), .C2(new_n426), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n427), .A2(new_n290), .B1(new_n263), .B2(new_n346), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n295), .A2(G77), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n259), .A2(G238), .A3(G1698), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n259), .A2(G232), .A3(new_n261), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n431), .B(new_n432), .C1(new_n237), .C2(new_n259), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n267), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n269), .A2(G244), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n307), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n396), .ZN(new_n437));
  INV_X1    g0237(.A(new_n436), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n398), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n430), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n422), .A2(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n308), .A2(G169), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n308), .A2(new_n398), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n297), .A3(new_n443), .ZN(new_n444));
  XOR2_X1   g0244(.A(new_n444), .B(KEYINPUT69), .Z(new_n445));
  NAND2_X1  g0245(.A1(new_n438), .A2(G190), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n436), .A2(G200), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n428), .A2(new_n446), .A3(new_n447), .A4(new_n429), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n359), .A2(new_n441), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT5), .B(G41), .ZN(new_n451));
  INV_X1    g0251(.A(G45), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(G1), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n451), .A2(new_n453), .B1(new_n223), .B2(new_n265), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n251), .A2(G45), .ZN(new_n455));
  OR2_X1    g0255(.A1(KEYINPUT5), .A2(G41), .ZN(new_n456));
  NAND2_X1  g0256(.A1(KEYINPUT5), .A2(G41), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n454), .A2(G270), .B1(G274), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(G257), .B(new_n261), .C1(new_n320), .C2(new_n321), .ZN(new_n460));
  OAI211_X1 g0260(.A(G264), .B(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n257), .A2(G303), .A3(new_n258), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n267), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT82), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT82), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n459), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G200), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n244), .A2(G20), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G283), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n472), .B(new_n274), .C1(G33), .C2(new_n239), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n290), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT20), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n290), .A2(KEYINPUT20), .A3(new_n471), .A4(new_n473), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n256), .A2(G1), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n290), .A2(new_n346), .A3(new_n478), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n476), .A2(new_n477), .B1(G116), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n346), .A2(new_n244), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G190), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n470), .B(new_n483), .C1(new_n484), .C2(new_n469), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n469), .A2(G169), .A3(new_n482), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT21), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n459), .A2(G179), .A3(new_n464), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n469), .A2(new_n482), .A3(KEYINPUT21), .A4(G169), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n485), .A2(new_n488), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G116), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(G20), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n274), .B(G87), .C1(new_n320), .C2(new_n321), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT22), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT22), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n259), .A2(new_n498), .A3(new_n274), .A4(G87), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT24), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n274), .A2(G107), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n502), .B(KEYINPUT23), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n501), .B1(new_n500), .B2(new_n503), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n290), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n479), .A2(G107), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n292), .A2(G107), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n508), .B(KEYINPUT25), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(G257), .B(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n511));
  OAI211_X1 g0311(.A(G250), .B(new_n261), .C1(new_n320), .C2(new_n321), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G294), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(new_n267), .B1(new_n454), .B2(G264), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n458), .A2(G274), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n250), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n516), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n484), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n510), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT83), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n515), .A2(G179), .A3(new_n516), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n396), .B1(new_n515), .B2(new_n516), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n518), .A2(G169), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n515), .A2(G179), .A3(new_n516), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(KEYINPUT83), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT84), .B1(new_n528), .B2(new_n510), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(KEYINPUT84), .A3(new_n510), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n520), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(G244), .B(new_n261), .C1(new_n320), .C2(new_n321), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n261), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n259), .A2(G250), .A3(G1698), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n472), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n267), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT77), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n451), .A2(new_n453), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(new_n266), .A3(G257), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n516), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n535), .A2(new_n536), .A3(new_n472), .A4(new_n538), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT77), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(new_n547), .A3(new_n267), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n541), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n544), .B1(new_n267), .B2(new_n546), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n549), .A2(G200), .B1(G190), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(G107), .B1(new_n405), .B2(new_n406), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT76), .B1(new_n279), .B2(G77), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT6), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n238), .A2(new_n240), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n237), .A2(KEYINPUT6), .A3(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n553), .B1(new_n557), .B2(G20), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n279), .A2(KEYINPUT76), .A3(G77), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n552), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n290), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n346), .A2(new_n239), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n479), .A2(G97), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n551), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT78), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n540), .A2(new_n545), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n396), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n541), .A2(new_n398), .A3(new_n545), .A4(new_n548), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n560), .A2(new_n290), .B1(G97), .B2(new_n479), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(KEYINPUT78), .A3(new_n562), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n568), .A2(new_n570), .A3(new_n571), .A4(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(G33), .A2(G41), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n455), .B(G250), .C1(new_n575), .C2(new_n222), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n453), .A2(G274), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(G244), .B(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n579));
  OAI211_X1 g0379(.A(G238), .B(new_n261), .C1(new_n320), .C2(new_n321), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n580), .A3(new_n494), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n578), .B1(new_n581), .B2(new_n267), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n582), .A2(G169), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n398), .ZN(new_n585));
  AND2_X1   g0385(.A1(KEYINPUT79), .A2(G87), .ZN(new_n586));
  NOR2_X1   g0386(.A1(KEYINPUT79), .A2(G87), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n239), .B(new_n237), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n324), .A2(new_n274), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(KEYINPUT19), .A3(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n274), .B(G68), .C1(new_n320), .C2(new_n321), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT80), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n259), .A2(KEYINPUT80), .A3(new_n274), .A4(G68), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT19), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n275), .B2(new_n239), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n590), .A2(new_n593), .A3(new_n594), .A4(new_n596), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n597), .A2(new_n290), .B1(new_n346), .B2(new_n426), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT81), .ZN(new_n599));
  INV_X1    g0399(.A(new_n426), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n479), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n599), .B1(new_n598), .B2(new_n601), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n584), .B(new_n585), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n582), .A2(new_n250), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(G190), .B2(new_n582), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n479), .A2(G87), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n598), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n566), .A2(new_n574), .A3(new_n604), .A4(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n450), .A2(new_n493), .A3(new_n532), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n611), .B(KEYINPUT85), .ZN(G372));
  NAND2_X1  g0412(.A1(new_n315), .A2(KEYINPUT10), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT73), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT10), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT72), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n315), .B2(KEYINPUT10), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n614), .A2(new_n615), .B1(new_n617), .B2(new_n310), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n418), .A2(new_n421), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n357), .A2(new_n349), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n440), .ZN(new_n621));
  INV_X1    g0421(.A(new_n351), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n619), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n402), .A2(new_n403), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n618), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT86), .ZN(new_n626));
  INV_X1    g0426(.A(new_n445), .ZN(new_n627));
  OR3_X1    g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n625), .B2(new_n627), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(KEYINPUT78), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT78), .B1(new_n572), .B2(new_n562), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n571), .A2(new_n570), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n633), .A2(new_n634), .B1(new_n565), .B2(new_n551), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n525), .A2(new_n526), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n510), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n637), .A2(new_n488), .A3(new_n490), .A4(new_n491), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n604), .A2(new_n608), .ZN(new_n639));
  OR3_X1    g0439(.A1(new_n510), .A2(new_n517), .A3(new_n519), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n635), .A2(new_n638), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n604), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n633), .A2(new_n604), .A3(new_n608), .A4(new_n634), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(KEYINPUT26), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n604), .A2(new_n608), .A3(new_n634), .A4(new_n564), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n645), .A2(KEYINPUT26), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n641), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n450), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n630), .A2(new_n648), .ZN(G369));
  NAND3_X1  g0449(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n650));
  INV_X1    g0450(.A(G13), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(G20), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n251), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n650), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n532), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n637), .B2(new_n658), .ZN(new_n662));
  XOR2_X1   g0462(.A(new_n662), .B(KEYINPUT87), .Z(new_n663));
  NOR2_X1   g0463(.A1(new_n483), .A2(new_n659), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n650), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n492), .B2(new_n664), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n528), .A2(new_n510), .A3(new_n658), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n528), .A2(KEYINPUT84), .A3(new_n510), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n640), .B1(new_n669), .B2(new_n529), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n510), .A2(new_n658), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n663), .A2(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n219), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G1), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n588), .A2(G116), .ZN(new_n679));
  OAI22_X1  g0479(.A1(new_n678), .A2(new_n679), .B1(new_n226), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  NOR4_X1   g0481(.A1(new_n670), .A2(new_n609), .A3(new_n492), .A4(new_n658), .ZN(new_n682));
  AOI21_X1  g0482(.A(G179), .B1(new_n466), .B2(new_n468), .ZN(new_n683));
  INV_X1    g0483(.A(new_n582), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n683), .A2(new_n518), .A3(new_n549), .A4(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT30), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT88), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n515), .A2(new_n582), .A3(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n489), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n687), .B1(new_n515), .B2(new_n582), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(new_n569), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n686), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n489), .A2(new_n688), .ZN(new_n693));
  NOR4_X1   g0493(.A1(new_n693), .A2(new_n569), .A3(new_n690), .A4(KEYINPUT30), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n685), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(KEYINPUT89), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n515), .A2(new_n582), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT88), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n489), .A3(new_n550), .A4(new_n688), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT30), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n689), .A2(new_n691), .A3(new_n686), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT89), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(new_n685), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n698), .A2(new_n658), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT31), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n697), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n682), .B1(new_n709), .B2(KEYINPUT90), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n704), .A2(new_n705), .A3(new_n685), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n705), .B1(new_n704), .B2(new_n685), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n711), .A2(new_n712), .A3(new_n659), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n696), .B1(new_n713), .B2(KEYINPUT31), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT90), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n710), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G330), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n647), .A2(new_n659), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT29), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n643), .A2(KEYINPUT26), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n642), .B1(new_n645), .B2(KEYINPUT26), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n650), .B1(new_n530), .B2(new_n531), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n635), .A2(new_n640), .A3(new_n639), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n723), .B(new_n724), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n722), .B1(new_n727), .B2(new_n659), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n719), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n681), .B1(new_n730), .B2(G1), .ZN(G364));
  NOR2_X1   g0531(.A1(new_n666), .A2(G330), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n251), .B1(new_n652), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n676), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n667), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT91), .Z(new_n737));
  NAND2_X1  g0537(.A1(new_n248), .A2(G45), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n675), .A2(new_n259), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n738), .B(new_n739), .C1(G45), .C2(new_n226), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n259), .A2(G355), .A3(new_n219), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n740), .B(new_n741), .C1(G116), .C2(new_n219), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n222), .B1(G20), .B2(new_n396), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n274), .A2(G179), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(G190), .A3(G200), .ZN(new_n750));
  OR3_X1    g0550(.A1(new_n750), .A2(new_n587), .A3(new_n586), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n749), .A2(new_n484), .A3(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G190), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(KEYINPUT92), .B(G159), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n751), .B1(new_n237), .B2(new_n752), .C1(KEYINPUT32), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n274), .A2(new_n398), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(G190), .A3(new_n250), .ZN(new_n760));
  INV_X1    g0560(.A(G58), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n259), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n759), .A2(new_n753), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n762), .B1(G77), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n759), .A2(new_n484), .A3(G200), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n757), .A2(KEYINPUT32), .B1(new_n767), .B2(G68), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n484), .A2(G179), .A3(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n274), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n765), .B(new_n768), .C1(new_n239), .C2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n759), .A2(G190), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n758), .B(new_n771), .C1(G50), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(G326), .ZN(new_n775));
  INV_X1    g0575(.A(G294), .ZN(new_n776));
  XOR2_X1   g0576(.A(KEYINPUT33), .B(G317), .Z(new_n777));
  OAI221_X1 g0577(.A(new_n775), .B1(new_n776), .B2(new_n770), .C1(new_n766), .C2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G322), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n760), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G283), .ZN(new_n781));
  INV_X1    g0581(.A(G303), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n781), .A2(new_n752), .B1(new_n750), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G329), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n366), .B1(new_n754), .B2(new_n784), .C1(new_n785), .C2(new_n763), .ZN(new_n786));
  NOR4_X1   g0586(.A1(new_n778), .A2(new_n780), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n746), .B1(new_n774), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n748), .A2(new_n735), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT93), .ZN(new_n790));
  INV_X1    g0590(.A(new_n745), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n790), .B1(new_n666), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n737), .A2(new_n792), .ZN(G396));
  OR2_X1    g0593(.A1(new_n440), .A2(new_n658), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n430), .A2(new_n658), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n448), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n440), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n720), .B(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n718), .B(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n735), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n773), .A2(G137), .B1(new_n764), .B2(new_n756), .ZN(new_n803));
  INV_X1    g0603(.A(G150), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n804), .B2(new_n766), .ZN(new_n805));
  INV_X1    g0605(.A(new_n760), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(G143), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT95), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT34), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n752), .A2(new_n338), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n259), .B1(new_n770), .B2(new_n761), .ZN(new_n811));
  INV_X1    g0611(.A(new_n750), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n810), .B(new_n811), .C1(G50), .C2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(G132), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n809), .B(new_n813), .C1(new_n814), .C2(new_n754), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n366), .B1(new_n763), .B2(new_n244), .C1(new_n776), .C2(new_n760), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n752), .A2(new_n242), .ZN(new_n817));
  INV_X1    g0617(.A(new_n770), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(G97), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n782), .B2(new_n772), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n816), .B(new_n820), .C1(G311), .C2(new_n755), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n767), .A2(KEYINPUT94), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n767), .A2(KEYINPUT94), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n821), .B1(new_n237), .B2(new_n750), .C1(new_n781), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n815), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n746), .A2(new_n743), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n826), .A2(new_n746), .B1(new_n263), .B2(new_n827), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n828), .B(new_n735), .C1(new_n744), .C2(new_n798), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n802), .A2(new_n829), .ZN(G384));
  OAI211_X1 g0630(.A(G20), .B(new_n223), .C1(new_n557), .C2(KEYINPUT35), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n244), .B(new_n831), .C1(KEYINPUT35), .C2(new_n557), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT36), .Z(new_n833));
  NAND2_X1  g0633(.A1(new_n361), .A2(G77), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n226), .A2(new_n834), .B1(G50), .B2(new_n338), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n835), .A2(G1), .A3(new_n651), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT96), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT101), .ZN(new_n839));
  NOR4_X1   g0639(.A1(new_n412), .A2(new_n378), .A3(new_n383), .A4(new_n416), .ZN(new_n840));
  INV_X1    g0640(.A(new_n656), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n840), .A2(new_n415), .B1(new_n385), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT100), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n842), .B(new_n400), .C1(new_n843), .C2(KEYINPUT37), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n410), .A2(new_n411), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n383), .B1(new_n845), .B2(new_n290), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n846), .A2(new_n379), .A3(new_n415), .A4(new_n417), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n385), .A2(new_n841), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n400), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n847), .A2(new_n848), .A3(new_n843), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT37), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n844), .B(new_n852), .C1(new_n422), .C2(new_n848), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n839), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n844), .A2(new_n852), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n624), .A2(new_n619), .ZN(new_n857));
  INV_X1    g0657(.A(new_n848), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n856), .A2(KEYINPUT101), .A3(KEYINPUT38), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n853), .A2(new_n854), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n855), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT102), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n619), .A2(new_n864), .B1(new_n402), .B2(new_n403), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n418), .A2(new_n421), .A3(KEYINPUT102), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n848), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n844), .A2(new_n852), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n854), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT39), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n856), .A2(KEYINPUT38), .A3(new_n859), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n863), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n620), .A2(new_n658), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n624), .A2(new_n841), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n620), .A2(new_n659), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n349), .A2(new_n658), .ZN(new_n880));
  AND4_X1   g0680(.A1(KEYINPUT97), .A2(new_n620), .A3(new_n622), .A4(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT97), .B1(new_n358), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT98), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n620), .A2(new_n622), .A3(new_n880), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT97), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n358), .A2(KEYINPUT97), .A3(new_n880), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT98), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(new_n890), .A3(new_n879), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n884), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n647), .A2(new_n798), .A3(new_n659), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n794), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT99), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n884), .A2(new_n891), .B1(new_n893), .B2(new_n794), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT99), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n897), .A2(new_n899), .A3(new_n862), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n875), .A2(new_n877), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n450), .B1(new_n721), .B2(new_n728), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n630), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n901), .B(new_n903), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n532), .A2(new_n610), .A3(new_n493), .A4(new_n659), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n707), .A2(new_n708), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n658), .A4(new_n706), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n794), .A2(new_n797), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n884), .B2(new_n891), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n862), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n890), .B1(new_n889), .B2(new_n879), .ZN(new_n913));
  AOI211_X1 g0713(.A(KEYINPUT98), .B(new_n878), .C1(new_n887), .C2(new_n888), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n798), .B(new_n908), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n912), .B1(new_n869), .B2(new_n871), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n911), .A2(new_n912), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n450), .A2(new_n908), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n918), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(G330), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n904), .A2(new_n921), .B1(new_n251), .B2(new_n652), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT103), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n904), .A2(new_n921), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n838), .B1(new_n923), .B2(new_n924), .ZN(G367));
  AOI21_X1  g0725(.A(new_n635), .B1(new_n564), .B2(new_n658), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n634), .A2(new_n565), .A3(new_n659), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OR4_X1    g0729(.A1(KEYINPUT107), .A2(new_n663), .A3(KEYINPUT44), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n663), .A2(new_n929), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT45), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n663), .A2(KEYINPUT45), .A3(new_n929), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n663), .B2(new_n929), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n672), .A2(new_n660), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n667), .B1(new_n939), .B2(new_n661), .ZN(new_n940));
  INV_X1    g0740(.A(new_n673), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n729), .B(new_n719), .C1(new_n938), .C2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n676), .B(KEYINPUT41), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n733), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OR3_X1    g0746(.A1(new_n928), .A2(KEYINPUT42), .A3(new_n661), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n530), .A2(new_n531), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n574), .B1(new_n928), .B2(new_n948), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n947), .A2(KEYINPUT105), .B1(new_n659), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT42), .B1(new_n928), .B2(new_n661), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n950), .B(new_n951), .C1(KEYINPUT105), .C2(new_n947), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n952), .A2(KEYINPUT106), .ZN(new_n953));
  INV_X1    g0753(.A(new_n639), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n659), .B1(new_n598), .B2(new_n607), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT104), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n642), .A2(new_n955), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(KEYINPUT104), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT43), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n952), .A2(KEYINPUT106), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n953), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n673), .A2(new_n928), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n953), .B2(new_n962), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n965), .B1(new_n964), .B2(new_n967), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n946), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n739), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n747), .B1(new_n219), .B2(new_n426), .C1(new_n235), .C2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n824), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n756), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n752), .A2(new_n263), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n770), .A2(new_n338), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n975), .B(new_n976), .C1(G58), .C2(new_n812), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n773), .A2(G143), .ZN(new_n978));
  INV_X1    g0778(.A(G137), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n259), .B1(new_n754), .B2(new_n979), .C1(new_n760), .C2(new_n804), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(G50), .B2(new_n764), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n974), .A2(new_n977), .A3(new_n978), .A4(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n750), .A2(new_n244), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT46), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n772), .A2(new_n785), .B1(new_n752), .B2(new_n239), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n366), .B1(new_n760), .B2(new_n782), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n770), .A2(new_n237), .B1(new_n763), .B2(new_n781), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT108), .Z(new_n989));
  OAI211_X1 g0789(.A(new_n987), .B(new_n989), .C1(new_n776), .C2(new_n824), .ZN(new_n990));
  INV_X1    g0790(.A(G317), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n754), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n982), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT47), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n801), .B1(new_n994), .B2(new_n746), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n972), .B(new_n995), .C1(new_n960), .C2(new_n791), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n970), .A2(new_n996), .ZN(G387));
  OAI22_X1  g0797(.A1(new_n824), .A2(new_n785), .B1(new_n779), .B2(new_n772), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT112), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n782), .B2(new_n763), .C1(new_n991), .C2(new_n760), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT48), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n781), .B2(new_n770), .C1(new_n776), .C2(new_n750), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT49), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n752), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n259), .B1(new_n1006), .B2(G116), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1004), .B(new_n1008), .C1(G326), .C2(new_n755), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n750), .A2(new_n263), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G97), .B2(new_n1006), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n370), .B2(new_n772), .C1(new_n284), .C2(new_n766), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n600), .A2(new_n818), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n366), .B1(new_n806), .B2(G50), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(new_n804), .C2(new_n754), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1012), .B(new_n1015), .C1(G68), .C2(new_n764), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT111), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n746), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n672), .A2(new_n791), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n232), .A2(G45), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT109), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n423), .A2(new_n204), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1022), .A2(KEYINPUT50), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(KEYINPUT50), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n679), .B1(G68), .B2(G77), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1024), .A2(new_n452), .A3(new_n1025), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1021), .B(new_n739), .C1(new_n1023), .C2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n679), .A2(new_n219), .A3(new_n259), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(G107), .C2(new_n219), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT110), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(KEYINPUT110), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n747), .A3(new_n1031), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1018), .A2(new_n735), .A3(new_n1019), .A4(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n942), .A2(new_n734), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n730), .A2(new_n942), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n730), .A2(new_n942), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1035), .A2(new_n676), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1033), .A2(new_n1034), .A3(new_n1037), .ZN(G393));
  XNOR2_X1  g0838(.A(new_n938), .B(new_n941), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n677), .B1(new_n1039), .B2(new_n1036), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n938), .A2(new_n730), .A3(new_n942), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1039), .A2(new_n733), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n928), .A2(new_n745), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n973), .A2(G303), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n812), .A2(G283), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n760), .A2(new_n785), .B1(new_n772), .B2(new_n991), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT52), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n366), .B1(new_n754), .B2(new_n779), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n770), .A2(new_n244), .B1(new_n752), .B2(new_n237), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G294), .C2(new_n764), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .A4(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n366), .B1(new_n755), .B2(G143), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n338), .B2(new_n750), .C1(new_n242), .C2(new_n752), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT114), .Z(new_n1055));
  OAI22_X1  g0855(.A1(new_n760), .A2(new_n370), .B1(new_n772), .B2(new_n804), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT51), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n973), .A2(G50), .B1(new_n423), .B2(new_n764), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n770), .A2(new_n263), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1052), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n746), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n747), .B1(new_n239), .B2(new_n219), .C1(new_n245), .C2(new_n971), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n735), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT113), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1044), .A2(new_n1062), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1042), .A2(new_n1043), .A3(new_n1066), .ZN(G390));
  INV_X1    g0867(.A(KEYINPUT117), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n798), .A2(G330), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n892), .B1(new_n717), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n913), .A2(new_n914), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n908), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n894), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n906), .A2(KEYINPUT90), .A3(new_n696), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n905), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n709), .A2(KEYINPUT90), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n892), .B(new_n1069), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n727), .A2(new_n659), .A3(new_n797), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1079), .A2(new_n794), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1074), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n450), .A2(G330), .A3(new_n908), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n630), .A2(new_n902), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT116), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT116), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1088), .B(new_n1085), .C1(new_n1074), .C2(new_n1082), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT115), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n898), .B2(new_n874), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n874), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n895), .A2(KEYINPUT115), .A3(new_n1092), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1091), .A2(new_n1093), .A3(new_n863), .A4(new_n872), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n874), .B1(new_n869), .B2(new_n871), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n1071), .B2(new_n1080), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1078), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1073), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n1087), .A2(new_n1089), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n894), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1069), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n1071), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n892), .A2(new_n908), .A3(new_n1069), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1101), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1086), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n1088), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1096), .B1(new_n1109), .B2(new_n873), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1104), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1083), .A2(KEYINPUT116), .A3(new_n1086), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1108), .A2(new_n1111), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1100), .A2(new_n1114), .A3(new_n676), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n863), .A2(new_n743), .A3(new_n872), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n366), .B1(new_n763), .B2(new_n239), .C1(new_n244), .C2(new_n760), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1060), .A2(new_n810), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n781), .B2(new_n772), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1117), .B(new_n1119), .C1(G294), .C2(new_n755), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n242), .B2(new_n750), .C1(new_n237), .C2(new_n824), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n770), .A2(new_n370), .B1(new_n752), .B2(new_n204), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n366), .B1(new_n755), .B2(G125), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n814), .B2(new_n760), .ZN(new_n1124));
  XOR2_X1   g0924(.A(KEYINPUT54), .B(G143), .Z(new_n1125));
  AOI211_X1 g0925(.A(new_n1122), .B(new_n1124), .C1(new_n764), .C2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(G128), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n772), .C1(new_n979), .C2(new_n824), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n812), .A2(G150), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT53), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1121), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1131), .A2(new_n746), .B1(new_n284), .B2(new_n827), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1116), .A2(new_n735), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n734), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1068), .B1(new_n1115), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1115), .A2(new_n1068), .A3(new_n1135), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(G378));
  AND3_X1   g0939(.A1(new_n897), .A2(new_n899), .A3(new_n862), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1092), .B1(new_n863), .B2(new_n872), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1140), .A2(new_n1141), .A3(new_n876), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n297), .A2(new_n841), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n444), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n618), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n319), .A2(new_n444), .A3(new_n1143), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT55), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT56), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n618), .A2(new_n1145), .A3(new_n1144), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1143), .B1(new_n319), .B2(new_n444), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT55), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT56), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n918), .B2(G330), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n855), .A2(new_n860), .A3(new_n861), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n912), .B1(new_n1160), .B2(new_n915), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n916), .A2(new_n917), .ZN(new_n1162));
  AND4_X1   g0962(.A1(G330), .A2(new_n1161), .A3(new_n1158), .A4(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1142), .B1(new_n1159), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1161), .A2(new_n1162), .A3(G330), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1158), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n918), .A2(G330), .A3(new_n1158), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1167), .A2(new_n901), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1164), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n734), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n827), .A2(new_n204), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G41), .B(new_n976), .C1(G107), .C2(new_n806), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G97), .A2(new_n767), .B1(new_n1006), .B2(G58), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n600), .A2(new_n764), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n259), .B(new_n1010), .C1(G283), .C2(new_n755), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G116), .B2(new_n773), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT58), .Z(new_n1179));
  OAI21_X1  g0979(.A(new_n204), .B1(new_n320), .B2(G41), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n812), .A2(new_n1125), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT118), .Z(new_n1182));
  NAND2_X1  g0982(.A1(new_n806), .A2(G128), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G150), .A2(new_n818), .B1(new_n773), .B2(G125), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n767), .A2(G132), .B1(new_n764), .B2(G137), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(G33), .B1(new_n755), .B2(G124), .ZN(new_n1189));
  AOI21_X1  g0989(.A(G41), .B1(new_n1006), .B2(new_n756), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1179), .A2(new_n1180), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n801), .B1(new_n1192), .B2(new_n746), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1172), .B(new_n1193), .C1(new_n1166), .C2(new_n744), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT120), .Z(new_n1195));
  NAND2_X1  g0995(.A1(new_n1171), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1100), .A2(new_n1086), .B1(new_n1169), .B2(new_n1164), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n676), .B1(new_n1198), .B2(KEYINPUT57), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1108), .A2(new_n1113), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1200));
  OAI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1200), .B2(new_n1085), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1164), .A2(KEYINPUT121), .A3(new_n1169), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT121), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1167), .A2(new_n901), .A3(new_n1168), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1197), .B1(new_n1199), .B2(new_n1206), .ZN(G375));
  NOR2_X1   g1007(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n1085), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1108), .A2(new_n1209), .A3(new_n1113), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(new_n945), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT122), .Z(new_n1212));
  NAND2_X1  g1012(.A1(new_n973), .A2(new_n1125), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n818), .A2(G50), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n259), .B1(new_n754), .B2(new_n1127), .C1(new_n760), .C2(new_n979), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G150), .B2(new_n764), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n761), .A2(new_n752), .B1(new_n750), .B2(new_n370), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G132), .B2(new_n773), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1213), .A2(new_n1214), .A3(new_n1216), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n973), .A2(G116), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n750), .A2(new_n239), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n975), .B(new_n1221), .C1(G294), .C2(new_n773), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n366), .B1(new_n760), .B2(new_n781), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G107), .B2(new_n764), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1220), .A2(new_n1013), .A3(new_n1222), .A4(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n754), .A2(new_n782), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1219), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1227), .A2(new_n746), .B1(new_n338), .B2(new_n827), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n735), .B(new_n1228), .C1(new_n892), .C2(new_n744), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1208), .B2(new_n733), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1212), .A2(new_n1231), .ZN(G381));
  INV_X1    g1032(.A(new_n1066), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1234), .A2(new_n996), .A3(new_n970), .A4(new_n1043), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1235), .A2(G396), .A3(G393), .ZN(new_n1236));
  INV_X1    g1036(.A(G384), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1236), .A2(new_n1237), .A3(new_n1231), .A4(new_n1212), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(KEYINPUT123), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(KEYINPUT123), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1115), .A2(new_n1135), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(G375), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1239), .A2(new_n1240), .A3(new_n1242), .ZN(G407));
  INV_X1    g1043(.A(G213), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1242), .B2(new_n657), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(G407), .A2(new_n1245), .ZN(G409));
  NAND3_X1  g1046(.A1(new_n1202), .A2(new_n734), .A3(new_n1204), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1100), .A2(new_n1086), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1170), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1195), .B(new_n1247), .C1(new_n1249), .C2(new_n945), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1241), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1115), .A2(new_n1068), .A3(new_n1135), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(new_n1136), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1252), .B1(G375), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT60), .B1(new_n1208), .B2(new_n1085), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n677), .B(new_n1256), .C1(new_n1210), .C2(KEYINPUT60), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1237), .B1(new_n1257), .B2(new_n1230), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1256), .B1(new_n1210), .B2(KEYINPUT60), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n676), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(G384), .A3(new_n1231), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1244), .A2(G343), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1255), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT62), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(G2897), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1258), .A2(new_n1261), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1268), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT57), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n677), .B1(new_n1249), .B2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1248), .A2(KEYINPUT57), .A3(new_n1204), .A4(new_n1202), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1196), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1275), .A2(G378), .B1(new_n1251), .B2(new_n1250), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1271), .B1(new_n1276), .B2(new_n1263), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1255), .A2(new_n1278), .A3(new_n1262), .A4(new_n1264), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1266), .A2(new_n1267), .A3(new_n1277), .A4(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT125), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1255), .A2(new_n1264), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT61), .B1(new_n1283), .B2(new_n1271), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1284), .A2(new_n1266), .A3(KEYINPUT125), .A4(new_n1279), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(G393), .B(G396), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(KEYINPUT124), .B1(G390), .B2(G387), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n1234), .A2(new_n1043), .B1(new_n970), .B2(new_n996), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1287), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT126), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G390), .A2(G387), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1292), .A2(new_n1235), .A3(KEYINPUT124), .A4(new_n1286), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1290), .A2(new_n1291), .A3(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1291), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1282), .A2(new_n1285), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1277), .A2(KEYINPUT63), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1298), .B2(new_n1265), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1255), .A2(KEYINPUT63), .A3(new_n1262), .A4(new_n1264), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1297), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(KEYINPUT127), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT127), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1297), .A2(new_n1302), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(G405));
  NAND2_X1  g1107(.A1(G375), .A2(new_n1251), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1308), .B1(new_n1254), .B2(G375), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1309), .B(new_n1262), .ZN(new_n1310));
  XOR2_X1   g1110(.A(new_n1310), .B(new_n1301), .Z(G402));
endmodule


