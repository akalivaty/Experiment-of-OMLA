//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1284, new_n1285,
    new_n1286, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(G50), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G77), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT64), .ZN(G353));
  NOR2_X1   g0008(.A1(G97), .A2(G107), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G87), .ZN(G355));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT65), .Z(new_n213));
  XOR2_X1   g0013(.A(KEYINPUT67), .B(G244), .Z(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G107), .A2(G264), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n213), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n213), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n204), .A2(KEYINPUT66), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n204), .A2(KEYINPUT66), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n230), .A2(G50), .A3(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n223), .B(new_n226), .C1(new_n229), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n205), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n202), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n246), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G223), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT68), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(KEYINPUT68), .A3(G1698), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n253), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(G1698), .B1(new_n262), .B2(new_n263), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G222), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(new_n215), .B2(new_n264), .ZN(new_n269));
  OR3_X1    g0069(.A1(new_n266), .A2(new_n269), .A3(KEYINPUT69), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT69), .B1(new_n266), .B2(new_n269), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n271), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n276), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n277), .B1(G226), .B2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G179), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n228), .A2(new_n261), .A3(KEYINPUT72), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT72), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(G20), .B2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n206), .A2(G20), .B1(new_n287), .B2(G150), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT71), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT8), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G58), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT70), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(KEYINPUT70), .A3(G58), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n294), .A2(new_n289), .A3(new_n295), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n228), .A2(G33), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n288), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n227), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n275), .A2(G13), .A3(G20), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(new_n227), .A3(new_n302), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT73), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT73), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n306), .A2(new_n309), .B1(new_n275), .B2(G20), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  MUX2_X1   g0111(.A(new_n305), .B(new_n311), .S(G50), .Z(new_n312));
  NAND2_X1  g0112(.A1(new_n304), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n283), .B(new_n313), .C1(G169), .C2(new_n281), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT75), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n304), .A2(new_n315), .A3(new_n312), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n315), .B1(new_n304), .B2(new_n312), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT9), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n318), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT9), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(new_n316), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT10), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(new_n273), .B2(new_n280), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n326), .B1(G190), .B2(new_n281), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n323), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n324), .B1(new_n323), .B2(new_n327), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n314), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT13), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n267), .A2(G226), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G97), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n264), .A2(G232), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n333), .B(new_n334), .C1(new_n258), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n271), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n277), .B1(G238), .B2(new_n279), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n332), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(new_n332), .A3(new_n338), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G200), .ZN(new_n343));
  AOI211_X1 g0143(.A(new_n202), .B(new_n306), .C1(new_n275), .C2(G20), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT76), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n284), .A2(new_n286), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(new_n205), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n300), .A2(new_n215), .B1(new_n228), .B2(G68), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n303), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT11), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n305), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n202), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT12), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n349), .A2(new_n350), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n345), .A2(new_n351), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n340), .A2(G190), .A3(new_n341), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n343), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n341), .ZN(new_n360));
  OAI21_X1  g0160(.A(G169), .B1(new_n360), .B2(new_n339), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT14), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT14), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n342), .A2(new_n363), .A3(G169), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n340), .A2(G179), .A3(new_n341), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n359), .B1(new_n366), .B2(new_n356), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G33), .A2(G41), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(G1), .A3(G13), .ZN(new_n369));
  OAI211_X1 g0169(.A(G226), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT78), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n264), .A2(KEYINPUT78), .A3(G226), .A4(G1698), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(G223), .B(new_n258), .C1(new_n255), .C2(new_n256), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G87), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n376), .A2(KEYINPUT79), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(KEYINPUT79), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n369), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n277), .ZN(new_n381));
  INV_X1    g0181(.A(new_n279), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n381), .B1(new_n382), .B2(new_n236), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n325), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G190), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n277), .B1(G232), .B2(new_n279), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n372), .B2(new_n373), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n385), .B(new_n386), .C1(new_n388), .C2(new_n369), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n257), .B2(new_n228), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n262), .A2(KEYINPUT7), .A3(new_n228), .A4(new_n263), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G58), .A2(G68), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n203), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G20), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT77), .ZN(new_n398));
  INV_X1    g0198(.A(G159), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n397), .B(new_n398), .C1(new_n346), .C2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n284), .B2(new_n286), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n228), .B1(new_n203), .B2(new_n395), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT77), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n394), .A2(new_n400), .A3(KEYINPUT16), .A4(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n262), .A2(new_n228), .A3(new_n263), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n202), .B1(new_n408), .B2(new_n392), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n397), .B1(new_n346), .B2(new_n399), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n405), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n404), .A2(new_n303), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n297), .A2(new_n308), .A3(new_n310), .A4(new_n298), .ZN(new_n413));
  INV_X1    g0213(.A(new_n298), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n352), .B1(new_n414), .B2(new_n296), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n390), .A2(KEYINPUT80), .A3(new_n412), .A4(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n412), .A2(new_n416), .ZN(new_n420));
  OAI21_X1  g0220(.A(G169), .B1(new_n380), .B2(new_n383), .ZN(new_n421));
  OAI211_X1 g0221(.A(G179), .B(new_n386), .C1(new_n388), .C2(new_n369), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT18), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n412), .A2(new_n416), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n426), .A2(KEYINPUT80), .A3(KEYINPUT17), .A4(new_n390), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n420), .A2(new_n423), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n419), .A2(new_n425), .A3(new_n427), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n259), .A2(new_n265), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n432), .A2(G238), .ZN(new_n433));
  INV_X1    g0233(.A(G107), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n335), .A2(G1698), .B1(new_n434), .B2(new_n264), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n271), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n214), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n277), .B1(new_n437), .B2(new_n279), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G169), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n436), .A2(new_n282), .A3(new_n438), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n290), .A2(new_n292), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n346), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT15), .B(G87), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n446), .A2(new_n300), .B1(new_n228), .B2(new_n215), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n303), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n215), .B1(new_n275), .B2(G20), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n307), .A2(new_n449), .B1(new_n215), .B2(new_n352), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n441), .A2(new_n442), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n325), .B1(new_n436), .B2(new_n438), .ZN(new_n453));
  OR3_X1    g0253(.A1(new_n453), .A2(KEYINPUT74), .A3(new_n451), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT74), .B1(new_n453), .B2(new_n451), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n436), .A2(G190), .A3(new_n438), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n367), .A2(new_n431), .A3(new_n452), .A4(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT81), .B1(new_n331), .B2(new_n458), .ZN(new_n459));
  AND4_X1   g0259(.A1(new_n431), .A2(new_n367), .A3(new_n452), .A4(new_n457), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n323), .A2(new_n327), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT10), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n328), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT81), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n460), .A2(new_n463), .A3(new_n464), .A4(new_n314), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n459), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n264), .A2(G264), .A3(G1698), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n264), .A2(G257), .A3(new_n258), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n257), .A2(G303), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n271), .ZN(new_n471));
  INV_X1    g0271(.A(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G1), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT5), .B(G41), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n271), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n271), .A2(new_n274), .ZN(new_n476));
  AND2_X1   g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n475), .A2(G270), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n440), .B1(new_n471), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT21), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n302), .A2(new_n227), .B1(G20), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  INV_X1    g0286(.A(G97), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n486), .B(new_n228), .C1(G33), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT20), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n485), .A2(KEYINPUT20), .A3(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n305), .A2(new_n484), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n261), .A2(G1), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n306), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n496), .B2(new_n484), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n483), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n482), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT85), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT86), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n471), .A2(new_n481), .A3(G179), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n493), .A2(new_n497), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n482), .A2(KEYINPUT85), .A3(new_n498), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n501), .A2(new_n502), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT85), .B1(new_n482), .B2(new_n498), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT86), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT21), .B1(new_n482), .B2(new_n504), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n474), .A2(G274), .A3(new_n369), .A4(new_n473), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n479), .A2(new_n369), .ZN(new_n514));
  INV_X1    g0314(.A(G270), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n271), .B2(new_n470), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G190), .ZN(new_n518));
  INV_X1    g0318(.A(new_n504), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n518), .B(new_n519), .C1(new_n325), .C2(new_n517), .ZN(new_n520));
  AND4_X1   g0320(.A1(new_n507), .A2(new_n510), .A3(new_n512), .A4(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT25), .B1(new_n352), .B2(new_n434), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n352), .A2(KEYINPUT25), .A3(new_n434), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n523), .A2(new_n524), .B1(new_n496), .B2(G107), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n479), .A2(G264), .A3(new_n369), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT90), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT90), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n479), .A2(new_n528), .A3(G264), .A4(new_n369), .ZN(new_n529));
  OAI211_X1 g0329(.A(G257), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n530));
  OAI211_X1 g0330(.A(G250), .B(new_n258), .C1(new_n255), .C2(new_n256), .ZN(new_n531));
  INV_X1    g0331(.A(G294), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n530), .B(new_n531), .C1(new_n261), .C2(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n527), .A2(new_n529), .B1(new_n533), .B2(new_n271), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n513), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n325), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n526), .A2(new_n513), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n271), .B2(new_n533), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n385), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT89), .ZN(new_n541));
  OAI21_X1  g0341(.A(KEYINPUT23), .B1(new_n228), .B2(G107), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT23), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n434), .A3(G20), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n228), .A2(G33), .A3(G116), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT88), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT88), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n542), .A2(new_n544), .A3(new_n545), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n228), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT22), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT22), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n264), .A2(new_n553), .A3(new_n228), .A4(G87), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g0356(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n550), .A2(new_n555), .A3(new_n557), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n541), .B1(new_n561), .B2(new_n303), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n550), .A2(new_n555), .A3(new_n557), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n557), .B1(new_n550), .B2(new_n555), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n541), .B(new_n303), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n525), .B(new_n540), .C1(new_n562), .C2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n535), .A2(new_n282), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n538), .A2(new_n440), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n525), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n303), .B1(new_n563), .B2(new_n564), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT89), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n571), .B1(new_n573), .B2(new_n565), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n567), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n305), .A2(G97), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n496), .B2(G97), .ZN(new_n577));
  OAI21_X1  g0377(.A(G107), .B1(new_n391), .B2(new_n393), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n215), .B1(new_n284), .B2(new_n286), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT6), .ZN(new_n580));
  AND2_X1   g0380(.A1(G97), .A2(G107), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(new_n209), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n434), .A2(KEYINPUT6), .A3(G97), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n579), .B1(new_n584), .B2(G20), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT82), .B1(new_n586), .B2(new_n303), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT82), .ZN(new_n588));
  INV_X1    g0388(.A(new_n303), .ZN(new_n589));
  AOI211_X1 g0389(.A(new_n588), .B(new_n589), .C1(new_n578), .C2(new_n585), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n577), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(G257), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n513), .B1(new_n514), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(G244), .B(new_n258), .C1(new_n255), .C2(new_n256), .ZN(new_n595));
  XOR2_X1   g0395(.A(KEYINPUT83), .B(KEYINPUT4), .Z(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT84), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(G250), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT4), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n486), .B(new_n599), .C1(new_n595), .C2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT84), .B1(new_n595), .B2(new_n596), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n594), .B1(new_n603), .B2(new_n369), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n440), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n595), .A2(new_n596), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT84), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n267), .A2(KEYINPUT4), .A3(G244), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n599), .A2(new_n486), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n608), .A2(new_n597), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n593), .B1(new_n611), .B2(new_n271), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n282), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n591), .A2(new_n605), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n577), .ZN(new_n615));
  INV_X1    g0415(.A(new_n579), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n434), .A2(KEYINPUT6), .A3(G97), .ZN(new_n617));
  XNOR2_X1  g0417(.A(G97), .B(G107), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n580), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n616), .B1(new_n619), .B2(new_n228), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n434), .B1(new_n408), .B2(new_n392), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n303), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n588), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n586), .A2(KEYINPUT82), .A3(new_n303), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n615), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AOI211_X1 g0425(.A(G190), .B(new_n593), .C1(new_n611), .C2(new_n271), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n611), .A2(new_n271), .ZN(new_n627));
  AOI21_X1  g0427(.A(G200), .B1(new_n627), .B2(new_n594), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n625), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(G238), .B(new_n258), .C1(new_n255), .C2(new_n256), .ZN(new_n630));
  OAI211_X1 g0430(.A(G244), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n631));
  NAND2_X1  g0431(.A1(G33), .A2(G116), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n271), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n369), .A2(G274), .A3(new_n473), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n275), .A2(G45), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n369), .A2(G250), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G200), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n264), .A2(new_n228), .A3(G68), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT19), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n228), .B1(new_n334), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(G87), .B2(new_n210), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n643), .B1(new_n300), .B2(new_n487), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n642), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n647), .A2(new_n303), .B1(new_n352), .B2(new_n446), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n638), .B1(new_n271), .B2(new_n633), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G190), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n496), .A2(G87), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n641), .A2(new_n648), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(new_n303), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n446), .A2(new_n352), .ZN(new_n654));
  INV_X1    g0454(.A(new_n446), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n496), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n649), .A2(new_n282), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n657), .B(new_n658), .C1(G169), .C2(new_n649), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n652), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n614), .A2(new_n629), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n575), .A2(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n466), .A2(new_n521), .A3(new_n662), .ZN(G372));
  INV_X1    g0463(.A(new_n659), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n652), .A2(new_n659), .ZN(new_n666));
  OR3_X1    g0466(.A1(new_n614), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n665), .B1(new_n614), .B2(new_n666), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n614), .A2(new_n629), .A3(new_n660), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n567), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n501), .A2(new_n505), .A3(new_n506), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(new_n511), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n574), .A2(new_n570), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n669), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n466), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n329), .A2(new_n330), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n425), .A2(new_n429), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n366), .A2(new_n356), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n359), .B2(new_n452), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n419), .A2(new_n427), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n314), .B1(new_n678), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT91), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI211_X1 g0486(.A(KEYINPUT91), .B(new_n314), .C1(new_n678), .C2(new_n683), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n677), .A2(new_n688), .ZN(G369));
  NAND3_X1  g0489(.A1(new_n275), .A2(new_n228), .A3(G13), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n519), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n673), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n511), .B1(new_n672), .B2(KEYINPUT86), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n507), .A3(new_n520), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n698), .B1(new_n700), .B2(new_n697), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G330), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n574), .A2(new_n696), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n525), .B1(new_n562), .B2(new_n566), .ZN(new_n705));
  INV_X1    g0505(.A(new_n570), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n575), .A2(new_n704), .B1(new_n707), .B2(new_n696), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n695), .B1(new_n699), .B2(new_n507), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(new_n707), .A3(new_n567), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n674), .A2(new_n696), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n709), .A2(new_n713), .ZN(G399));
  INV_X1    g0514(.A(new_n224), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G87), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n209), .A2(new_n718), .A3(new_n484), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT92), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(G1), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n232), .B2(new_n717), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n661), .B1(new_n574), .B2(new_n540), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(new_n674), .B2(new_n673), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n695), .B1(new_n725), .B2(new_n669), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n699), .A2(new_n707), .A3(new_n507), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT95), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT95), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n699), .A2(new_n707), .A3(new_n731), .A4(new_n507), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(new_n724), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n695), .B1(new_n733), .B2(new_n669), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n728), .B1(new_n734), .B2(new_n727), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT30), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n517), .A2(G179), .A3(new_n534), .A4(new_n649), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n736), .B1(new_n737), .B2(new_n604), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n634), .A2(new_n639), .A3(KEYINPUT93), .ZN(new_n739));
  AOI21_X1  g0539(.A(KEYINPUT93), .B1(new_n634), .B2(new_n639), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(G179), .B1(new_n471), .B2(new_n481), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n741), .A2(new_n604), .A3(new_n535), .A4(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n534), .A2(new_n649), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(KEYINPUT30), .A3(new_n503), .A4(new_n612), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n738), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT31), .B1(new_n746), .B2(new_n695), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT94), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n670), .A2(new_n707), .A3(new_n567), .A4(new_n696), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n751), .B1(new_n752), .B2(new_n700), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n662), .A2(KEYINPUT94), .A3(new_n521), .A4(new_n696), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G330), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n735), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n723), .B1(new_n758), .B2(G1), .ZN(G364));
  AND2_X1   g0559(.A1(new_n228), .A2(G13), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n275), .B1(new_n760), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n716), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n703), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(G330), .B2(new_n701), .ZN(new_n765));
  INV_X1    g0565(.A(new_n763), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n227), .B1(G20), .B2(new_n440), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G190), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n487), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n325), .A2(G179), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(G20), .A3(G190), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n769), .A2(G20), .A3(new_n385), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G159), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n264), .B1(new_n775), .B2(new_n718), .C1(new_n778), .C2(KEYINPUT32), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n773), .B(new_n779), .C1(KEYINPUT32), .C2(new_n778), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n228), .A2(new_n282), .A3(KEYINPUT97), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT97), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(G20), .B2(G179), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n784), .A2(new_n385), .A3(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G58), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n774), .A2(G20), .A3(new_n385), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT99), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(KEYINPUT99), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n434), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n784), .A2(G190), .A3(G200), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n791), .B1(G77), .B2(new_n792), .ZN(new_n793));
  AND3_X1   g0593(.A1(new_n780), .A2(new_n786), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(G200), .B1(new_n781), .B2(new_n783), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT98), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n385), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n796), .A2(G190), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n794), .B1(new_n205), .B2(new_n798), .C1(new_n202), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n785), .ZN(new_n802));
  INV_X1    g0602(.A(G322), .ZN(new_n803));
  INV_X1    g0603(.A(G283), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n802), .A2(new_n803), .B1(new_n790), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G311), .B2(new_n792), .ZN(new_n806));
  XNOR2_X1  g0606(.A(KEYINPUT33), .B(G317), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n799), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n797), .A2(G326), .ZN(new_n809));
  INV_X1    g0609(.A(G329), .ZN(new_n810));
  INV_X1    g0610(.A(G303), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n257), .B1(new_n776), .B2(new_n810), .C1(new_n775), .C2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G294), .B2(new_n771), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n806), .A2(new_n808), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n768), .B1(new_n801), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(G13), .A2(G33), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G20), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n767), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n224), .A2(G355), .A3(new_n264), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n715), .A2(new_n264), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n472), .B2(new_n233), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n824), .A2(KEYINPUT96), .B1(new_n472), .B2(new_n251), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n824), .A2(KEYINPUT96), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n820), .B1(G116), .B2(new_n224), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n766), .B(new_n815), .C1(new_n819), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n818), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n701), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n765), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G396));
  INV_X1    g0632(.A(new_n792), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n484), .A2(new_n833), .B1(new_n802), .B2(new_n532), .ZN(new_n834));
  INV_X1    g0634(.A(G311), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n257), .B1(new_n776), .B2(new_n835), .C1(new_n775), .C2(new_n434), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n790), .A2(new_n718), .ZN(new_n837));
  NOR4_X1   g0637(.A1(new_n834), .A2(new_n773), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n838), .B1(new_n798), .B2(new_n811), .C1(new_n804), .C2(new_n800), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G143), .A2(new_n785), .B1(new_n792), .B2(G159), .ZN(new_n840));
  INV_X1    g0640(.A(G137), .ZN(new_n841));
  INV_X1    g0641(.A(G150), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n840), .B1(new_n798), .B2(new_n841), .C1(new_n842), .C2(new_n800), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT34), .Z(new_n844));
  INV_X1    g0644(.A(new_n790), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(G68), .ZN(new_n846));
  INV_X1    g0646(.A(G132), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n264), .B1(new_n776), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n775), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(G50), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n846), .B(new_n850), .C1(new_n201), .C2(new_n772), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n839), .B1(new_n844), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n767), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n767), .A2(new_n816), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n766), .B1(new_n215), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n452), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n451), .A2(new_n695), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n457), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n452), .A2(new_n695), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n853), .B(new_n855), .C1(new_n817), .C2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n860), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n726), .B(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n757), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n763), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n864), .A2(new_n865), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n861), .B1(new_n867), .B2(new_n868), .ZN(G384));
  INV_X1    g0669(.A(new_n693), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n420), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n430), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n390), .A2(new_n412), .A3(new_n416), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(new_n424), .A3(new_n871), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT37), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n874), .A2(new_n424), .A3(new_n871), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT39), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n413), .A2(new_n415), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n404), .A2(new_n303), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n394), .A2(new_n403), .A3(new_n400), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n405), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n884), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n423), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n874), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n888), .A2(new_n693), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n878), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n430), .A2(new_n891), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT38), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n882), .A2(new_n883), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT100), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n893), .A2(new_n894), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n881), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT100), .A4(KEYINPUT38), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n897), .B1(KEYINPUT39), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n366), .A2(new_n356), .A3(new_n696), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n359), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n356), .A2(new_n695), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n680), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n356), .B(new_n695), .C1(new_n359), .C2(new_n366), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n676), .A2(new_n860), .A3(new_n696), .ZN(new_n913));
  INV_X1    g0713(.A(new_n859), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n903), .ZN(new_n916));
  INV_X1    g0716(.A(new_n679), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n916), .B1(new_n917), .B2(new_n870), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n906), .A2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n466), .A2(new_n735), .B1(new_n686), .B2(new_n687), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n919), .B(new_n920), .Z(new_n921));
  INV_X1    g0721(.A(KEYINPUT102), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n749), .B1(new_n747), .B2(new_n922), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n746), .A2(KEYINPUT102), .A3(KEYINPUT31), .A4(new_n695), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n575), .A2(new_n661), .A3(new_n695), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT94), .B1(new_n927), .B2(new_n521), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n752), .A2(new_n751), .A3(new_n700), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n911), .A2(new_n860), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT103), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n925), .B1(new_n753), .B2(new_n754), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n911), .A2(new_n860), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT103), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n882), .B2(new_n895), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n933), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n903), .A2(new_n930), .A3(new_n931), .ZN(new_n940));
  XOR2_X1   g0740(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n466), .A2(new_n930), .ZN(new_n944));
  OAI21_X1  g0744(.A(G330), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n921), .A2(new_n946), .B1(new_n275), .B2(new_n760), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n921), .B2(new_n946), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n584), .A2(KEYINPUT35), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n584), .A2(KEYINPUT35), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n949), .A2(new_n950), .A3(G116), .A4(new_n229), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT36), .Z(new_n952));
  NAND3_X1  g0752(.A1(new_n233), .A2(G77), .A3(new_n395), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n275), .B(G13), .C1(new_n953), .C2(new_n247), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n948), .A2(new_n952), .A3(new_n954), .ZN(G367));
  OR2_X1    g0755(.A1(new_n614), .A2(new_n696), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n614), .B(new_n629), .C1(new_n625), .C2(new_n696), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n711), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT42), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n614), .B1(new_n957), .B2(new_n707), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n961), .A2(KEYINPUT42), .B1(new_n696), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n648), .A2(new_n651), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n695), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n660), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n659), .A2(new_n966), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n962), .A2(new_n964), .B1(KEYINPUT43), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n970), .B(new_n971), .Z(new_n972));
  NOR2_X1   g0772(.A1(new_n709), .A2(new_n959), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT104), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n713), .A2(new_n958), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT44), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n978), .B2(new_n977), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n977), .A2(new_n976), .A3(new_n978), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n713), .A2(new_n958), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT45), .Z(new_n983));
  NAND3_X1  g0783(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT105), .ZN(new_n985));
  INV_X1    g0785(.A(new_n709), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n711), .B1(new_n708), .B2(new_n710), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n703), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n758), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n709), .A2(KEYINPUT105), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n980), .A2(new_n709), .A3(new_n981), .A4(new_n983), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n987), .A2(new_n991), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n758), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n716), .B(KEYINPUT41), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n762), .B1(new_n998), .B2(KEYINPUT106), .ZN(new_n999));
  AOI211_X1 g0799(.A(KEYINPUT106), .B(new_n996), .C1(new_n994), .C2(new_n758), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n975), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G283), .A2(new_n792), .B1(new_n785), .B2(G303), .ZN(new_n1003));
  XOR2_X1   g0803(.A(KEYINPUT107), .B(G317), .Z(new_n1004));
  OAI21_X1  g0804(.A(new_n257), .B1(new_n1004), .B2(new_n776), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n775), .A2(new_n484), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n1006), .A2(KEYINPUT46), .B1(new_n772), .B2(new_n434), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1005), .B(new_n1007), .C1(KEYINPUT46), .C2(new_n1006), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n790), .A2(new_n487), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n1003), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n798), .B2(new_n835), .C1(new_n532), .C2(new_n800), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n799), .A2(G159), .B1(G50), .B2(new_n792), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n1014), .A2(KEYINPUT108), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n257), .B1(new_n849), .B2(G58), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n771), .A2(G68), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n841), .C2(new_n776), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n802), .A2(new_n842), .B1(new_n790), .B2(new_n215), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(new_n797), .C2(G143), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n1014), .B2(KEYINPUT108), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1012), .B1(new_n1015), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT47), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n768), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n1023), .B2(new_n1022), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n967), .A2(new_n818), .A3(new_n968), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n821), .A2(new_n242), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n818), .B(new_n767), .C1(new_n715), .C2(new_n655), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n766), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AND3_X1   g0829(.A1(new_n1025), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1002), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(G387));
  NAND2_X1  g0832(.A1(new_n989), .A2(new_n762), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT109), .Z(new_n1034));
  OR2_X1    g0834(.A1(new_n708), .A2(new_n829), .ZN(new_n1035));
  OR3_X1    g0835(.A1(new_n239), .A2(new_n472), .A3(new_n264), .ZN(new_n1036));
  OAI21_X1  g0836(.A(KEYINPUT50), .B1(new_n444), .B2(G50), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1037), .B(new_n472), .C1(new_n202), .C2(new_n215), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n444), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n257), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n720), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n715), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n819), .B1(new_n224), .B2(new_n434), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n763), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n257), .B1(new_n849), .B2(G77), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n842), .B2(new_n776), .C1(new_n446), .C2(new_n772), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1010), .B1(new_n205), .B2(new_n802), .C1(new_n202), .C2(new_n833), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n299), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1046), .B(new_n1047), .C1(new_n799), .C2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n399), .B2(new_n798), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n772), .A2(new_n804), .B1(new_n775), .B2(new_n532), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1004), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G303), .A2(new_n792), .B1(new_n785), .B2(new_n1052), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n798), .B2(new_n803), .C1(new_n835), .C2(new_n800), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1055), .B2(new_n1054), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT49), .Z(new_n1058));
  AOI21_X1  g0858(.A(new_n264), .B1(new_n777), .B2(G326), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n790), .B2(new_n484), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1050), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1044), .B1(new_n1061), .B2(new_n767), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1034), .B1(new_n1035), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(KEYINPUT110), .B1(new_n990), .B2(new_n716), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n990), .A2(KEYINPUT110), .A3(new_n716), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n758), .B2(new_n989), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1063), .B1(new_n1064), .B2(new_n1066), .ZN(G393));
  NOR2_X1   g0867(.A1(new_n822), .A2(new_n246), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n819), .B1(new_n224), .B2(new_n487), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n763), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n791), .B1(G294), .B2(new_n792), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n257), .B1(new_n775), .B2(new_n804), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G322), .B2(new_n777), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(new_n484), .C2(new_n772), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n799), .B2(G303), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n797), .A2(G317), .B1(G311), .B2(new_n785), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT52), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1075), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1080), .A2(KEYINPUT112), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n797), .A2(G150), .B1(G159), .B2(new_n785), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT51), .Z(new_n1083));
  AOI22_X1  g0883(.A1(new_n799), .A2(G50), .B1(new_n443), .B2(new_n792), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1084), .A2(KEYINPUT111), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(KEYINPUT111), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n257), .B1(new_n777), .B2(G143), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n771), .A2(G77), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(new_n202), .C2(new_n775), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n837), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .A4(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1080), .A2(KEYINPUT112), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1081), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1070), .B1(new_n1093), .B2(new_n767), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n829), .B2(new_n958), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n984), .A2(new_n986), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n993), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1095), .B1(new_n1097), .B2(new_n761), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT113), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n990), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1100), .A2(new_n716), .A3(new_n994), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1099), .A2(new_n1101), .ZN(G390));
  INV_X1    g0902(.A(new_n905), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n882), .B2(new_n895), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n858), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n859), .B1(new_n734), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1104), .B1(new_n1106), .B2(new_n912), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n903), .A2(KEYINPUT39), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1108), .B(new_n896), .C1(new_n915), .C2(new_n1103), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n755), .A2(new_n756), .A3(new_n862), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n911), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1107), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n753), .A2(new_n754), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n756), .B1(new_n1113), .B2(new_n926), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n931), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n762), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n854), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n763), .B1(new_n1048), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n846), .B1(new_n532), .B2(new_n776), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1121), .A2(KEYINPUT117), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(KEYINPUT117), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n264), .B1(new_n849), .B2(G87), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1088), .B(new_n1124), .C1(new_n802), .C2(new_n484), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G97), .B2(new_n792), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1122), .A2(new_n1123), .A3(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n434), .A2(new_n800), .B1(new_n798), .B2(new_n804), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n264), .B1(new_n790), .B2(new_n205), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT116), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1132));
  INV_X1    g0932(.A(G125), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n772), .A2(new_n399), .B1(new_n1133), .B2(new_n776), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT53), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n775), .B2(new_n842), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n849), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G132), .A2(new_n785), .B1(new_n792), .B2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1131), .A2(new_n1132), .A3(new_n1138), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(G128), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1143), .A2(new_n798), .B1(new_n800), .B2(new_n841), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n1127), .A2(new_n1128), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1120), .B1(new_n1145), .B2(new_n767), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n904), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n817), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1118), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1114), .A2(new_n860), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n912), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1151), .A2(new_n1111), .A3(new_n1106), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n750), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1113), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(G330), .A3(new_n860), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1155), .A2(new_n912), .B1(new_n931), .B2(new_n1114), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT114), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n859), .B1(new_n726), .B2(new_n860), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1115), .B1(new_n1110), .B2(new_n911), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n913), .A2(new_n914), .ZN(new_n1161));
  AOI21_X1  g0961(.A(KEYINPUT114), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1152), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n466), .A2(new_n1114), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n920), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1163), .A2(new_n1117), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT115), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1157), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1160), .A2(KEYINPUT114), .A3(new_n1161), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1165), .B1(new_n1171), .B2(new_n1152), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT115), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n1173), .A3(new_n1117), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1168), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1172), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1107), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n905), .B1(new_n1158), .B2(new_n912), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n695), .B(new_n858), .C1(new_n733), .C2(new_n669), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n911), .B1(new_n1179), .B2(new_n859), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n904), .A2(new_n1178), .B1(new_n1180), .B2(new_n1104), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1177), .B1(new_n1181), .B2(new_n1115), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n717), .B1(new_n1176), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1149), .B1(new_n1175), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(G378));
  AOI21_X1  g0985(.A(new_n693), .B1(new_n320), .B2(new_n316), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n331), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1186), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n463), .A2(new_n314), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1187), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n816), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n763), .B1(G50), .B2(new_n1119), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1017), .B1(new_n802), .B2(new_n434), .C1(new_n446), .C2(new_n833), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n264), .A2(G41), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n215), .B2(new_n775), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n790), .A2(new_n201), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(G283), .C2(new_n777), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT118), .Z(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n484), .B2(new_n798), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1198), .B(new_n1204), .C1(G97), .C2(new_n799), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1205), .A2(KEYINPUT58), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n772), .A2(new_n842), .B1(new_n1139), .B2(new_n775), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n802), .A2(new_n1143), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(G137), .C2(new_n792), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n798), .B2(new_n1133), .C1(new_n847), .C2(new_n800), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n845), .A2(G159), .ZN(new_n1213));
  AOI211_X1 g1013(.A(G33), .B(G41), .C1(new_n777), .C2(G124), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1205), .A2(KEYINPUT58), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1199), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n205), .C1(G33), .C2(G41), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1206), .A2(new_n1215), .A3(new_n1216), .A4(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1197), .B1(new_n1219), .B2(new_n767), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1196), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT119), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n939), .A2(new_n942), .A3(G330), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1195), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1226), .A2(new_n939), .A3(new_n942), .A4(G330), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n919), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1223), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1225), .A2(new_n919), .A3(new_n1227), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT120), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT120), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1225), .A2(new_n919), .A3(new_n1233), .A4(new_n1227), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1230), .A2(new_n1232), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1232), .A2(new_n1234), .B1(new_n1236), .B2(KEYINPUT119), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1222), .B1(new_n1238), .B2(new_n762), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1173), .B1(new_n1172), .B2(new_n1117), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1111), .A2(new_n1106), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1169), .A2(new_n1170), .B1(new_n1151), .B2(new_n1241), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(new_n1242), .A2(new_n1182), .A3(new_n1165), .A4(KEYINPUT115), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1166), .B1(new_n1240), .B2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT57), .B1(new_n1238), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1165), .B1(new_n1168), .B2(new_n1174), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT121), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1231), .A2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1225), .A2(new_n919), .A3(KEYINPUT121), .A4(new_n1227), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n1236), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT57), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n716), .B1(new_n1246), .B2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1239), .B1(new_n1245), .B2(new_n1252), .ZN(G375));
  AOI21_X1  g1053(.A(new_n766), .B1(new_n202), .B2(new_n854), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n797), .A2(G294), .B1(G107), .B2(new_n792), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n484), .B2(new_n800), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT122), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n785), .A2(G283), .B1(new_n655), .B2(new_n771), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT123), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n257), .B1(new_n776), .B2(new_n811), .C1(new_n775), .C2(new_n487), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n845), .B2(G77), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1257), .A2(new_n1259), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT124), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n264), .B1(new_n776), .B2(new_n1143), .C1(new_n775), .C2(new_n399), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1201), .B1(G137), .B2(new_n785), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n842), .B2(new_n833), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n1265), .B(new_n1267), .C1(G50), .C2(new_n771), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1268), .B1(new_n847), .B2(new_n798), .C1(new_n800), .C2(new_n1139), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1264), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1254), .B1(new_n817), .B2(new_n911), .C1(new_n1271), .C2(new_n768), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1242), .B2(new_n761), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1172), .A2(new_n996), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1242), .A2(new_n1165), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(G381));
  INV_X1    g1077(.A(G390), .ZN(new_n1278));
  INV_X1    g1078(.A(G384), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NOR4_X1   g1080(.A1(new_n1280), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1281));
  INV_X1    g1081(.A(G375), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1031), .A3(new_n1184), .A4(new_n1282), .ZN(G407));
  NAND2_X1  g1083(.A1(new_n694), .A2(G213), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1282), .A2(new_n1184), .A3(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(G407), .A2(G213), .A3(new_n1286), .ZN(G409));
  INV_X1    g1087(.A(KEYINPUT61), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G378), .B(new_n1239), .C1(new_n1245), .C2(new_n1252), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1230), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1230), .A2(new_n1232), .A3(new_n1234), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1294), .A2(new_n1246), .A3(new_n996), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1250), .A2(new_n762), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1221), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1184), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1285), .B1(new_n1289), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1285), .A2(G2897), .ZN(new_n1300));
  XOR2_X1   g1100(.A(new_n1300), .B(KEYINPUT126), .Z(new_n1301));
  NOR2_X1   g1101(.A1(new_n1172), .A2(new_n717), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT60), .B1(new_n1275), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT60), .ZN(new_n1305));
  AOI211_X1 g1105(.A(KEYINPUT125), .B(new_n1305), .C1(new_n1242), .C2(new_n1165), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1302), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1273), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(G384), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G384), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1301), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1311), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1301), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1313), .A2(new_n1309), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1312), .A2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1288), .B1(new_n1299), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1299), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n996), .B1(new_n994), .B2(new_n758), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT106), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n761), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n974), .B1(new_n1325), .B2(new_n1000), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1030), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1326), .A2(G390), .A3(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(G390), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1330));
  XNOR2_X1  g1130(.A(G393), .B(new_n831), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  NOR3_X1   g1132(.A1(new_n1329), .A2(new_n1330), .A3(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1278), .B1(new_n1002), .B2(new_n1030), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1331), .B1(new_n1334), .B2(new_n1328), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1299), .A2(KEYINPUT63), .A3(new_n1319), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1318), .A2(new_n1322), .A3(new_n1336), .A4(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT62), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1299), .A2(new_n1339), .A3(new_n1319), .ZN(new_n1340));
  XOR2_X1   g1140(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1341));
  AOI21_X1  g1141(.A(new_n1341), .B1(new_n1299), .B2(new_n1319), .ZN(new_n1342));
  NOR3_X1   g1142(.A1(new_n1340), .A2(new_n1317), .A3(new_n1342), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1338), .B1(new_n1343), .B2(new_n1336), .ZN(G405));
  NAND2_X1  g1144(.A1(G375), .A2(new_n1184), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n1289), .ZN(new_n1346));
  OR2_X1    g1146(.A1(new_n1346), .A2(new_n1319), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1319), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1336), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1347), .A2(new_n1336), .A3(new_n1348), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1351), .A2(new_n1352), .ZN(G402));
endmodule


