//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n556, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n576, new_n577, new_n578, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n640, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n461), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n465), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n471), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n461), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n471), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n471), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n472), .B(KEYINPUT69), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  AOI21_X1  g064(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(new_n491), .A3(G138), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n491), .B1(new_n490), .B2(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n471), .A2(G126), .A3(G2105), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n495), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(G50), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT72), .A2(G651), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(KEYINPUT71), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n518), .B1(KEYINPUT72), .B2(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT6), .B1(new_n507), .B2(KEYINPUT71), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n508), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n521), .A2(KEYINPUT73), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n526), .B(new_n517), .C1(new_n519), .C2(new_n520), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n525), .A2(G543), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n515), .A2(KEYINPUT71), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n534), .B(KEYINPUT6), .C1(KEYINPUT71), .C2(new_n507), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n512), .B1(new_n535), .B2(new_n517), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n533), .B1(G89), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n529), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(G168));
  NAND2_X1  g114(.A1(new_n528), .A2(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n512), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n536), .A2(G90), .B1(G651), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n540), .A2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  NAND2_X1  g121(.A1(new_n528), .A2(G43), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n512), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n536), .A2(G81), .B1(G651), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT74), .Z(G188));
  AND2_X1   g134(.A1(G53), .A2(G543), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n525), .A2(new_n527), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(KEYINPUT75), .B(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n525), .A2(new_n527), .A3(new_n560), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n567), .B1(new_n510), .B2(new_n511), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n503), .A2(KEYINPUT76), .A3(new_n504), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G65), .ZN(new_n571));
  INV_X1    g146(.A(G78), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(new_n502), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(G91), .B2(new_n536), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n566), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n529), .A2(new_n576), .A3(new_n537), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n576), .B1(new_n529), .B2(new_n537), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(G286));
  OAI21_X1  g154(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT78), .Z(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(G87), .B2(new_n536), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n528), .A2(G49), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G288));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OR3_X1    g160(.A1(new_n512), .A2(KEYINPUT79), .A3(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT79), .B1(new_n512), .B2(new_n585), .ZN(new_n588));
  INV_X1    g163(.A(G73), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(new_n502), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n592), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n521), .A2(G48), .A3(G543), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n536), .A2(G86), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n594), .A2(new_n595), .A3(new_n598), .A4(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(G72), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G60), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n512), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n536), .A2(G85), .B1(G651), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n525), .A2(G543), .A3(new_n527), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(G290));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NOR2_X1   g185(.A1(G301), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n606), .A2(KEYINPUT83), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT83), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n525), .A2(new_n613), .A3(G543), .A4(new_n527), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n612), .A2(G54), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n536), .A2(KEYINPUT10), .A3(G92), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n521), .A2(new_n505), .ZN(new_n618));
  INV_X1    g193(.A(G92), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n570), .A2(G66), .ZN(new_n621));
  NAND2_X1  g196(.A1(G79), .A2(G543), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n616), .A2(new_n620), .B1(new_n623), .B2(G651), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n615), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n625), .A2(KEYINPUT84), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n625), .A2(KEYINPUT84), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n611), .B1(new_n629), .B2(new_n610), .ZN(G284));
  AOI21_X1  g205(.A(new_n611), .B1(new_n629), .B2(new_n610), .ZN(G321));
  NOR2_X1   g206(.A1(G286), .A2(new_n610), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n570), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n633));
  INV_X1    g208(.A(G91), .ZN(new_n634));
  OAI22_X1  g209(.A1(new_n633), .A2(new_n507), .B1(new_n634), .B2(new_n618), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n563), .B2(new_n565), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT85), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n632), .B1(new_n610), .B2(new_n637), .ZN(G297));
  AOI21_X1  g213(.A(new_n632), .B1(new_n610), .B2(new_n637), .ZN(G280));
  NOR2_X1   g214(.A1(new_n628), .A2(G559), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(G860), .B2(new_n629), .ZN(G148));
  NAND2_X1  g216(.A1(new_n552), .A2(new_n610), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n640), .B2(new_n610), .ZN(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g219(.A1(new_n482), .A2(G123), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n484), .A2(G135), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n461), .A2(G111), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n645), .B(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT86), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(G2096), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n464), .A2(new_n471), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT12), .Z(new_n653));
  XOR2_X1   g228(.A(KEYINPUT13), .B(G2100), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(new_n655), .ZN(G156));
  XNOR2_X1  g231(.A(G2427), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2430), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(KEYINPUT14), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT88), .ZN(new_n663));
  XOR2_X1   g238(.A(G1341), .B(G1348), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2451), .B(G2454), .Z(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n665), .B(new_n668), .Z(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n665), .B(new_n668), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(new_n670), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n674), .A3(G14), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G401));
  XOR2_X1   g251(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2084), .B(G2090), .Z(new_n679));
  XNOR2_X1  g254(.A(G2067), .B(G2678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(KEYINPUT17), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n678), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2072), .B(G2078), .Z(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n681), .B2(new_n677), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2096), .B(G2100), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1961), .B(G1966), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT90), .ZN(new_n693));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT91), .B(KEYINPUT20), .Z(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n693), .A2(new_n694), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n691), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n698), .A2(new_n695), .A3(new_n691), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n696), .B1(new_n695), .B2(new_n691), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT92), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n705), .B(new_n707), .Z(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n705), .B(new_n707), .ZN(new_n711));
  INV_X1    g286(.A(new_n709), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n710), .A2(new_n713), .ZN(G229));
  MUX2_X1   g289(.A(G6), .B(G305), .S(G16), .Z(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT32), .B(G1981), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G288), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G16), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G16), .B2(G23), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT33), .B(G1976), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT94), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n720), .A2(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G22), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G166), .B2(new_n725), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1971), .ZN(new_n728));
  NOR4_X1   g303(.A1(new_n717), .A2(new_n723), .A3(new_n724), .A4(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT34), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  MUX2_X1   g307(.A(G24), .B(G290), .S(G16), .Z(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(G1986), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(G1986), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n482), .A2(G119), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n484), .A2(G131), .ZN(new_n737));
  OR2_X1    g312(.A1(G95), .A2(G2105), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n738), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT93), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n736), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  MUX2_X1   g316(.A(G25), .B(new_n741), .S(G29), .Z(new_n742));
  XOR2_X1   g317(.A(KEYINPUT35), .B(G1991), .Z(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n742), .B(new_n744), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n734), .A2(new_n735), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n731), .A2(new_n732), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT36), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT95), .ZN(new_n749));
  OR3_X1    g324(.A1(new_n749), .A2(G4), .A3(G16), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(G4), .B2(G16), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n750), .B(new_n751), .C1(new_n628), .C2(new_n725), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1348), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT25), .Z(new_n755));
  AOI22_X1  g330(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(new_n461), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G139), .B2(new_n484), .ZN(new_n758));
  INV_X1    g333(.A(G29), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n759), .B2(G33), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(G2072), .ZN(new_n763));
  NOR2_X1   g338(.A1(G164), .A2(new_n759), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G27), .B2(new_n759), .ZN(new_n765));
  INV_X1    g340(.A(G2078), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n762), .A2(G2072), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n763), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT31), .B(G11), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT100), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT30), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n759), .B1(new_n773), .B2(G28), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n773), .B2(G28), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT24), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n759), .B1(new_n776), .B2(G34), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n776), .B2(G34), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G160), .B2(G29), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n772), .B(new_n775), .C1(new_n779), .C2(G2084), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n780), .B1(G2084), .B2(new_n779), .C1(new_n650), .C2(new_n759), .ZN(new_n781));
  NOR2_X1   g356(.A1(G16), .A2(G19), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n553), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1341), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n770), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G2090), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n759), .A2(G35), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT101), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G162), .B2(new_n759), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT29), .Z(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT27), .B(G1996), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n484), .A2(G141), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n464), .A2(G105), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(KEYINPUT97), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT97), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n464), .A2(new_n795), .A3(G105), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n479), .A2(G129), .A3(new_n480), .ZN(new_n799));
  NAND3_X1  g374(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT26), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(KEYINPUT98), .B1(new_n798), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  AOI22_X1  g379(.A1(G141), .A2(new_n484), .B1(new_n794), .B2(new_n796), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT98), .ZN(new_n806));
  INV_X1    g381(.A(new_n802), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n804), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G29), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G29), .B2(G32), .ZN(new_n812));
  OAI221_X1 g387(.A(new_n785), .B1(new_n786), .B2(new_n790), .C1(new_n791), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n791), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT99), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n790), .A2(new_n786), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(KEYINPUT102), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(KEYINPUT102), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n725), .A2(G20), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT23), .Z(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G299), .B2(G16), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1956), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n817), .A2(new_n818), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n759), .A2(G26), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT28), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n482), .A2(G128), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n484), .A2(G140), .ZN(new_n827));
  OR2_X1    g402(.A1(G104), .A2(G2105), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n828), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n825), .B1(new_n831), .B2(new_n759), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT96), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G2067), .ZN(new_n834));
  NOR2_X1   g409(.A1(G5), .A2(G16), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G171), .B2(G16), .ZN(new_n836));
  INV_X1    g411(.A(G1961), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(G16), .A2(G21), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G168), .B2(G16), .ZN(new_n840));
  INV_X1    g415(.A(G1966), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n834), .A2(new_n838), .A3(new_n842), .ZN(new_n843));
  NOR4_X1   g418(.A1(new_n813), .A2(new_n815), .A3(new_n823), .A4(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n748), .A2(new_n753), .A3(new_n844), .ZN(G150));
  INV_X1    g420(.A(G150), .ZN(G311));
  NAND2_X1  g421(.A1(new_n528), .A2(G55), .ZN(new_n847));
  NAND2_X1  g422(.A1(G80), .A2(G543), .ZN(new_n848));
  INV_X1    g423(.A(G67), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n512), .B2(new_n849), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n536), .A2(G93), .B1(G651), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G860), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT104), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT37), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n629), .A2(G559), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT38), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n552), .A2(new_n852), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n547), .A2(new_n847), .A3(new_n551), .A4(new_n851), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n857), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT103), .ZN(new_n864));
  INV_X1    g439(.A(G860), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n861), .B2(new_n862), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n855), .B1(new_n864), .B2(new_n866), .ZN(G145));
  INV_X1    g442(.A(G37), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n650), .B(G160), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n488), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT108), .B1(new_n803), .B2(new_n808), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT105), .B1(new_n493), .B2(new_n494), .ZN(new_n873));
  INV_X1    g448(.A(new_n494), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n875), .A3(new_n492), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n496), .A2(KEYINPUT106), .A3(new_n498), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT106), .B1(new_n496), .B2(new_n498), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n877), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n878), .B1(new_n877), .B2(new_n881), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n830), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n875), .B1(new_n874), .B2(new_n492), .ZN(new_n886));
  NOR3_X1   g461(.A1(new_n493), .A2(KEYINPUT105), .A3(new_n494), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n881), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT107), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n889), .A2(new_n831), .A3(new_n882), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n803), .A2(new_n808), .A3(KEYINPUT108), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n872), .A2(new_n885), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n831), .B1(new_n889), .B2(new_n882), .ZN(new_n893));
  INV_X1    g468(.A(new_n890), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n803), .A2(KEYINPUT108), .A3(new_n808), .ZN(new_n895));
  OAI22_X1  g470(.A1(new_n893), .A2(new_n894), .B1(new_n895), .B2(new_n871), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n892), .A2(new_n896), .A3(new_n758), .ZN(new_n897));
  INV_X1    g472(.A(new_n758), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n805), .A2(new_n807), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n885), .A2(new_n899), .A3(new_n890), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n885), .B2(new_n890), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT109), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n899), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n894), .B2(new_n893), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n900), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(KEYINPUT109), .A3(new_n898), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n897), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n741), .B(new_n653), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n484), .A2(G142), .ZN(new_n912));
  OR2_X1    g487(.A1(G106), .A2(G2105), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n913), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n915), .B1(G130), .B2(new_n482), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n911), .B(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n870), .B1(new_n910), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n917), .ZN(new_n919));
  AOI211_X1 g494(.A(new_n919), .B(new_n897), .C1(new_n905), .C2(new_n909), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n868), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n910), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n892), .A2(new_n896), .A3(new_n758), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT109), .B1(new_n908), .B2(new_n898), .ZN(new_n927));
  AOI211_X1 g502(.A(new_n904), .B(new_n758), .C1(new_n907), .C2(new_n900), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n926), .B(new_n924), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n869), .B(G162), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n925), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n922), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g510(.A1(new_n852), .A2(new_n610), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n640), .B(new_n860), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT111), .B1(new_n625), .B2(new_n636), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n939));
  NAND4_X1  g514(.A1(G299), .A2(new_n939), .A3(new_n615), .A4(new_n624), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n938), .A2(KEYINPUT112), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT112), .B1(new_n938), .B2(new_n940), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n625), .A2(new_n636), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n937), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n938), .A2(new_n940), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n938), .A2(new_n940), .A3(KEYINPUT112), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n943), .A2(KEYINPUT41), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n947), .A2(new_n943), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT41), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n946), .B1(new_n937), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n718), .B(G305), .ZN(new_n959));
  XNOR2_X1  g534(.A(G290), .B(G303), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n959), .B(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT42), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n958), .B(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n936), .B1(new_n963), .B2(new_n610), .ZN(G295));
  OAI21_X1  g539(.A(new_n936), .B1(new_n963), .B2(new_n610), .ZN(G331));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n967));
  OAI21_X1  g542(.A(G171), .B1(new_n577), .B2(new_n578), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n538), .A2(G301), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n860), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n860), .B1(new_n968), .B2(new_n969), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n941), .A2(new_n942), .A3(new_n951), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT41), .B1(new_n947), .B2(new_n943), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n967), .B(new_n973), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT113), .B1(new_n945), .B2(new_n973), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n968), .A2(new_n969), .ZN(new_n978));
  INV_X1    g553(.A(new_n860), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n970), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(new_n953), .B2(new_n956), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n976), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n961), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n983), .A2(KEYINPUT115), .A3(new_n984), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n984), .B1(new_n983), .B2(KEYINPUT114), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n949), .A2(new_n943), .A3(new_n950), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n967), .B1(new_n992), .B2(new_n981), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(new_n995), .A3(new_n976), .ZN(new_n996));
  AOI21_X1  g571(.A(G37), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n966), .B1(new_n989), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n973), .A2(new_n947), .A3(new_n952), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n992), .A2(new_n955), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n999), .B(new_n1000), .C1(new_n945), .C2(new_n973), .ZN(new_n1001));
  AOI21_X1  g576(.A(G37), .B1(new_n1001), .B2(new_n961), .ZN(new_n1002));
  AOI211_X1 g577(.A(new_n986), .B(new_n961), .C1(new_n994), .C2(new_n976), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT115), .B1(new_n983), .B2(new_n984), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n966), .B(new_n1002), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n998), .A2(new_n1006), .A3(KEYINPUT44), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n989), .A2(new_n997), .A3(new_n966), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1008), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT116), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT44), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n990), .A2(new_n996), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n868), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT43), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(new_n1008), .A3(new_n1005), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1015), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1013), .A2(new_n1022), .ZN(G397));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n889), .A2(new_n1024), .A3(new_n882), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G160), .A2(G40), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G2067), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n831), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n830), .A2(G2067), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1029), .B1(new_n1034), .B2(new_n899), .ZN(new_n1035));
  INV_X1    g610(.A(G1996), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1029), .A2(new_n1036), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1037), .A2(KEYINPUT46), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(KEYINPUT46), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1035), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g615(.A(new_n1040), .B(KEYINPUT47), .Z(new_n1041));
  NOR2_X1   g616(.A1(G290), .A2(G1986), .ZN(new_n1042));
  XOR2_X1   g617(.A(new_n1042), .B(KEYINPUT117), .Z(new_n1043));
  INV_X1    g618(.A(new_n1029), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(KEYINPUT48), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1045), .A2(KEYINPUT48), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n810), .A2(new_n1036), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n899), .A2(G1996), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n1033), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n741), .A2(new_n744), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n741), .A2(new_n744), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI211_X1 g629(.A(new_n1046), .B(new_n1047), .C1(new_n1029), .C2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1031), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n1041), .B(new_n1055), .C1(new_n1029), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1028), .ZN(new_n1058));
  NOR2_X1   g633(.A1(G164), .A2(G1384), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n888), .A2(new_n1024), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT118), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n888), .A2(new_n1064), .A3(new_n1024), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1061), .B1(new_n1066), .B2(new_n1060), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1028), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n1067), .A2(G1348), .B1(new_n1069), .B2(G2067), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1070), .A2(KEYINPUT60), .A3(new_n628), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1065), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1064), .B1(new_n888), .B2(new_n1024), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1060), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1061), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1348), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1077), .A2(new_n1078), .B1(new_n1030), .B2(new_n1068), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1072), .B1(new_n1079), .B2(new_n629), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1070), .A2(new_n628), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1071), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(G299), .B(KEYINPUT123), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT122), .B1(new_n563), .B2(new_n565), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(KEYINPUT57), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1083), .B(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n889), .A2(KEYINPUT45), .A3(new_n1024), .A4(new_n882), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1026), .B1(G164), .B2(G1384), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1058), .A3(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT56), .B(G2072), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1063), .A2(KEYINPUT50), .A3(new_n1065), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1028), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1095));
  AOI21_X1  g670(.A(G1956), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1087), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1083), .B(new_n1085), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1096), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT61), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1097), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .A4(KEYINPUT61), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n1069), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1088), .A2(new_n1036), .A3(new_n1058), .A4(new_n1089), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n552), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1109), .B(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1082), .A2(new_n1105), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1097), .A2(KEYINPUT125), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT124), .B1(new_n1079), .B2(new_n628), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT125), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1087), .B(new_n1115), .C1(new_n1096), .C2(new_n1093), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1070), .A2(new_n1117), .A3(new_n629), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1101), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1112), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT50), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1122), .A2(G2084), .A3(new_n1061), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1028), .B1(new_n1059), .B2(KEYINPUT45), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1066), .B2(KEYINPUT45), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1123), .A2(KEYINPUT120), .B1(new_n841), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1077), .B2(G2084), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1126), .A2(G168), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(G8), .ZN(new_n1130));
  AOI21_X1  g705(.A(G168), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT51), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT51), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1129), .A2(new_n1133), .A3(G8), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT49), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n598), .A2(new_n599), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(new_n593), .ZN(new_n1138));
  INV_X1    g713(.A(G1981), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1138), .A2(new_n1139), .A3(new_n595), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1138), .B2(new_n595), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1136), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1142), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1144), .A2(KEYINPUT49), .A3(new_n1140), .ZN(new_n1145));
  INV_X1    g720(.A(G8), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1068), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1143), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT119), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1143), .A2(new_n1145), .A3(new_n1147), .A4(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(G303), .A2(G8), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT55), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(G1971), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1156), .A2(new_n786), .B1(new_n1157), .B2(new_n1090), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1154), .B1(new_n1158), .B2(new_n1146), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1090), .A2(new_n1157), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n1077), .B2(G2090), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1154), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1161), .A2(G8), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT52), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n718), .A2(G1976), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1147), .B2(new_n1165), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1147), .A2(new_n1165), .ZN(new_n1167));
  INV_X1    g742(.A(G1976), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT52), .B1(G288), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1166), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1152), .A2(new_n1159), .A3(new_n1163), .A4(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1088), .A2(new_n766), .A3(new_n1058), .A4(new_n1089), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT53), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1173), .A2(G2078), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1124), .B(new_n1175), .C1(new_n1066), .C2(KEYINPUT45), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1174), .B(new_n1176), .C1(G1961), .C2(new_n1067), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT54), .B1(new_n1177), .B2(G171), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1077), .A2(new_n837), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1027), .A2(new_n1058), .A3(new_n1175), .A4(new_n1088), .ZN(new_n1180));
  AOI21_X1  g755(.A(G301), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1177), .A2(G171), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1179), .A2(G301), .A3(new_n1180), .ZN(new_n1184));
  AOI21_X1  g759(.A(KEYINPUT54), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1171), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1121), .A2(new_n1135), .A3(new_n1186), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1152), .A2(new_n1170), .A3(new_n1163), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1189));
  NOR2_X1   g764(.A1(G286), .A2(new_n1146), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1189), .A2(KEYINPUT63), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1161), .A2(G8), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1193), .A2(new_n1154), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1188), .A2(new_n1192), .A3(KEYINPUT121), .A4(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT63), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1196), .B1(new_n1171), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT121), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1194), .A2(new_n1189), .A3(KEYINPUT63), .A4(new_n1190), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1152), .A2(new_n1170), .A3(new_n1163), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1195), .A2(new_n1198), .A3(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1152), .A2(new_n1168), .A3(new_n718), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1140), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1163), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1152), .A2(new_n1170), .ZN(new_n1207));
  AOI22_X1  g782(.A1(new_n1205), .A2(new_n1147), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1187), .A2(new_n1203), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1132), .A2(new_n1210), .A3(new_n1134), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1171), .A2(new_n1183), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  OR2_X1    g788(.A1(new_n1213), .A2(KEYINPUT126), .ZN(new_n1214));
  AOI22_X1  g789(.A1(new_n1213), .A2(KEYINPUT126), .B1(KEYINPUT62), .B2(new_n1135), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1209), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1054), .B1(G1986), .B2(G290), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1044), .B1(new_n1217), .B2(new_n1043), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1057), .B1(new_n1216), .B2(new_n1218), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n1221));
  NAND2_X1  g795(.A1(new_n1019), .A2(new_n1005), .ZN(new_n1222));
  INV_X1    g796(.A(new_n459), .ZN(new_n1223));
  OR2_X1    g797(.A1(new_n1223), .A2(G227), .ZN(new_n1224));
  AOI21_X1  g798(.A(new_n1224), .B1(new_n710), .B2(new_n713), .ZN(new_n1225));
  AND2_X1   g799(.A1(new_n1225), .A2(new_n675), .ZN(new_n1226));
  OAI21_X1  g800(.A(new_n1226), .B1(new_n921), .B2(new_n932), .ZN(new_n1227));
  INV_X1    g801(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g802(.A(new_n1221), .B1(new_n1222), .B2(new_n1228), .ZN(new_n1229));
  AOI211_X1 g803(.A(KEYINPUT127), .B(new_n1227), .C1(new_n1019), .C2(new_n1005), .ZN(new_n1230));
  NOR2_X1   g804(.A1(new_n1229), .A2(new_n1230), .ZN(G308));
  NAND2_X1  g805(.A1(new_n1222), .A2(new_n1228), .ZN(G225));
endmodule


