//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n210), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(new_n215), .A2(new_n216), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n221), .B1(new_n215), .B2(new_n216), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n223), .B1(new_n202), .B2(new_n224), .C1(new_n203), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n212), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n222), .A2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n224), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n244), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(KEYINPUT77), .ZN(new_n250));
  AND2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G223), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n250), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G226), .A3(G1698), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G87), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n254), .A2(G223), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n264), .B(KEYINPUT77), .C1(new_n252), .C2(new_n251), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n256), .A2(new_n262), .A3(new_n263), .A4(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G179), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  INV_X1    g0070(.A(new_n217), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n274), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n276), .B1(new_n278), .B2(new_n224), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n268), .A2(new_n269), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT78), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n279), .B1(new_n266), .B2(new_n267), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(KEYINPUT78), .A3(new_n269), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n268), .A2(new_n280), .ZN(new_n286));
  INV_X1    g0086(.A(G169), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n283), .A2(new_n285), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT69), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n202), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n217), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(G1), .B2(new_n210), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n297), .B1(new_n294), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT16), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n259), .A2(new_n210), .A3(new_n260), .ZN(new_n304));
  AND2_X1   g0104(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n305));
  NOR2_X1   g0105(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n251), .A2(new_n252), .A3(G20), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n308), .A2(KEYINPUT76), .B1(KEYINPUT7), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT76), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n304), .A2(new_n311), .A3(new_n307), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n203), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n202), .A2(new_n203), .ZN(new_n314));
  NOR2_X1   g0114(.A1(G58), .A2(G68), .ZN(new_n315));
  OAI21_X1  g0115(.A(G20), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(G20), .A2(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G159), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n303), .B1(new_n313), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n309), .A2(new_n307), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n203), .B1(new_n304), .B2(KEYINPUT7), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n300), .B1(new_n323), .B2(KEYINPUT16), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n302), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT18), .B1(new_n289), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT76), .B1(new_n309), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n309), .A2(KEYINPUT7), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n312), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n319), .B1(new_n330), .B2(G68), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n324), .B1(new_n331), .B2(KEYINPUT16), .ZN(new_n332));
  INV_X1    g0132(.A(new_n302), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT18), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n281), .A2(new_n282), .B1(new_n286), .B2(new_n287), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .A4(new_n285), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n326), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT79), .ZN(new_n339));
  INV_X1    g0139(.A(G190), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n268), .A2(new_n340), .A3(new_n280), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(G200), .B2(new_n284), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(new_n332), .A3(new_n333), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT17), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT17), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n325), .A2(new_n345), .A3(new_n342), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(new_n346), .A3(KEYINPUT80), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT80), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n343), .A2(KEYINPUT17), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n345), .B1(new_n325), .B2(new_n342), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT79), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n326), .A2(new_n352), .A3(new_n337), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n339), .A2(new_n347), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT13), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n224), .A2(new_n254), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n261), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT72), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G97), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n261), .A2(G226), .A3(new_n254), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT72), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n261), .A2(new_n362), .A3(new_n357), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n359), .A2(new_n360), .A3(new_n361), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n267), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n276), .B1(new_n278), .B2(new_n225), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n356), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  AOI211_X1 g0168(.A(KEYINPUT13), .B(new_n366), .C1(new_n364), .C2(new_n267), .ZN(new_n369));
  OAI21_X1  g0169(.A(G200), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n363), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n362), .B1(new_n261), .B2(new_n357), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n361), .A2(new_n360), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n277), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT13), .B1(new_n375), .B2(new_n366), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n365), .A2(new_n356), .A3(new_n367), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(G190), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT12), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n295), .B2(G68), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n296), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(new_n381), .C1(new_n301), .C2(new_n203), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT73), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n383), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n317), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n258), .A2(G20), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G77), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n390), .A2(new_n299), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n391), .A2(KEYINPUT11), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(KEYINPUT11), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n384), .A2(new_n385), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n370), .A2(new_n378), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT14), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n398), .B(G169), .C1(new_n368), .C2(new_n369), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n376), .A2(G179), .A3(new_n377), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n287), .B1(new_n376), .B2(new_n377), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n402), .A2(KEYINPUT74), .A3(new_n398), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT74), .ZN(new_n404));
  OAI21_X1  g0204(.A(G169), .B1(new_n368), .B2(new_n369), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n404), .B1(new_n405), .B2(KEYINPUT14), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n401), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n397), .B1(new_n407), .B2(new_n394), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n254), .A2(G222), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G223), .A2(G1698), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n261), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n411), .B(new_n267), .C1(G77), .C2(new_n261), .ZN(new_n412));
  XOR2_X1   g0212(.A(KEYINPUT68), .B(G226), .Z(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(new_n276), .C1(new_n278), .C2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(new_n340), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(G200), .B2(new_n414), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n292), .A2(new_n387), .A3(new_n293), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n317), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n300), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n296), .A2(new_n201), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n301), .B2(new_n201), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT9), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n416), .A2(new_n424), .ZN(new_n425));
  OR2_X1    g0225(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n426));
  NAND2_X1  g0226(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n416), .A2(new_n424), .A3(KEYINPUT71), .A4(KEYINPUT10), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n414), .A2(G179), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n287), .B2(new_n414), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n419), .B2(new_n421), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT15), .B(G87), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT70), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n435), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n387), .ZN(new_n439));
  INV_X1    g0239(.A(new_n290), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n440), .A2(new_n317), .B1(G20), .B2(G77), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n300), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n296), .A2(new_n389), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n301), .B2(new_n389), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G238), .A2(G1698), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n261), .B(new_n446), .C1(new_n224), .C2(G1698), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n447), .B(new_n267), .C1(G107), .C2(new_n261), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n277), .A2(G244), .A3(new_n274), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n276), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G200), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n450), .A2(new_n340), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n445), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n287), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n448), .A2(new_n269), .A3(new_n276), .A4(new_n449), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n445), .A2(new_n457), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n433), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n355), .A2(new_n408), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT87), .ZN(new_n461));
  INV_X1    g0261(.A(G41), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n209), .B(G45), .C1(new_n462), .C2(KEYINPUT5), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT5), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G41), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n273), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n277), .B(G270), .C1(new_n463), .C2(new_n466), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(G264), .A2(G1698), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n261), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT86), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n261), .A2(G257), .A3(new_n254), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n253), .A2(G303), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n261), .A2(KEYINPUT86), .A3(new_n471), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n474), .A2(new_n475), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n470), .B1(new_n478), .B2(new_n267), .ZN(new_n479));
  INV_X1    g0279(.A(G116), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n296), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n209), .A2(G33), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n295), .A2(new_n482), .A3(new_n217), .A4(new_n298), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n483), .B2(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n210), .C1(G33), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n480), .A2(G20), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n487), .A2(new_n488), .A3(new_n299), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT20), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n490), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n484), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n479), .A2(new_n287), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n461), .B1(new_n494), .B2(KEYINPUT21), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n478), .A2(new_n267), .ZN(new_n496));
  INV_X1    g0296(.A(new_n470), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n493), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(G169), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT21), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(KEYINPUT87), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n498), .A2(KEYINPUT21), .A3(new_n499), .A4(G169), .ZN(new_n504));
  AOI211_X1 g0304(.A(new_n269), .B(new_n470), .C1(new_n478), .C2(new_n267), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n499), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n499), .B1(new_n498), .B2(G200), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n340), .B2(new_n498), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n503), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT82), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n209), .A2(G45), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G250), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n512), .B1(new_n267), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n513), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n273), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G244), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G1698), .ZN(new_n520));
  OAI221_X1 g0320(.A(new_n520), .B1(G238), .B2(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G116), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n267), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n277), .A2(KEYINPUT82), .A3(G250), .A4(new_n513), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n518), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n287), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n515), .A2(new_n517), .A3(new_n525), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n277), .B1(new_n521), .B2(new_n522), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n269), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n295), .B1(new_n436), .B2(new_n437), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n360), .A2(new_n210), .ZN(new_n534));
  AND2_X1   g0334(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n535));
  NOR2_X1   g0335(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n536));
  INV_X1    g0336(.A(G87), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n486), .ZN(new_n538));
  OAI221_X1 g0338(.A(new_n534), .B1(new_n535), .B2(new_n536), .C1(G107), .C2(new_n538), .ZN(new_n539));
  XOR2_X1   g0339(.A(KEYINPUT83), .B(KEYINPUT19), .Z(new_n540));
  NAND2_X1  g0340(.A1(new_n387), .A2(G97), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT84), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n261), .A2(new_n544), .A3(new_n210), .A4(G68), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n261), .A2(new_n210), .A3(G68), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT84), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n533), .B1(new_n548), .B2(new_n300), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT85), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n436), .A2(new_n437), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(new_n483), .ZN(new_n552));
  INV_X1    g0352(.A(new_n483), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n436), .A2(new_n553), .A3(KEYINPUT85), .A4(new_n437), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n527), .B(new_n531), .C1(new_n549), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n547), .A2(new_n545), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n539), .A2(new_n542), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n532), .B1(new_n559), .B2(new_n299), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n526), .A2(G200), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n553), .A2(G87), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n530), .A2(G190), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n560), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n556), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n261), .A2(G257), .A3(G1698), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n261), .A2(G250), .A3(new_n254), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G294), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n267), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n267), .B1(new_n464), .B2(new_n467), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G264), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n468), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G169), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n569), .A2(new_n267), .B1(new_n571), .B2(G264), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(G179), .A3(new_n468), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n210), .B(G87), .C1(new_n251), .C2(new_n252), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT22), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT22), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n261), .A2(new_n580), .A3(new_n210), .A4(G87), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g0382(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT89), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n522), .B2(G20), .ZN(new_n585));
  OR3_X1    g0385(.A1(new_n210), .A2(KEYINPUT23), .A3(G107), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n210), .A2(KEYINPUT89), .A3(G33), .A4(G116), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT23), .B1(new_n210), .B2(G107), .ZN(new_n588));
  AND4_X1   g0388(.A1(new_n585), .A2(new_n586), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n582), .A2(new_n583), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n583), .B1(new_n582), .B2(new_n589), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n299), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT25), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n295), .B2(G107), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n295), .A2(new_n593), .A3(G107), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n594), .A2(new_n596), .B1(new_n553), .B2(G107), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n577), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n573), .A2(G190), .ZN(new_n600));
  AOI21_X1  g0400(.A(G200), .B1(new_n575), .B2(new_n468), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n592), .B(new_n597), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(G107), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n310), .B2(new_n312), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n317), .A2(G77), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT6), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n606), .A2(new_n486), .A3(G107), .ZN(new_n607));
  XNOR2_X1  g0407(.A(G97), .B(G107), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n607), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n605), .B1(new_n609), .B2(new_n210), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n299), .B1(new_n604), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n295), .A2(G97), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n553), .B2(G97), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n277), .B(G257), .C1(new_n463), .C2(new_n466), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n468), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n254), .A2(G244), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n261), .B(new_n617), .C1(KEYINPUT81), .C2(KEYINPUT4), .ZN(new_n618));
  NOR2_X1   g0418(.A1(KEYINPUT81), .A2(KEYINPUT4), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n253), .B2(new_n616), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n618), .A2(new_n620), .A3(new_n485), .A4(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n615), .B1(new_n622), .B2(new_n267), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n623), .A2(G200), .ZN(new_n624));
  AOI211_X1 g0424(.A(G190), .B(new_n615), .C1(new_n622), .C2(new_n267), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n611), .B(new_n613), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n610), .B1(new_n330), .B2(G107), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n613), .B1(new_n627), .B2(new_n300), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n623), .A2(new_n269), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n622), .A2(new_n267), .ZN(new_n630));
  INV_X1    g0430(.A(new_n615), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n287), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n628), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n599), .A2(new_n602), .A3(new_n626), .A4(new_n634), .ZN(new_n635));
  NOR4_X1   g0435(.A1(new_n460), .A2(new_n511), .A3(new_n565), .A4(new_n635), .ZN(G372));
  INV_X1    g0436(.A(new_n432), .ZN(new_n637));
  INV_X1    g0437(.A(new_n338), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n344), .A2(KEYINPUT80), .A3(new_n346), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT80), .B1(new_n344), .B2(new_n346), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n407), .A2(new_n394), .B1(new_n396), .B2(new_n458), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n638), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n428), .A2(new_n429), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n637), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT26), .B1(new_n565), .B2(new_n634), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n628), .A2(new_n633), .A3(new_n629), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n518), .A2(KEYINPUT90), .A3(new_n525), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT90), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n529), .B1(new_n528), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n287), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n653), .B(new_n531), .C1(new_n549), .C2(new_n555), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n652), .A2(G200), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n656), .A2(new_n560), .A3(new_n562), .A4(new_n563), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n648), .A2(new_n654), .A3(new_n655), .A4(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n647), .A2(new_n658), .A3(new_n654), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n577), .A2(new_n598), .A3(KEYINPUT91), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT91), .B1(new_n577), .B2(new_n598), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n503), .B(new_n508), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n602), .A2(new_n626), .A3(new_n634), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n531), .B1(new_n549), .B2(new_n555), .ZN(new_n664));
  INV_X1    g0464(.A(new_n653), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n666));
  INV_X1    g0466(.A(G200), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(new_n649), .B2(new_n651), .ZN(new_n668));
  OAI22_X1  g0468(.A1(new_n664), .A2(new_n665), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n659), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n646), .B1(new_n460), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT92), .ZN(G369));
  INV_X1    g0475(.A(G330), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n511), .B(KEYINPUT93), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n677), .B1(new_n493), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n507), .B1(new_n495), .B2(new_n502), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(new_n499), .A3(new_n683), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n676), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT94), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n599), .B2(new_n684), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n598), .A2(new_n683), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n599), .A2(new_n692), .A3(new_n602), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n577), .A2(new_n598), .A3(KEYINPUT94), .A4(new_n683), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n686), .A2(new_n683), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n695), .ZN(new_n698));
  OR3_X1    g0498(.A1(new_n660), .A2(new_n661), .A3(new_n683), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n696), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n213), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n538), .A2(G107), .A3(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n219), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT95), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n503), .A2(new_n508), .A3(new_n599), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n670), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT26), .B1(new_n669), .B2(new_n634), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n648), .A2(new_n655), .A3(new_n556), .A4(new_n564), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(new_n654), .A3(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(KEYINPUT29), .B(new_n684), .C1(new_n712), .C2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n683), .B1(new_n659), .B2(new_n671), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(KEYINPUT29), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n635), .A2(new_n565), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n719), .A2(new_n686), .A3(new_n510), .A4(new_n684), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n479), .A2(G179), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(new_n573), .A3(new_n632), .A4(new_n652), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n479), .A2(G179), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n623), .A2(new_n530), .A3(new_n575), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n575), .A2(new_n530), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(new_n505), .A3(KEYINPUT30), .A4(new_n623), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n722), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT31), .B1(new_n729), .B2(new_n683), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n676), .B1(new_n720), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n718), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n710), .B1(new_n735), .B2(G1), .ZN(G364));
  AND2_X1   g0536(.A1(new_n210), .A2(G13), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G45), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n705), .A2(G1), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n689), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n685), .A2(new_n676), .A3(new_n688), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n685), .A2(new_n688), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n210), .A2(G190), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G179), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G159), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT32), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n210), .A2(new_n340), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n667), .A2(G179), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n537), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n748), .A2(new_n755), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n757), .B1(G107), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n269), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n748), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n760), .B(new_n261), .C1(new_n389), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n754), .A2(new_n761), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT97), .Z(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n753), .B(new_n763), .C1(G58), .C2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n210), .B1(new_n749), .B2(G190), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n486), .ZN(new_n769));
  NAND3_X1  g0569(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n340), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n201), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n770), .A2(G190), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n769), .B(new_n773), .C1(G68), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G303), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n776), .A2(new_n756), .B1(new_n764), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G283), .ZN(new_n779));
  INV_X1    g0579(.A(new_n774), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT33), .B(G317), .Z(new_n781));
  OAI221_X1 g0581(.A(new_n253), .B1(new_n758), .B2(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n778), .B(new_n782), .C1(G329), .C2(new_n751), .ZN(new_n783));
  INV_X1    g0583(.A(new_n762), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n784), .A2(G311), .B1(G326), .B2(new_n771), .ZN(new_n785));
  INV_X1    g0585(.A(G294), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n786), .B2(new_n768), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT98), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n767), .A2(new_n775), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n217), .B1(G20), .B2(new_n287), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n740), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n746), .A2(new_n790), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n248), .A2(G45), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT96), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n703), .A2(new_n261), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n795), .B(new_n796), .C1(G45), .C2(new_n219), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n703), .A2(new_n253), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n798), .A2(G355), .B1(new_n480), .B2(new_n703), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n792), .B1(new_n793), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n747), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n743), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(G396));
  NAND2_X1  g0604(.A1(new_n458), .A2(KEYINPUT99), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT99), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n445), .B2(new_n457), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n454), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n672), .A2(new_n684), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n683), .B1(new_n442), .B2(new_n444), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n805), .A2(new_n453), .A3(new_n811), .A4(new_n807), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n458), .A2(new_n683), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n810), .B1(new_n717), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n740), .B1(new_n815), .B2(new_n734), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n734), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n790), .A2(new_n744), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n740), .B1(G77), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n764), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n261), .B(new_n769), .C1(G294), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n758), .A2(new_n537), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G311), .B2(new_n751), .ZN(new_n824));
  INV_X1    g0624(.A(new_n756), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G107), .A2(new_n825), .B1(new_n784), .B2(G116), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G283), .A2(new_n774), .B1(new_n771), .B2(G303), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n822), .A2(new_n824), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n784), .A2(G159), .B1(G150), .B2(new_n774), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  INV_X1    g0630(.A(G143), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(new_n830), .B2(new_n772), .C1(new_n765), .C2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n261), .B1(new_n756), .B2(new_n201), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n759), .A2(G68), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n837), .B2(new_n750), .ZN(new_n838));
  INV_X1    g0638(.A(new_n768), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n835), .B(new_n838), .C1(G58), .C2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n832), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n828), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n820), .B1(new_n843), .B2(new_n790), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n814), .B2(new_n745), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n817), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G384));
  INV_X1    g0647(.A(new_n609), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n848), .A2(KEYINPUT35), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(KEYINPUT35), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n849), .A2(G116), .A3(new_n218), .A4(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT36), .Z(new_n852));
  OAI211_X1 g0652(.A(new_n220), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n201), .A2(G68), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n209), .B(G13), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NOR4_X1   g0656(.A1(new_n511), .A2(new_n635), .A3(new_n565), .A4(new_n683), .ZN(new_n857));
  INV_X1    g0657(.A(new_n731), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n814), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n399), .A2(new_n400), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT74), .B1(new_n402), .B2(new_n398), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n405), .A2(new_n404), .A3(KEYINPUT14), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n394), .A2(new_n683), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n408), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(G58), .B(G68), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n870), .A2(G20), .B1(G159), .B2(new_n317), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT7), .ZN(new_n872));
  OAI21_X1  g0672(.A(G68), .B1(new_n309), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n304), .A2(new_n327), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n299), .B1(new_n875), .B2(new_n303), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n323), .A2(KEYINPUT16), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n333), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n681), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n354), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n878), .A2(new_n283), .A3(new_n285), .A4(new_n288), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(new_n343), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n334), .A2(new_n285), .A3(new_n336), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n334), .A2(new_n879), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .A4(new_n343), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n882), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n893), .B(new_n890), .C1(new_n354), .C2(new_n881), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n869), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT40), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n349), .A2(new_n350), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n334), .B(new_n879), .C1(new_n898), .C2(new_n338), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n886), .A2(new_n343), .A3(new_n887), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n889), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT38), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n890), .B1(new_n354), .B2(new_n881), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(new_n904), .B2(KEYINPUT38), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n720), .A2(new_n732), .B1(new_n813), .B2(new_n812), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n396), .B(new_n866), .C1(new_n865), .C2(new_n395), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n407), .A2(new_n394), .A3(new_n683), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n906), .A2(KEYINPUT40), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n897), .B1(new_n905), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n857), .A2(new_n860), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n460), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n913), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(G330), .A3(new_n915), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n865), .A2(new_n395), .A3(new_n683), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n326), .A2(new_n352), .A3(new_n337), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n352), .B1(new_n326), .B2(new_n337), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n880), .B1(new_n921), .B2(new_n641), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n893), .B1(new_n922), .B2(new_n890), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n882), .A2(KEYINPUT38), .A3(new_n891), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n894), .A2(KEYINPUT39), .A3(new_n903), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n917), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n808), .A2(new_n684), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT100), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n808), .A2(KEYINPUT100), .A3(new_n684), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n717), .B2(new_n809), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n933), .A2(new_n868), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n923), .A2(new_n924), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n934), .A2(new_n935), .B1(new_n338), .B2(new_n681), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n927), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n646), .B1(new_n718), .B2(new_n460), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n916), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n209), .B2(new_n737), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n916), .A2(new_n939), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n856), .B1(new_n941), .B2(new_n942), .ZN(G367));
  NAND2_X1  g0743(.A1(new_n438), .A2(new_n703), .ZN(new_n944));
  INV_X1    g0744(.A(new_n793), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n796), .B2(new_n239), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n739), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n758), .A2(new_n389), .B1(new_n750), .B2(new_n830), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n261), .B1(new_n768), .B2(new_n203), .C1(new_n201), .C2(new_n762), .ZN(new_n949));
  INV_X1    g0749(.A(G159), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n780), .A2(new_n950), .B1(new_n772), .B2(new_n831), .ZN(new_n951));
  INV_X1    g0751(.A(G150), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n202), .A2(new_n756), .B1(new_n764), .B2(new_n952), .ZN(new_n953));
  OR4_X1    g0753(.A1(new_n948), .A2(new_n949), .A3(new_n951), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n766), .A2(G303), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n756), .A2(new_n480), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(KEYINPUT46), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(G294), .B2(new_n774), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n839), .A2(G107), .B1(G311), .B2(new_n771), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n956), .A2(KEYINPUT46), .B1(new_n784), .B2(G283), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n955), .A2(new_n958), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(G317), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n253), .B1(new_n750), .B2(new_n962), .C1(new_n486), .C2(new_n758), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT105), .Z(new_n964));
  OAI21_X1  g0764(.A(new_n954), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT47), .Z(new_n966));
  AOI21_X1  g0766(.A(new_n684), .B1(new_n560), .B2(new_n562), .ZN(new_n967));
  MUX2_X1   g0767(.A(new_n669), .B(new_n654), .S(new_n967), .Z(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT101), .Z(new_n969));
  INV_X1    g0769(.A(new_n746), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n947), .B1(new_n791), .B2(new_n966), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n738), .A2(G1), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n697), .B(new_n695), .Z(new_n973));
  OR2_X1    g0773(.A1(new_n689), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n689), .A2(new_n973), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n974), .A2(new_n735), .A3(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT104), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n648), .A2(new_n683), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n628), .A2(new_n683), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n626), .A2(new_n634), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT44), .B1(new_n700), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n700), .A2(KEYINPUT44), .A3(new_n982), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n984), .A2(KEYINPUT103), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n701), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT45), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n700), .B2(new_n982), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT103), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n983), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n977), .B1(new_n987), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n976), .B1(new_n995), .B2(new_n696), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n696), .B2(new_n995), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n735), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n704), .B(KEYINPUT41), .Z(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n972), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n697), .A2(new_n695), .A3(new_n981), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(KEYINPUT42), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n980), .A2(new_n599), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n683), .B1(new_n1004), .B2(new_n634), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n1002), .B2(KEYINPUT42), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n969), .A2(KEYINPUT43), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  OR3_X1    g0808(.A1(new_n696), .A2(KEYINPUT102), .A3(new_n982), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(KEYINPUT102), .B1(new_n696), .B2(new_n982), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1011), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1008), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1015), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1017), .A2(new_n1007), .A3(new_n1013), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n971), .B1(new_n1001), .B2(new_n1019), .ZN(G387));
  AND2_X1   g0820(.A1(new_n974), .A2(new_n975), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n972), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT106), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n976), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1024), .A2(new_n705), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n735), .B2(new_n1021), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n798), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n1027), .A2(new_n706), .B1(G107), .B2(new_n213), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT107), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n440), .A2(new_n201), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT50), .ZN(new_n1031));
  AOI21_X1  g0831(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n706), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n796), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT108), .Z(new_n1035));
  NAND2_X1  g0835(.A1(new_n236), .A2(G45), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1029), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n740), .B1(new_n1037), .B2(new_n945), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n784), .A2(G303), .B1(G311), .B2(new_n774), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n777), .B2(new_n772), .C1(new_n765), .C2(new_n962), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n825), .A2(G294), .B1(new_n839), .B2(G283), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT49), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n758), .A2(new_n480), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n261), .B(new_n1049), .C1(G326), .C2(new_n751), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n551), .A2(new_n768), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n294), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1052), .B1(new_n1053), .B2(new_n774), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n261), .B1(new_n758), .B2(new_n486), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n764), .A2(new_n201), .B1(new_n762), .B2(new_n203), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(G159), .C2(new_n771), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n756), .A2(new_n389), .B1(new_n750), .B2(new_n952), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT109), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1054), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1051), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1038), .B1(new_n1061), .B2(new_n790), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n695), .B2(new_n970), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1023), .A2(new_n1026), .A3(new_n1063), .ZN(G393));
  OAI211_X1 g0864(.A(new_n689), .B(new_n695), .C1(new_n987), .C2(new_n994), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(KEYINPUT110), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n991), .A2(new_n696), .A3(new_n986), .A4(new_n993), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1065), .A2(KEYINPUT110), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n976), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(new_n704), .A3(new_n997), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(KEYINPUT113), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT113), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1070), .A2(new_n1073), .A3(new_n704), .A4(new_n997), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1069), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1075), .A2(new_n972), .A3(new_n1067), .A4(new_n1066), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n244), .A2(new_n703), .A3(new_n261), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n793), .B1(new_n486), .B2(new_n213), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n740), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n821), .A2(G311), .B1(G317), .B2(new_n771), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n1081));
  XNOR2_X1  g0881(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n756), .A2(new_n779), .B1(new_n762), .B2(new_n786), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G322), .B2(new_n751), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n253), .B1(new_n758), .B2(new_n603), .C1(new_n780), .C2(new_n776), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G116), .B2(new_n839), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1082), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n784), .A2(new_n440), .B1(G50), .B2(new_n774), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1089), .A2(KEYINPUT111), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(KEYINPUT111), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n756), .A2(new_n203), .B1(new_n750), .B2(new_n831), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n768), .A2(new_n389), .ZN(new_n1093));
  NOR4_X1   g0893(.A1(new_n1092), .A2(new_n823), .A3(new_n1093), .A4(new_n253), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1090), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n821), .A2(G159), .B1(G150), .B2(new_n771), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT51), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1087), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1079), .B1(new_n790), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n981), .B2(new_n970), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1076), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1072), .A2(new_n1074), .A3(new_n1102), .ZN(G390));
  OAI21_X1  g0903(.A(KEYINPUT39), .B1(new_n892), .B2(new_n894), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n905), .A2(new_n918), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n407), .A2(new_n394), .A3(new_n684), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n933), .B2(new_n868), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT116), .ZN(new_n1109));
  AND4_X1   g0909(.A1(new_n1109), .A2(new_n733), .A3(new_n814), .A4(new_n909), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n917), .A2(KEYINPUT114), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT114), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1106), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n903), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1114), .B1(new_n924), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n684), .B(new_n809), .C1(new_n712), .C2(new_n715), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n930), .A2(new_n931), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n909), .A2(KEYINPUT115), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT115), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n907), .B2(new_n908), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1119), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1110), .B1(new_n1116), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n733), .A2(new_n909), .A3(new_n814), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT116), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1108), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1126), .B1(new_n1108), .B2(new_n1124), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n733), .A2(new_n355), .A3(new_n408), .A4(new_n459), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n646), .B(new_n1131), .C1(new_n718), .C2(new_n460), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n868), .A2(new_n1121), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n733), .A2(new_n814), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1122), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1136), .A2(new_n1118), .A3(new_n1125), .A4(new_n1117), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n810), .A2(new_n1118), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1125), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n909), .B1(new_n733), .B2(new_n814), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1132), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1128), .A2(new_n1130), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1142), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1144), .A2(new_n704), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(G125), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n758), .A2(new_n201), .B1(new_n750), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n825), .A2(G150), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT53), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT54), .B(G143), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1148), .B(new_n1150), .C1(new_n784), .C2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n780), .A2(new_n830), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n261), .B1(new_n768), .B2(new_n950), .C1(new_n837), .C2(new_n764), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(G128), .C2(new_n771), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n772), .A2(new_n779), .B1(new_n762), .B2(new_n486), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G107), .B2(new_n774), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT117), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n836), .B1(new_n480), .B2(new_n764), .C1(new_n786), .C2(new_n750), .ZN(new_n1160));
  NOR4_X1   g0960(.A1(new_n1160), .A2(new_n261), .A3(new_n757), .A4(new_n1093), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1153), .A2(new_n1156), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n740), .B1(new_n1053), .B2(new_n819), .C1(new_n1162), .C2(new_n791), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1163), .B1(new_n1165), .B2(new_n744), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1166), .B1(new_n1167), .B2(new_n972), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1146), .A2(new_n1168), .ZN(G378));
  OAI22_X1  g0969(.A1(new_n772), .A2(new_n1147), .B1(new_n768), .B2(new_n952), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G128), .A2(new_n821), .B1(new_n825), .B2(new_n1152), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n830), .B2(new_n762), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(G132), .C2(new_n774), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n759), .A2(G159), .ZN(new_n1177));
  AOI211_X1 g0977(.A(G33), .B(G41), .C1(new_n751), .C2(G124), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n253), .A2(new_n462), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G77), .B2(new_n825), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n202), .B2(new_n758), .C1(new_n779), .C2(new_n750), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT118), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n764), .A2(new_n603), .B1(new_n768), .B2(new_n203), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n780), .A2(new_n486), .B1(new_n772), .B2(new_n480), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(new_n438), .C2(new_n784), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(KEYINPUT58), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1180), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1187), .A2(KEYINPUT58), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1179), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n790), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n739), .B1(new_n201), .B2(new_n818), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n433), .B(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n422), .A2(new_n681), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1195), .B(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1192), .B(new_n1193), .C1(new_n1198), .C2(new_n745), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1106), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n892), .A2(new_n894), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1138), .A2(new_n909), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1201), .A2(new_n1202), .B1(new_n638), .B2(new_n879), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT40), .B1(new_n935), .B2(new_n869), .ZN(new_n1205));
  OAI21_X1  g1005(.A(G330), .B1(new_n905), .B2(new_n910), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1205), .A2(new_n1206), .A3(new_n1198), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n924), .A2(new_n1115), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n906), .A2(KEYINPUT40), .A3(new_n909), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n676), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1197), .B1(new_n897), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1204), .B1(new_n1207), .B2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n897), .A2(new_n1210), .A3(new_n1197), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1198), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n937), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(KEYINPUT119), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT119), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1204), .B(new_n1217), .C1(new_n1207), .C2(new_n1211), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n972), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1199), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1132), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1145), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1212), .A2(KEYINPUT120), .A3(new_n1215), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT120), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n937), .A2(new_n1214), .A3(new_n1225), .A4(new_n1213), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(KEYINPUT57), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT57), .B1(new_n1145), .B2(new_n1222), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(new_n1218), .A3(new_n1216), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1221), .B1(new_n1231), .B2(new_n704), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(G375));
  NAND2_X1  g1033(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n972), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1133), .A2(new_n744), .A3(new_n1135), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n765), .A2(new_n830), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n253), .B1(new_n759), .B2(G58), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n201), .B2(new_n768), .C1(new_n780), .C2(new_n1151), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(G150), .A2(new_n784), .B1(new_n751), .B2(G128), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n950), .B2(new_n756), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n771), .A2(G132), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT121), .ZN(new_n1243));
  NOR4_X1   g1043(.A1(new_n1237), .A2(new_n1239), .A3(new_n1241), .A4(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n261), .B1(new_n759), .B2(G77), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1245), .B1(new_n772), .B2(new_n786), .C1(new_n480), .C2(new_n780), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n756), .A2(new_n486), .B1(new_n750), .B2(new_n776), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n764), .A2(new_n779), .B1(new_n762), .B2(new_n603), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1246), .A2(new_n1052), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n790), .B1(new_n1244), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n739), .B1(new_n203), .B2(new_n818), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1236), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1235), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1137), .A2(new_n1141), .A3(new_n1132), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1143), .A2(new_n1000), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(G381));
  NOR3_X1   g1057(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1258), .B(KEYINPUT122), .Z(new_n1259));
  NOR3_X1   g1059(.A1(new_n1259), .A2(G378), .A3(G381), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(G390), .A2(G387), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1232), .A3(new_n1261), .ZN(G407));
  INV_X1    g1062(.A(G378), .ZN(new_n1263));
  INV_X1    g1063(.A(G213), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1264), .A2(G343), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1232), .A2(new_n1263), .A3(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(G407), .A2(G213), .A3(new_n1266), .ZN(G409));
  INV_X1    g1067(.A(new_n1265), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT60), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1255), .B1(new_n1142), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n704), .B1(new_n1255), .B2(new_n1269), .ZN(new_n1272));
  OAI21_X1  g1072(.A(KEYINPUT124), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1272), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT124), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1270), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1277), .B2(new_n1254), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n846), .B(new_n1253), .C1(new_n1273), .C2(new_n1276), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n705), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1281), .A2(new_n1263), .A3(new_n1221), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(KEYINPUT123), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT123), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1224), .A2(new_n1285), .A3(new_n1226), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1284), .A2(new_n972), .A3(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1199), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n999), .B1(new_n1145), .B2(new_n1222), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1288), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G378), .B1(new_n1287), .B2(new_n1291), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1268), .B(new_n1280), .C1(new_n1282), .C2(new_n1292), .ZN(new_n1293));
  XOR2_X1   g1093(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1277), .A2(new_n1254), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n846), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1277), .A2(G384), .A3(new_n1254), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1265), .A2(G2897), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1298), .A2(new_n1299), .A3(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1300), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1292), .B1(new_n1232), .B2(G378), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1304), .B1(new_n1305), .B2(new_n1265), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1287), .A2(new_n1291), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1263), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1221), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1229), .A2(new_n1289), .B1(new_n1227), .B2(KEYINPUT57), .ZN(new_n1310));
  OAI211_X1 g1110(.A(G378), .B(new_n1309), .C1(new_n1310), .C2(new_n705), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT62), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1312), .A2(new_n1313), .A3(new_n1268), .A4(new_n1280), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1295), .A2(new_n1296), .A3(new_n1306), .A4(new_n1314), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(G393), .B(G396), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1101), .B1(new_n1071), .B2(KEYINPUT113), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n999), .B1(new_n997), .B2(new_n735), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1018), .B(new_n1016), .C1(new_n1319), .C2(new_n972), .ZN(new_n1320));
  AOI22_X1  g1120(.A1(new_n1318), .A2(new_n1074), .B1(new_n1320), .B2(new_n971), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1317), .B1(new_n1261), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(G390), .A2(G387), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1318), .A2(new_n1320), .A3(new_n971), .A4(new_n1074), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1323), .A2(new_n1324), .A3(new_n1316), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1322), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1315), .A2(new_n1326), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(KEYINPUT61), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT63), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1293), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT125), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1304), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1302), .A2(new_n1303), .A3(KEYINPUT125), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1332), .B(new_n1333), .C1(new_n1305), .C2(new_n1265), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1312), .A2(KEYINPUT63), .A3(new_n1268), .A4(new_n1280), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1328), .A2(new_n1330), .A3(new_n1334), .A4(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1327), .A2(new_n1336), .ZN(G405));
  NAND2_X1  g1137(.A1(new_n1280), .A2(KEYINPUT127), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1323), .A2(new_n1324), .A3(new_n1316), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1316), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1339), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1322), .A2(new_n1325), .A3(new_n1338), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1280), .A2(KEYINPUT127), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(G375), .A2(new_n1263), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1345), .B1(new_n1346), .B2(new_n1311), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(new_n1344), .B(new_n1347), .ZN(G402));
endmodule


