

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755;

  AND2_X1 U369 ( .A1(n598), .A2(n597), .ZN(n600) );
  INV_X1 U370 ( .A(G953), .ZN(n741) );
  XNOR2_X1 U371 ( .A(n347), .B(KEYINPUT36), .ZN(n585) );
  NOR2_X2 U372 ( .A1(n582), .A2(n583), .ZN(n347) );
  XNOR2_X2 U373 ( .A(n375), .B(KEYINPUT73), .ZN(n700) );
  XNOR2_X1 U374 ( .A(G104), .B(G101), .ZN(n438) );
  XNOR2_X1 U375 ( .A(n438), .B(n437), .ZN(n725) );
  NOR2_X2 U376 ( .A1(n739), .A2(n373), .ZN(n372) );
  INV_X1 U377 ( .A(n659), .ZN(n655) );
  XNOR2_X2 U378 ( .A(n550), .B(n551), .ZN(n701) );
  XNOR2_X2 U379 ( .A(n601), .B(KEYINPUT40), .ZN(n755) );
  NOR2_X2 U380 ( .A1(n755), .A2(n751), .ZN(n607) );
  INV_X1 U381 ( .A(G143), .ZN(n406) );
  XNOR2_X1 U382 ( .A(n406), .B(G128), .ZN(n506) );
  XNOR2_X1 U383 ( .A(KEYINPUT4), .B(KEYINPUT66), .ZN(n408) );
  XNOR2_X1 U384 ( .A(n370), .B(KEYINPUT32), .ZN(n547) );
  XNOR2_X1 U385 ( .A(n603), .B(KEYINPUT41), .ZN(n702) );
  NOR2_X1 U386 ( .A1(n575), .A2(n574), .ZN(n604) );
  XNOR2_X1 U387 ( .A(n666), .B(n385), .ZN(n588) );
  NOR2_X1 U388 ( .A1(n483), .A2(n523), .ZN(n596) );
  XNOR2_X1 U389 ( .A(n390), .B(KEYINPUT67), .ZN(n580) );
  XNOR2_X1 U390 ( .A(n541), .B(n522), .ZN(n549) );
  BUF_X1 U391 ( .A(n541), .Z(n542) );
  XNOR2_X1 U392 ( .A(n502), .B(n501), .ZN(n535) );
  NOR2_X2 U393 ( .A1(n620), .A2(G902), .ZN(n474) );
  XNOR2_X1 U394 ( .A(n387), .B(n386), .ZN(n718) );
  XNOR2_X1 U395 ( .A(n408), .B(n441), .ZN(n509) );
  XNOR2_X2 U396 ( .A(n738), .B(G146), .ZN(n471) );
  XNOR2_X2 U397 ( .A(n407), .B(n488), .ZN(n738) );
  NAND2_X1 U398 ( .A1(n680), .A2(n391), .ZN(n390) );
  NOR2_X1 U399 ( .A1(n523), .A2(n679), .ZN(n391) );
  INV_X1 U400 ( .A(n730), .ZN(n374) );
  AND2_X1 U401 ( .A1(n588), .A2(n384), .ZN(n589) );
  INV_X1 U402 ( .A(KEYINPUT47), .ZN(n384) );
  NOR2_X1 U403 ( .A1(KEYINPUT17), .A2(G953), .ZN(n398) );
  XNOR2_X1 U404 ( .A(n509), .B(n442), .ZN(n407) );
  INV_X1 U405 ( .A(G137), .ZN(n442) );
  XNOR2_X1 U406 ( .A(n365), .B(n364), .ZN(n363) );
  INV_X1 U407 ( .A(KEYINPUT104), .ZN(n364) );
  NAND2_X1 U408 ( .A1(n564), .A2(n588), .ZN(n365) );
  NAND2_X1 U409 ( .A1(n661), .A2(n647), .ZN(n564) );
  INV_X1 U410 ( .A(KEYINPUT44), .ZN(n424) );
  XNOR2_X1 U411 ( .A(KEYINPUT10), .B(n505), .ZN(n490) );
  XNOR2_X1 U412 ( .A(n725), .B(n439), .ZN(n513) );
  NOR2_X1 U413 ( .A1(n630), .A2(G902), .ZN(n502) );
  OR2_X1 U414 ( .A1(n709), .A2(G902), .ZN(n409) );
  INV_X1 U415 ( .A(G469), .ZN(n444) );
  XNOR2_X1 U416 ( .A(n350), .B(n463), .ZN(n680) );
  XNOR2_X1 U417 ( .A(n462), .B(KEYINPUT25), .ZN(n463) );
  XNOR2_X1 U418 ( .A(n506), .B(n405), .ZN(n488) );
  INV_X1 U419 ( .A(G134), .ZN(n405) );
  XNOR2_X1 U420 ( .A(n389), .B(n388), .ZN(n478) );
  NAND2_X1 U421 ( .A1(G237), .A2(G234), .ZN(n388) );
  XNOR2_X1 U422 ( .A(KEYINPUT14), .B(KEYINPUT94), .ZN(n389) );
  NAND2_X1 U423 ( .A1(n552), .A2(KEYINPUT22), .ZN(n433) );
  INV_X1 U424 ( .A(n549), .ZN(n429) );
  NOR2_X1 U425 ( .A1(n539), .A2(KEYINPUT22), .ZN(n430) );
  NOR2_X1 U426 ( .A1(n718), .A2(G902), .ZN(n489) );
  XNOR2_X1 U427 ( .A(n460), .B(n459), .ZN(n723) );
  XNOR2_X1 U428 ( .A(n451), .B(n450), .ZN(n460) );
  XNOR2_X1 U429 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U430 ( .A(n449), .B(KEYINPUT97), .ZN(n450) );
  AND2_X1 U431 ( .A1(n697), .A2(n611), .ZN(n615) );
  XNOR2_X1 U432 ( .A(n624), .B(KEYINPUT91), .ZN(n724) );
  NAND2_X1 U433 ( .A1(n348), .A2(KEYINPUT47), .ZN(n394) );
  INV_X1 U434 ( .A(KEYINPUT79), .ZN(n385) );
  INV_X1 U435 ( .A(KEYINPUT64), .ZN(n441) );
  INV_X1 U436 ( .A(G237), .ZN(n475) );
  XNOR2_X1 U437 ( .A(G131), .B(G116), .ZN(n465) );
  XOR2_X1 U438 ( .A(KEYINPUT5), .B(G101), .Z(n466) );
  XNOR2_X1 U439 ( .A(KEYINPUT92), .B(KEYINPUT15), .ZN(n445) );
  AND2_X1 U440 ( .A1(n402), .A2(n401), .ZN(n400) );
  NAND2_X1 U441 ( .A1(KEYINPUT17), .A2(G953), .ZN(n401) );
  XNOR2_X1 U442 ( .A(KEYINPUT74), .B(KEYINPUT18), .ZN(n504) );
  INV_X1 U443 ( .A(KEYINPUT2), .ZN(n373) );
  XNOR2_X1 U444 ( .A(n537), .B(n536), .ZN(n669) );
  INV_X1 U445 ( .A(n417), .ZN(n414) );
  NAND2_X1 U446 ( .A1(n516), .A2(G214), .ZN(n665) );
  INV_X1 U447 ( .A(KEYINPUT48), .ZN(n420) );
  XNOR2_X1 U448 ( .A(n464), .B(G119), .ZN(n511) );
  XNOR2_X1 U449 ( .A(G113), .B(KEYINPUT3), .ZN(n464) );
  XNOR2_X1 U450 ( .A(n455), .B(n454), .ZN(n458) );
  XNOR2_X1 U451 ( .A(G119), .B(G128), .ZN(n454) );
  XNOR2_X1 U452 ( .A(G137), .B(G110), .ZN(n452) );
  XNOR2_X1 U453 ( .A(n490), .B(KEYINPUT23), .ZN(n451) );
  XNOR2_X1 U454 ( .A(n419), .B(n737), .ZN(n630) );
  XNOR2_X1 U455 ( .A(n471), .B(n443), .ZN(n709) );
  XOR2_X1 U456 ( .A(n572), .B(KEYINPUT28), .Z(n575) );
  AND2_X1 U457 ( .A1(n542), .A2(n580), .ZN(n572) );
  XNOR2_X1 U458 ( .A(n535), .B(n422), .ZN(n562) );
  INV_X1 U459 ( .A(KEYINPUT102), .ZN(n422) );
  XNOR2_X1 U460 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U461 ( .A(n512), .B(n511), .ZN(n727) );
  XNOR2_X1 U462 ( .A(n510), .B(KEYINPUT16), .ZN(n512) );
  XNOR2_X1 U463 ( .A(n488), .B(n487), .ZN(n386) );
  XNOR2_X1 U464 ( .A(n486), .B(n485), .ZN(n387) );
  XNOR2_X1 U465 ( .A(n630), .B(KEYINPUT59), .ZN(n631) );
  NAND2_X1 U466 ( .A1(n351), .A2(n428), .ZN(n370) );
  AND2_X1 U467 ( .A1(n352), .A2(n540), .ZN(n371) );
  XNOR2_X1 U468 ( .A(n559), .B(n378), .ZN(n661) );
  INV_X1 U469 ( .A(KEYINPUT31), .ZN(n378) );
  NOR2_X1 U470 ( .A1(n427), .A2(n426), .ZN(n565) );
  XNOR2_X1 U471 ( .A(n722), .B(n723), .ZN(n379) );
  NOR2_X1 U472 ( .A1(n705), .A2(G953), .ZN(n706) );
  OR2_X1 U473 ( .A1(n396), .A2(n395), .ZN(n348) );
  XOR2_X1 U474 ( .A(n518), .B(n517), .Z(n349) );
  OR2_X1 U475 ( .A1(G902), .A2(n723), .ZN(n350) );
  BUF_X1 U476 ( .A(n552), .Z(n557) );
  AND2_X1 U477 ( .A1(n433), .A2(n371), .ZN(n351) );
  AND2_X1 U478 ( .A1(n432), .A2(n429), .ZN(n352) );
  OR2_X1 U479 ( .A1(n533), .A2(n532), .ZN(n353) );
  AND2_X1 U480 ( .A1(n549), .A2(n581), .ZN(n354) );
  AND2_X1 U481 ( .A1(n416), .A2(n554), .ZN(n355) );
  AND2_X1 U482 ( .A1(n578), .A2(n394), .ZN(n356) );
  XOR2_X1 U483 ( .A(n444), .B(KEYINPUT68), .Z(n357) );
  AND2_X1 U484 ( .A1(G214), .A2(n498), .ZN(n358) );
  AND2_X1 U485 ( .A1(n604), .A2(n576), .ZN(n359) );
  AND2_X1 U486 ( .A1(n549), .A2(n655), .ZN(n360) );
  AND2_X1 U487 ( .A1(n433), .A2(n432), .ZN(n361) );
  NAND2_X1 U488 ( .A1(n659), .A2(n662), .ZN(n666) );
  INV_X1 U489 ( .A(n666), .ZN(n396) );
  NAND2_X1 U490 ( .A1(n366), .A2(n362), .ZN(n571) );
  NOR2_X1 U491 ( .A1(n363), .A2(n644), .ZN(n362) );
  XNOR2_X1 U492 ( .A(n367), .B(n424), .ZN(n366) );
  NAND2_X1 U493 ( .A1(n369), .A2(n368), .ZN(n367) );
  INV_X1 U494 ( .A(n754), .ZN(n368) );
  XNOR2_X1 U495 ( .A(n548), .B(n425), .ZN(n369) );
  NAND2_X1 U496 ( .A1(n431), .A2(n430), .ZN(n428) );
  NOR2_X2 U497 ( .A1(n730), .A2(n739), .ZN(n697) );
  NAND2_X1 U498 ( .A1(n374), .A2(n372), .ZN(n375) );
  NOR2_X2 U499 ( .A1(n616), .A2(n700), .ZN(n717) );
  XNOR2_X1 U500 ( .A(n376), .B(n508), .ZN(n515) );
  XNOR2_X1 U501 ( .A(n509), .B(n507), .ZN(n376) );
  NAND2_X1 U502 ( .A1(n400), .A2(n399), .ZN(n404) );
  INV_X2 U503 ( .A(G116), .ZN(n377) );
  XNOR2_X2 U504 ( .A(G110), .B(G107), .ZN(n437) );
  INV_X1 U505 ( .A(n651), .ZN(n546) );
  XNOR2_X2 U506 ( .A(n534), .B(KEYINPUT0), .ZN(n552) );
  XNOR2_X2 U507 ( .A(n377), .B(G122), .ZN(n510) );
  XNOR2_X1 U508 ( .A(n381), .B(n420), .ZN(n380) );
  NOR2_X1 U509 ( .A1(n379), .A2(n724), .ZN(G66) );
  NAND2_X1 U510 ( .A1(n380), .A2(n610), .ZN(n739) );
  NAND2_X1 U511 ( .A1(n383), .A2(n382), .ZN(n381) );
  XNOR2_X1 U512 ( .A(n607), .B(KEYINPUT46), .ZN(n382) );
  AND2_X1 U513 ( .A1(n592), .A2(n435), .ZN(n383) );
  NAND2_X1 U514 ( .A1(n356), .A2(n392), .ZN(n579) );
  NAND2_X1 U515 ( .A1(n393), .A2(KEYINPUT47), .ZN(n392) );
  INV_X1 U516 ( .A(n604), .ZN(n393) );
  INV_X1 U517 ( .A(n576), .ZN(n395) );
  NAND2_X1 U518 ( .A1(n576), .A2(n353), .ZN(n534) );
  XNOR2_X2 U519 ( .A(n581), .B(n423), .ZN(n576) );
  XNOR2_X2 U520 ( .A(n397), .B(KEYINPUT87), .ZN(n581) );
  NAND2_X2 U521 ( .A1(n530), .A2(n665), .ZN(n397) );
  INV_X1 U522 ( .A(n547), .ZN(n629) );
  NAND2_X1 U523 ( .A1(n398), .A2(G224), .ZN(n399) );
  INV_X1 U524 ( .A(G224), .ZN(n403) );
  NAND2_X1 U525 ( .A1(n403), .A2(KEYINPUT17), .ZN(n402) );
  XNOR2_X1 U526 ( .A(n404), .B(n504), .ZN(n508) );
  NOR2_X2 U527 ( .A1(n545), .A2(n544), .ZN(n651) );
  XNOR2_X2 U528 ( .A(n573), .B(KEYINPUT1), .ZN(n676) );
  XNOR2_X2 U529 ( .A(n409), .B(n357), .ZN(n573) );
  NAND2_X1 U530 ( .A1(n410), .A2(n355), .ZN(n556) );
  NAND2_X1 U531 ( .A1(n413), .A2(n411), .ZN(n410) );
  NAND2_X1 U532 ( .A1(n701), .A2(n412), .ZN(n411) );
  INV_X1 U533 ( .A(KEYINPUT34), .ZN(n412) );
  NAND2_X1 U534 ( .A1(n415), .A2(n414), .ZN(n413) );
  INV_X1 U535 ( .A(n701), .ZN(n415) );
  NAND2_X1 U536 ( .A1(n557), .A2(KEYINPUT34), .ZN(n416) );
  NOR2_X2 U537 ( .A1(n557), .A2(KEYINPUT34), .ZN(n417) );
  XNOR2_X1 U538 ( .A(n418), .B(n358), .ZN(n419) );
  XNOR2_X1 U539 ( .A(n497), .B(n496), .ZN(n418) );
  XNOR2_X2 U540 ( .A(n421), .B(KEYINPUT103), .ZN(n659) );
  NOR2_X1 U541 ( .A1(n562), .A2(n563), .ZN(n421) );
  NAND2_X1 U542 ( .A1(n655), .A2(n354), .ZN(n582) );
  NAND2_X1 U543 ( .A1(n525), .A2(n360), .ZN(n526) );
  INV_X1 U544 ( .A(KEYINPUT19), .ZN(n423) );
  INV_X1 U545 ( .A(KEYINPUT86), .ZN(n425) );
  NAND2_X1 U546 ( .A1(n352), .A2(n433), .ZN(n426) );
  INV_X1 U547 ( .A(n428), .ZN(n427) );
  NAND2_X1 U548 ( .A1(n361), .A2(n428), .ZN(n545) );
  INV_X1 U549 ( .A(n552), .ZN(n431) );
  NAND2_X1 U550 ( .A1(n539), .A2(KEYINPUT22), .ZN(n432) );
  NOR2_X1 U551 ( .A1(n652), .A2(n590), .ZN(n434) );
  XOR2_X1 U552 ( .A(n579), .B(KEYINPUT78), .Z(n435) );
  INV_X1 U553 ( .A(KEYINPUT83), .ZN(n587) );
  XNOR2_X1 U554 ( .A(n752), .B(n587), .ZN(n591) );
  NOR2_X1 U555 ( .A1(n591), .A2(n434), .ZN(n592) );
  INV_X1 U556 ( .A(KEYINPUT70), .ZN(n472) );
  XNOR2_X1 U557 ( .A(n472), .B(G472), .ZN(n473) );
  INV_X1 U558 ( .A(KEYINPUT96), .ZN(n449) );
  INV_X1 U559 ( .A(KEYINPUT45), .ZN(n570) );
  XNOR2_X1 U560 ( .A(KEYINPUT39), .B(KEYINPUT84), .ZN(n599) );
  XOR2_X1 U561 ( .A(G131), .B(G140), .Z(n491) );
  NAND2_X1 U562 ( .A1(G227), .A2(n741), .ZN(n436) );
  XNOR2_X1 U563 ( .A(n491), .B(n436), .ZN(n440) );
  INV_X1 U564 ( .A(KEYINPUT69), .ZN(n439) );
  XNOR2_X1 U565 ( .A(n440), .B(n513), .ZN(n443) );
  XNOR2_X1 U566 ( .A(n445), .B(G902), .ZN(n612) );
  NAND2_X1 U567 ( .A1(n612), .A2(G234), .ZN(n446) );
  XNOR2_X1 U568 ( .A(KEYINPUT20), .B(n446), .ZN(n461) );
  AND2_X1 U569 ( .A1(n461), .A2(G221), .ZN(n448) );
  INV_X1 U570 ( .A(KEYINPUT21), .ZN(n447) );
  XNOR2_X1 U571 ( .A(n448), .B(n447), .ZN(n679) );
  XNOR2_X2 U572 ( .A(G146), .B(G125), .ZN(n505) );
  XOR2_X1 U573 ( .A(KEYINPUT24), .B(G140), .Z(n453) );
  XNOR2_X1 U574 ( .A(n453), .B(n452), .ZN(n455) );
  NAND2_X1 U575 ( .A1(G234), .A2(n741), .ZN(n456) );
  XOR2_X1 U576 ( .A(KEYINPUT8), .B(n456), .Z(n484) );
  AND2_X1 U577 ( .A1(G221), .A2(n484), .ZN(n457) );
  NAND2_X1 U578 ( .A1(G217), .A2(n461), .ZN(n462) );
  NOR2_X1 U579 ( .A1(n679), .A2(n680), .ZN(n675) );
  NAND2_X1 U580 ( .A1(n573), .A2(n675), .ZN(n560) );
  XNOR2_X1 U581 ( .A(n560), .B(KEYINPUT107), .ZN(n598) );
  XNOR2_X1 U582 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U583 ( .A(n511), .B(n467), .Z(n469) );
  NOR2_X1 U584 ( .A1(G953), .A2(G237), .ZN(n498) );
  NAND2_X1 U585 ( .A1(n498), .A2(G210), .ZN(n468) );
  XNOR2_X1 U586 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U587 ( .A(n471), .B(n470), .ZN(n620) );
  XNOR2_X2 U588 ( .A(n474), .B(n473), .ZN(n541) );
  INV_X1 U589 ( .A(G902), .ZN(n476) );
  NAND2_X1 U590 ( .A1(n476), .A2(n475), .ZN(n516) );
  NAND2_X1 U591 ( .A1(n541), .A2(n665), .ZN(n477) );
  XNOR2_X1 U592 ( .A(KEYINPUT30), .B(n477), .ZN(n483) );
  NAND2_X1 U593 ( .A1(G952), .A2(n478), .ZN(n695) );
  NOR2_X1 U594 ( .A1(n695), .A2(G953), .ZN(n532) );
  NAND2_X1 U595 ( .A1(n478), .A2(G902), .ZN(n479) );
  XNOR2_X1 U596 ( .A(n479), .B(KEYINPUT95), .ZN(n531) );
  NAND2_X1 U597 ( .A1(G953), .A2(n531), .ZN(n480) );
  NOR2_X1 U598 ( .A1(G900), .A2(n480), .ZN(n481) );
  NOR2_X1 U599 ( .A1(n532), .A2(n481), .ZN(n482) );
  XOR2_X1 U600 ( .A(KEYINPUT75), .B(n482), .Z(n523) );
  NAND2_X1 U601 ( .A1(n598), .A2(n596), .ZN(n503) );
  XNOR2_X1 U602 ( .A(G107), .B(KEYINPUT9), .ZN(n487) );
  XOR2_X1 U603 ( .A(n510), .B(KEYINPUT7), .Z(n486) );
  NAND2_X1 U604 ( .A1(G217), .A2(n484), .ZN(n485) );
  XOR2_X1 U605 ( .A(G478), .B(n489), .Z(n563) );
  XNOR2_X1 U606 ( .A(n491), .B(n490), .ZN(n737) );
  XOR2_X1 U607 ( .A(G104), .B(G122), .Z(n493) );
  XNOR2_X1 U608 ( .A(G113), .B(G143), .ZN(n492) );
  XNOR2_X1 U609 ( .A(n493), .B(n492), .ZN(n497) );
  XOR2_X1 U610 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n495) );
  XNOR2_X1 U611 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n494) );
  XNOR2_X1 U612 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U613 ( .A(KEYINPUT100), .B(KEYINPUT13), .Z(n500) );
  XNOR2_X1 U614 ( .A(KEYINPUT101), .B(G475), .ZN(n499) );
  XNOR2_X1 U615 ( .A(n500), .B(n499), .ZN(n501) );
  NAND2_X1 U616 ( .A1(n563), .A2(n535), .ZN(n553) );
  NOR2_X1 U617 ( .A1(n503), .A2(n553), .ZN(n520) );
  XNOR2_X1 U618 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U619 ( .A(n727), .B(n513), .ZN(n514) );
  XNOR2_X1 U620 ( .A(n514), .B(n515), .ZN(n637) );
  NAND2_X1 U621 ( .A1(n637), .A2(n612), .ZN(n519) );
  NAND2_X1 U622 ( .A1(n516), .A2(G210), .ZN(n518) );
  INV_X1 U623 ( .A(KEYINPUT93), .ZN(n517) );
  XNOR2_X2 U624 ( .A(n519), .B(n349), .ZN(n530) );
  BUF_X1 U625 ( .A(n530), .Z(n528) );
  NAND2_X1 U626 ( .A1(n520), .A2(n528), .ZN(n577) );
  XOR2_X1 U627 ( .A(G143), .B(KEYINPUT113), .Z(n521) );
  XNOR2_X1 U628 ( .A(n577), .B(n521), .ZN(G45) );
  INV_X1 U629 ( .A(KEYINPUT6), .ZN(n522) );
  INV_X1 U630 ( .A(n679), .ZN(n538) );
  NAND2_X1 U631 ( .A1(n580), .A2(n665), .ZN(n524) );
  NOR2_X1 U632 ( .A1(n524), .A2(n676), .ZN(n525) );
  XNOR2_X1 U633 ( .A(KEYINPUT106), .B(n526), .ZN(n527) );
  XNOR2_X1 U634 ( .A(n527), .B(KEYINPUT43), .ZN(n529) );
  INV_X1 U635 ( .A(n528), .ZN(n594) );
  AND2_X1 U636 ( .A1(n529), .A2(n594), .ZN(n609) );
  XOR2_X1 U637 ( .A(n609), .B(G140), .Z(G42) );
  NOR2_X1 U638 ( .A1(G898), .A2(n741), .ZN(n728) );
  AND2_X1 U639 ( .A1(n531), .A2(n728), .ZN(n533) );
  NOR2_X1 U640 ( .A1(n563), .A2(n535), .ZN(n537) );
  INV_X1 U641 ( .A(KEYINPUT105), .ZN(n536) );
  NAND2_X1 U642 ( .A1(n669), .A2(n538), .ZN(n539) );
  INV_X1 U643 ( .A(n676), .ZN(n567) );
  INV_X1 U644 ( .A(n680), .ZN(n566) );
  NOR2_X1 U645 ( .A1(n567), .A2(n566), .ZN(n540) );
  NOR2_X1 U646 ( .A1(n542), .A2(n566), .ZN(n543) );
  NAND2_X1 U647 ( .A1(n567), .A2(n543), .ZN(n544) );
  NAND2_X1 U648 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U649 ( .A(KEYINPUT88), .B(KEYINPUT33), .Z(n551) );
  AND2_X1 U650 ( .A1(n676), .A2(n675), .ZN(n558) );
  NAND2_X1 U651 ( .A1(n558), .A2(n549), .ZN(n550) );
  INV_X1 U652 ( .A(n553), .ZN(n554) );
  XNOR2_X1 U653 ( .A(KEYINPUT82), .B(KEYINPUT35), .ZN(n555) );
  XNOR2_X1 U654 ( .A(n556), .B(n555), .ZN(n754) );
  AND2_X1 U655 ( .A1(n542), .A2(n558), .ZN(n687) );
  NAND2_X1 U656 ( .A1(n431), .A2(n687), .ZN(n559) );
  NOR2_X1 U657 ( .A1(n560), .A2(n542), .ZN(n561) );
  NAND2_X1 U658 ( .A1(n431), .A2(n561), .ZN(n647) );
  NAND2_X1 U659 ( .A1(n563), .A2(n562), .ZN(n662) );
  XNOR2_X1 U660 ( .A(n565), .B(KEYINPUT85), .ZN(n569) );
  NAND2_X1 U661 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U662 ( .A1(n569), .A2(n568), .ZN(n644) );
  XNOR2_X2 U663 ( .A(n571), .B(n570), .ZN(n730) );
  INV_X1 U664 ( .A(n573), .ZN(n574) );
  XNOR2_X1 U665 ( .A(n577), .B(KEYINPUT80), .ZN(n578) );
  INV_X1 U666 ( .A(n580), .ZN(n583) );
  NAND2_X1 U667 ( .A1(n585), .A2(n676), .ZN(n586) );
  XNOR2_X2 U668 ( .A(n586), .B(KEYINPUT109), .ZN(n752) );
  INV_X1 U669 ( .A(n359), .ZN(n652) );
  XNOR2_X1 U670 ( .A(n589), .B(KEYINPUT71), .ZN(n590) );
  XOR2_X1 U671 ( .A(KEYINPUT72), .B(KEYINPUT38), .Z(n593) );
  XNOR2_X1 U672 ( .A(n594), .B(n593), .ZN(n667) );
  INV_X1 U673 ( .A(n667), .ZN(n595) );
  AND2_X1 U674 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U675 ( .A(n600), .B(n599), .ZN(n608) );
  NOR2_X1 U676 ( .A1(n608), .A2(n659), .ZN(n601) );
  INV_X1 U677 ( .A(n669), .ZN(n602) );
  NOR2_X1 U678 ( .A1(n667), .A2(n602), .ZN(n673) );
  NAND2_X1 U679 ( .A1(n665), .A2(n673), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n604), .A2(n702), .ZN(n606) );
  XOR2_X1 U681 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n605) );
  XNOR2_X1 U682 ( .A(n606), .B(n605), .ZN(n751) );
  NOR2_X1 U683 ( .A1(n608), .A2(n662), .ZN(n664) );
  NOR2_X1 U684 ( .A1(n664), .A2(n609), .ZN(n610) );
  INV_X1 U685 ( .A(n612), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n612), .B(KEYINPUT81), .ZN(n613) );
  AND2_X1 U687 ( .A1(n613), .A2(KEYINPUT2), .ZN(n614) );
  NOR2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n717), .A2(G472), .ZN(n622) );
  XOR2_X1 U690 ( .A(KEYINPUT62), .B(KEYINPUT110), .Z(n618) );
  XNOR2_X1 U691 ( .A(KEYINPUT111), .B(KEYINPUT89), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n622), .B(n621), .ZN(n625) );
  INV_X1 U694 ( .A(G952), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n623), .A2(G953), .ZN(n624) );
  INV_X1 U696 ( .A(n724), .ZN(n640) );
  NAND2_X1 U697 ( .A1(n625), .A2(n640), .ZN(n627) );
  XNOR2_X1 U698 ( .A(KEYINPUT90), .B(KEYINPUT63), .ZN(n626) );
  XNOR2_X1 U699 ( .A(n627), .B(n626), .ZN(G57) );
  XNOR2_X1 U700 ( .A(G119), .B(KEYINPUT127), .ZN(n628) );
  XNOR2_X1 U701 ( .A(n629), .B(n628), .ZN(G21) );
  NAND2_X1 U702 ( .A1(n717), .A2(G475), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n632), .B(n631), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n633), .A2(n640), .ZN(n635) );
  XNOR2_X1 U705 ( .A(KEYINPUT65), .B(KEYINPUT60), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(G60) );
  NAND2_X1 U707 ( .A1(n717), .A2(G210), .ZN(n639) );
  XOR2_X1 U708 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n636) );
  XNOR2_X1 U709 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n639), .B(n638), .ZN(n641) );
  NAND2_X1 U711 ( .A1(n641), .A2(n640), .ZN(n643) );
  INV_X1 U712 ( .A(KEYINPUT56), .ZN(n642) );
  XNOR2_X1 U713 ( .A(n643), .B(n642), .ZN(G51) );
  XOR2_X1 U714 ( .A(G101), .B(n644), .Z(n645) );
  XNOR2_X1 U715 ( .A(KEYINPUT112), .B(n645), .ZN(G3) );
  NOR2_X1 U716 ( .A1(n659), .A2(n647), .ZN(n646) );
  XOR2_X1 U717 ( .A(G104), .B(n646), .Z(G6) );
  NOR2_X1 U718 ( .A1(n662), .A2(n647), .ZN(n649) );
  XNOR2_X1 U719 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U721 ( .A(G107), .B(n650), .ZN(G9) );
  XOR2_X1 U722 ( .A(G110), .B(n651), .Z(G12) );
  NOR2_X1 U723 ( .A1(n652), .A2(n662), .ZN(n654) );
  XNOR2_X1 U724 ( .A(G128), .B(KEYINPUT29), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n654), .B(n653), .ZN(G30) );
  XOR2_X1 U726 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n657) );
  NAND2_X1 U727 ( .A1(n359), .A2(n655), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U729 ( .A(G146), .B(n658), .ZN(G48) );
  NOR2_X1 U730 ( .A1(n659), .A2(n661), .ZN(n660) );
  XOR2_X1 U731 ( .A(G113), .B(n660), .Z(G15) );
  NOR2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U733 ( .A(G116), .B(n663), .Z(G18) );
  XOR2_X1 U734 ( .A(G134), .B(n664), .Z(G36) );
  INV_X1 U735 ( .A(n665), .ZN(n671) );
  NOR2_X1 U736 ( .A1(n667), .A2(n396), .ZN(n668) );
  NOR2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n701), .A2(n674), .ZN(n692) );
  XNOR2_X1 U741 ( .A(KEYINPUT117), .B(KEYINPUT50), .ZN(n678) );
  NOR2_X1 U742 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U743 ( .A(n678), .B(n677), .ZN(n684) );
  XOR2_X1 U744 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n682) );
  NAND2_X1 U745 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U746 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U748 ( .A1(n542), .A2(n685), .ZN(n686) );
  NOR2_X1 U749 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U750 ( .A(KEYINPUT51), .B(n688), .ZN(n689) );
  NAND2_X1 U751 ( .A1(n689), .A2(n702), .ZN(n690) );
  XOR2_X1 U752 ( .A(KEYINPUT118), .B(n690), .Z(n691) );
  NOR2_X1 U753 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U754 ( .A(n693), .B(KEYINPUT52), .ZN(n694) );
  OR2_X1 U755 ( .A1(n695), .A2(n694), .ZN(n707) );
  XOR2_X1 U756 ( .A(KEYINPUT2), .B(KEYINPUT77), .Z(n696) );
  NOR2_X1 U757 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U758 ( .A(n698), .B(KEYINPUT76), .ZN(n699) );
  OR2_X1 U759 ( .A1(n700), .A2(n699), .ZN(n704) );
  NAND2_X1 U760 ( .A1(n702), .A2(n415), .ZN(n703) );
  NAND2_X1 U761 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U762 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U763 ( .A(KEYINPUT53), .B(n708), .Z(G75) );
  XOR2_X1 U764 ( .A(KEYINPUT119), .B(KEYINPUT121), .Z(n711) );
  XNOR2_X1 U765 ( .A(n709), .B(KEYINPUT120), .ZN(n710) );
  XNOR2_X1 U766 ( .A(n711), .B(n710), .ZN(n713) );
  XOR2_X1 U767 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n712) );
  XNOR2_X1 U768 ( .A(n713), .B(n712), .ZN(n715) );
  NAND2_X1 U769 ( .A1(n717), .A2(G469), .ZN(n714) );
  XOR2_X1 U770 ( .A(n715), .B(n714), .Z(n716) );
  NOR2_X1 U771 ( .A1(n724), .A2(n716), .ZN(G54) );
  NAND2_X1 U772 ( .A1(n717), .A2(G478), .ZN(n720) );
  XNOR2_X1 U773 ( .A(n718), .B(KEYINPUT122), .ZN(n719) );
  XNOR2_X1 U774 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U775 ( .A1(n724), .A2(n721), .ZN(G63) );
  NAND2_X1 U776 ( .A1(n717), .A2(G217), .ZN(n722) );
  XNOR2_X1 U777 ( .A(n725), .B(KEYINPUT123), .ZN(n726) );
  XNOR2_X1 U778 ( .A(n727), .B(n726), .ZN(n729) );
  NOR2_X1 U779 ( .A1(n729), .A2(n728), .ZN(n736) );
  OR2_X1 U780 ( .A1(n730), .A2(G953), .ZN(n734) );
  NAND2_X1 U781 ( .A1(G953), .A2(G224), .ZN(n731) );
  XNOR2_X1 U782 ( .A(n731), .B(KEYINPUT61), .ZN(n732) );
  NAND2_X1 U783 ( .A1(n732), .A2(G898), .ZN(n733) );
  NAND2_X1 U784 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U785 ( .A(n736), .B(n735), .ZN(G69) );
  XOR2_X1 U786 ( .A(n738), .B(n737), .Z(n744) );
  INV_X1 U787 ( .A(n744), .ZN(n740) );
  XNOR2_X1 U788 ( .A(n740), .B(n739), .ZN(n742) );
  NAND2_X1 U789 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U790 ( .A(KEYINPUT124), .B(n743), .ZN(n750) );
  XNOR2_X1 U791 ( .A(n744), .B(G227), .ZN(n745) );
  XNOR2_X1 U792 ( .A(n745), .B(KEYINPUT125), .ZN(n746) );
  NAND2_X1 U793 ( .A1(n746), .A2(G900), .ZN(n747) );
  NAND2_X1 U794 ( .A1(G953), .A2(n747), .ZN(n748) );
  XNOR2_X1 U795 ( .A(KEYINPUT126), .B(n748), .ZN(n749) );
  NAND2_X1 U796 ( .A1(n750), .A2(n749), .ZN(G72) );
  XOR2_X1 U797 ( .A(G137), .B(n751), .Z(G39) );
  XNOR2_X1 U798 ( .A(n752), .B(G125), .ZN(n753) );
  XNOR2_X1 U799 ( .A(n753), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U800 ( .A(G122), .B(n754), .Z(G24) );
  XOR2_X1 U801 ( .A(n755), .B(G131), .Z(G33) );
endmodule

