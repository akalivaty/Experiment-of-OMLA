//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(G8gat), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G71gat), .A2(G78gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G71gat), .A2(G78gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n209), .A2(KEYINPUT9), .ZN(new_n212));
  XNOR2_X1  g011(.A(G57gat), .B(G64gat), .ZN(new_n213));
  OR3_X1    g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n207), .B1(KEYINPUT21), .B2(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n216), .A2(KEYINPUT21), .ZN(new_n220));
  NAND2_X1  g019(.A1(G231gat), .A2(G233gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n219), .B(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G183gat), .B(G211gat), .Z(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G127gat), .B(G155gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n223), .B(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(KEYINPUT96), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT95), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT96), .B1(new_n233), .B2(new_n231), .ZN(new_n234));
  MUX2_X1   g033(.A(new_n230), .B(new_n232), .S(new_n234), .Z(new_n235));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236));
  NAND2_X1  g035(.A1(G99gat), .A2(G106gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(KEYINPUT97), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(KEYINPUT97), .B2(new_n237), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT98), .B(G85gat), .ZN(new_n240));
  INV_X1    g039(.A(G92gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT99), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n239), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n243), .B1(new_n239), .B2(new_n242), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n235), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G99gat), .B(G106gat), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n247), .B(new_n235), .C1(new_n244), .C2(new_n245), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(KEYINPUT100), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT100), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n246), .A2(new_n252), .A3(new_n248), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT101), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT101), .B1(new_n251), .B2(new_n253), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT14), .ZN(new_n259));
  INV_X1    g058(.A(G29gat), .ZN(new_n260));
  INV_X1    g059(.A(G36gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n262), .A2(new_n263), .B1(G29gat), .B2(G36gat), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n264), .A2(KEYINPUT15), .ZN(new_n265));
  XNOR2_X1  g064(.A(G43gat), .B(G50gat), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n264), .A2(KEYINPUT15), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n258), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n270), .A2(KEYINPUT17), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(KEYINPUT17), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n273), .B(new_n274), .C1(new_n256), .C2(new_n257), .ZN(new_n275));
  AND2_X1   g074(.A1(G232gat), .A2(G233gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT41), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n272), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(G134gat), .B(G162gat), .Z(new_n279));
  AND2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n278), .A2(new_n279), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n276), .A2(KEYINPUT41), .ZN(new_n283));
  XNOR2_X1  g082(.A(G190gat), .B(G218gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n285), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(new_n280), .B2(new_n281), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT92), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT34), .ZN(new_n292));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT24), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G169gat), .ZN(new_n305));
  INV_X1    g104(.A(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g106(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(new_n295), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT25), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n298), .A2(new_n304), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  OR2_X1    g111(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n314));
  AOI21_X1  g113(.A(G190gat), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT28), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT67), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT67), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT28), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G190gat), .ZN(new_n322));
  AND2_X1   g121(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n321), .A2(new_n327), .A3(new_n299), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n329), .A2(new_n330), .A3(new_n293), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n330), .B1(new_n329), .B2(new_n293), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n307), .A2(KEYINPUT26), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n312), .B1(new_n328), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n299), .A2(KEYINPUT65), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT65), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(G183gat), .A3(G190gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n339), .A3(new_n300), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT66), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n337), .A2(new_n339), .A3(KEYINPUT66), .A4(new_n300), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n302), .A2(new_n303), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n298), .A2(new_n309), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT25), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n336), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n310), .B1(new_n345), .B2(new_n347), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n321), .A2(new_n327), .A3(new_n299), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n311), .B1(new_n353), .B2(new_n334), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT73), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n356));
  INV_X1    g155(.A(G113gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G120gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT71), .B(G120gat), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n359), .B1(new_n360), .B2(G113gat), .ZN(new_n361));
  INV_X1    g160(.A(G127gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G134gat), .ZN(new_n363));
  INV_X1    g162(.A(G134gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G127gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT1), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n356), .B1(new_n361), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT69), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n362), .A2(KEYINPUT69), .A3(G134gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n365), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G120gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G113gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT70), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n366), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n375), .B1(new_n358), .B2(new_n374), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n372), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n367), .ZN(new_n380));
  OR2_X1    g179(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n357), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n380), .B(KEYINPUT72), .C1(new_n383), .C2(new_n359), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n379), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n351), .A2(new_n355), .A3(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n336), .A2(new_n349), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n368), .A2(new_n379), .A3(new_n384), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(KEYINPUT73), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n292), .B1(new_n391), .B2(KEYINPUT32), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT74), .B(KEYINPUT33), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G15gat), .B(G43gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(G71gat), .B(G99gat), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n396), .B(new_n397), .Z(new_n398));
  NAND2_X1  g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n391), .A2(KEYINPUT32), .A3(new_n292), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n393), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n398), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n402), .B1(new_n391), .B2(new_n394), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n391), .A2(KEYINPUT32), .A3(new_n292), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(new_n404), .B2(new_n392), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n387), .B1(new_n386), .B2(new_n390), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(KEYINPUT75), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n401), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n401), .B2(new_n405), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n291), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n407), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n399), .B1(new_n393), .B2(new_n400), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n404), .A2(new_n392), .A3(new_n403), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n401), .A2(new_n405), .A3(new_n407), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(KEYINPUT92), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G141gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G148gat), .ZN(new_n418));
  INV_X1    g217(.A(G148gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G141gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G155gat), .B(G162gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(G155gat), .A2(G162gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT2), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n422), .B1(new_n424), .B2(new_n421), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT78), .B(G211gat), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT22), .B1(new_n428), .B2(G218gat), .ZN(new_n429));
  XOR2_X1   g228(.A(G197gat), .B(G204gat), .Z(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G211gat), .B(G218gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT3), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n427), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n433), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n424), .ZN(new_n441));
  OR2_X1    g240(.A1(G155gat), .A2(G162gat), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n442), .A2(new_n423), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n436), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n434), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n437), .B2(new_n438), .ZN(new_n449));
  INV_X1    g248(.A(G228gat), .ZN(new_n450));
  INV_X1    g249(.A(G233gat), .ZN(new_n451));
  OAI22_X1  g250(.A1(new_n439), .A2(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n437), .A2(KEYINPUT84), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n450), .A2(new_n451), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n437), .A2(KEYINPUT84), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n453), .A2(new_n454), .A3(new_n448), .A4(new_n455), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(G78gat), .B(G106gat), .Z(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(G22gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT31), .B(G50gat), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n459), .B(new_n460), .Z(new_n461));
  OR2_X1    g260(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n452), .A2(new_n456), .A3(new_n461), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n410), .A2(new_n416), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT91), .ZN(new_n466));
  XOR2_X1   g265(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n467));
  OAI21_X1  g266(.A(KEYINPUT3), .B1(new_n425), .B2(new_n426), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n446), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n389), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n427), .A2(new_n368), .A3(new_n379), .A4(new_n384), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(G225gat), .A2(G233gat), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT4), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n473), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n427), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n385), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n479), .A2(KEYINPUT81), .A3(new_n471), .ZN(new_n480));
  INV_X1    g279(.A(new_n473), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT81), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n385), .A2(new_n482), .A3(new_n478), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n477), .A2(KEYINPUT5), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n473), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(KEYINPUT4), .B(new_n471), .C1(new_n389), .C2(new_n469), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n471), .A2(new_n467), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G1gat), .B(G29gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(G85gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT0), .B(G57gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n492), .A2(KEYINPUT6), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT82), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT82), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n492), .A2(new_n499), .A3(KEYINPUT6), .A4(new_n496), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT88), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n486), .B1(new_n472), .B2(new_n476), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n490), .B1(new_n503), .B2(new_n484), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n496), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI211_X1 g305(.A(KEYINPUT87), .B(new_n490), .C1(new_n503), .C2(new_n484), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n492), .A2(KEYINPUT87), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n504), .A2(new_n505), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT88), .A4(new_n496), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n492), .A2(new_n496), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n501), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT79), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n336), .A2(new_n349), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT79), .B1(new_n352), .B2(new_n354), .ZN(new_n519));
  NAND2_X1  g318(.A1(G226gat), .A2(G233gat), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(KEYINPUT29), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n518), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n352), .A2(new_n354), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n521), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n440), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n518), .A2(new_n519), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n521), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n388), .A2(new_n522), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n440), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G8gat), .B(G36gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(G64gat), .B(G92gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n527), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n520), .B1(new_n518), .B2(new_n519), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n524), .A2(KEYINPUT29), .A3(new_n521), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n537), .A2(new_n538), .A3(new_n433), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n534), .B1(new_n539), .B2(new_n526), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n540), .A3(KEYINPUT30), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n539), .A2(new_n526), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(new_n543), .A3(new_n535), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n466), .B1(new_n516), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT35), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n513), .A2(new_n514), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n549), .B1(new_n508), .B2(new_n511), .ZN(new_n550));
  OAI211_X1 g349(.A(KEYINPUT91), .B(new_n545), .C1(new_n550), .C2(new_n501), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n465), .A2(new_n547), .A3(new_n548), .A4(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n408), .A2(new_n409), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n464), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n492), .A2(new_n496), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n515), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n501), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n545), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT35), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n552), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n512), .A2(new_n515), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT90), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT37), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n527), .B2(new_n531), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n566), .B2(new_n535), .ZN(new_n567));
  OAI211_X1 g366(.A(KEYINPUT90), .B(new_n534), .C1(new_n542), .C2(new_n565), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n542), .A2(new_n565), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT38), .ZN(new_n571));
  AOI211_X1 g370(.A(KEYINPUT38), .B(new_n535), .C1(new_n542), .C2(new_n565), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n529), .A2(new_n433), .A3(new_n530), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n523), .A2(new_n525), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n573), .B(KEYINPUT37), .C1(new_n433), .C2(new_n574), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n572), .A2(new_n575), .B1(new_n542), .B2(new_n535), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n563), .A2(new_n571), .A3(new_n558), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n480), .A2(new_n483), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n473), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n579), .A2(KEYINPUT86), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT39), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n581), .B1(new_n579), .B2(KEYINPUT86), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT85), .A4(new_n481), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n488), .A2(new_n489), .A3(new_n481), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT85), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n580), .A2(new_n582), .A3(new_n583), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n583), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n496), .B1(new_n588), .B2(new_n581), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(KEYINPUT40), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT89), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT40), .B1(new_n587), .B2(new_n589), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n545), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n590), .A2(new_n591), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n592), .A2(new_n594), .A3(new_n512), .A4(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n577), .A2(new_n464), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n464), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n560), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT77), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n601));
  NAND2_X1  g400(.A1(new_n553), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT36), .B1(new_n408), .B2(new_n409), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT77), .B1(new_n553), .B2(new_n601), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n597), .B(new_n599), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  AOI211_X1 g405(.A(new_n229), .B(new_n290), .C1(new_n562), .C2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n273), .A2(new_n206), .A3(new_n274), .ZN(new_n608));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n207), .A2(new_n271), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT18), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n206), .A2(new_n270), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n609), .B(KEYINPUT13), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G113gat), .B(G141gat), .ZN(new_n620));
  INV_X1    g419(.A(G197gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT11), .B(G169gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  XOR2_X1   g423(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n613), .A2(new_n614), .A3(new_n618), .A4(new_n625), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G204gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT104), .B(G176gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n249), .A2(new_n634), .A3(new_n250), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n246), .A2(KEYINPUT102), .A3(new_n248), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(new_n216), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n254), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n637), .B1(new_n638), .B2(new_n216), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n633), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(KEYINPUT103), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n637), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n216), .B1(new_n251), .B2(new_n253), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n216), .A2(KEYINPUT10), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n645), .A2(new_n650), .B1(new_n258), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n643), .B1(new_n652), .B2(new_n642), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n641), .B(KEYINPUT105), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n656), .B1(new_n642), .B2(new_n640), .ZN(new_n657));
  INV_X1    g456(.A(new_n633), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n607), .A2(new_n629), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(new_n557), .A3(new_n558), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n546), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT106), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT16), .B(G8gat), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n665), .A2(new_n664), .A3(new_n667), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n669), .B1(new_n666), .B2(G8gat), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(G1325gat));
  NOR2_X1   g470(.A1(new_n604), .A2(new_n605), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n661), .A2(G15gat), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n410), .ZN(new_n674));
  INV_X1    g473(.A(new_n416), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n661), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n677), .A2(G15gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n673), .B1(new_n678), .B2(KEYINPUT107), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(KEYINPUT107), .B2(new_n678), .ZN(G1326gat));
  NAND2_X1  g479(.A1(new_n661), .A2(new_n598), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NAND2_X1  g482(.A1(new_n562), .A2(new_n606), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n660), .A2(new_n229), .A3(new_n629), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n290), .A3(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n687), .A2(G29gat), .A3(new_n559), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT45), .Z(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n684), .B2(new_n290), .ZN(new_n691));
  AOI211_X1 g490(.A(KEYINPUT44), .B(new_n289), .C1(new_n562), .C2(new_n606), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n686), .ZN(new_n694));
  OAI21_X1  g493(.A(G29gat), .B1(new_n694), .B2(new_n559), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n689), .A2(new_n695), .ZN(G1328gat));
  OAI21_X1  g495(.A(G36gat), .B1(new_n694), .B2(new_n545), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n687), .A2(G36gat), .A3(new_n545), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT46), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(G1329gat));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n701));
  INV_X1    g500(.A(new_n676), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n687), .A2(G43gat), .A3(new_n702), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT109), .Z(new_n704));
  INV_X1    g503(.A(new_n672), .ZN(new_n705));
  OAI21_X1  g504(.A(G43gat), .B1(new_n694), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n701), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n598), .B(new_n686), .C1(new_n691), .C2(new_n692), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n710), .A2(G50gat), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n687), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n464), .A2(G50gat), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n289), .B1(new_n562), .B2(new_n606), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(KEYINPUT110), .A3(new_n686), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n709), .B1(new_n711), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n714), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n687), .B2(new_n712), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n722), .A2(KEYINPUT111), .A3(new_n717), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT111), .B1(new_n722), .B2(new_n717), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n709), .B1(new_n710), .B2(G50gat), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT112), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n715), .B2(new_n718), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n722), .A2(KEYINPUT111), .A3(new_n717), .ZN(new_n730));
  AND4_X1   g529(.A1(KEYINPUT112), .A2(new_n726), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n720), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT113), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT113), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n734), .B(new_n720), .C1(new_n727), .C2(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(G1331gat));
  NOR2_X1   g535(.A1(new_n660), .A2(new_n629), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n607), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(new_n559), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g539(.A(new_n738), .B(KEYINPUT114), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n546), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT49), .B(G64gat), .Z(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(G1333gat));
  NOR3_X1   g544(.A1(new_n738), .A2(G71gat), .A3(new_n702), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n741), .A2(new_n672), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n747), .B2(G71gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n741), .A2(new_n598), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g550(.A1(new_n693), .A2(new_n229), .A3(new_n737), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n752), .A2(new_n559), .A3(new_n240), .ZN(new_n753));
  INV_X1    g552(.A(new_n629), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n716), .A2(new_n229), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n660), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(new_n557), .A3(new_n558), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n753), .B1(new_n240), .B2(new_n760), .ZN(G1336gat));
  NAND2_X1  g560(.A1(new_n757), .A2(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n659), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n241), .B1(new_n763), .B2(new_n545), .ZN(new_n764));
  INV_X1    g563(.A(new_n752), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(G92gat), .A3(new_n546), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(G1337gat));
  OR3_X1    g568(.A1(new_n763), .A2(G99gat), .A3(new_n702), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n765), .A2(new_n672), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n771), .A2(KEYINPUT115), .ZN(new_n772));
  OAI21_X1  g571(.A(G99gat), .B1(new_n771), .B2(KEYINPUT115), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(G1338gat));
  INV_X1    g573(.A(G106gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n775), .A3(new_n598), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n693), .A2(new_n598), .A3(new_n229), .A4(new_n737), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G106gat), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n778), .A2(KEYINPUT116), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n779), .A2(new_n780), .A3(KEYINPUT53), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n776), .B(new_n778), .C1(KEYINPUT116), .C2(KEYINPUT53), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n781), .A2(new_n783), .ZN(G1339gat));
  INV_X1    g583(.A(new_n229), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n658), .B1(new_n656), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n645), .A2(new_n650), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n258), .A2(new_n651), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n655), .A3(new_n789), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n790), .B(KEYINPUT54), .C1(new_n642), .C2(new_n652), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT118), .ZN(new_n795));
  INV_X1    g594(.A(new_n628), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n609), .B1(new_n608), .B2(new_n610), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n797), .A2(KEYINPUT119), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n616), .A2(new_n617), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n797), .B2(KEYINPUT119), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n624), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT120), .B1(new_n796), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n798), .A2(new_n800), .ZN(new_n803));
  INV_X1    g602(.A(new_n624), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n806), .A3(new_n628), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(new_n286), .A3(new_n288), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n791), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(new_n653), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT55), .B1(new_n787), .B2(new_n791), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n795), .A2(new_n810), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT121), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n653), .B(new_n811), .C1(new_n813), .C2(new_n814), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT121), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n819), .A2(new_n820), .A3(new_n815), .A4(new_n810), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n795), .A2(new_n812), .A3(new_n629), .A4(new_n815), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n659), .A2(new_n628), .A3(new_n805), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n289), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n785), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n289), .A2(new_n785), .A3(new_n754), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n828), .A2(new_n659), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OR3_X1    g630(.A1(new_n828), .A2(new_n830), .A3(new_n659), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n827), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n559), .A2(new_n546), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n465), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n754), .ZN(new_n838));
  INV_X1    g637(.A(new_n555), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(new_n839), .A3(new_n836), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n629), .A2(new_n357), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(G1340gat));
  OAI21_X1  g641(.A(G120gat), .B1(new_n837), .B2(new_n660), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n659), .A2(new_n360), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n840), .B2(new_n844), .ZN(G1341gat));
  OAI21_X1  g644(.A(G127gat), .B1(new_n837), .B2(new_n229), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n229), .A2(G127gat), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n835), .A2(new_n839), .A3(new_n836), .A4(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n847), .B1(new_n846), .B2(new_n849), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(G1342gat));
  NAND2_X1  g651(.A1(new_n290), .A2(new_n364), .ZN(new_n853));
  OR3_X1    g652(.A1(new_n840), .A2(KEYINPUT56), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G134gat), .B1(new_n837), .B2(new_n289), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT56), .B1(new_n840), .B2(new_n853), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(G1343gat));
  NAND3_X1  g656(.A1(new_n812), .A2(new_n629), .A3(new_n794), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n824), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n289), .ZN(new_n860));
  AOI211_X1 g659(.A(KEYINPUT118), .B(KEYINPUT55), .C1(new_n787), .C2(new_n791), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n818), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n820), .B1(new_n862), .B2(new_n810), .ZN(new_n863));
  NOR4_X1   g662(.A1(new_n818), .A2(new_n809), .A3(new_n861), .A4(KEYINPUT121), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n833), .B1(new_n865), .B2(new_n229), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT57), .B1(new_n866), .B2(new_n464), .ZN(new_n867));
  OR3_X1    g666(.A1(new_n672), .A2(new_n559), .A3(new_n546), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n870), .B(new_n598), .C1(new_n827), .C2(new_n833), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n867), .A2(new_n629), .A3(new_n869), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(G141gat), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n834), .A2(new_n464), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n874), .A2(new_n417), .A3(new_n629), .A4(new_n869), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT58), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n873), .A2(new_n878), .A3(new_n875), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(G1344gat));
  NAND2_X1  g679(.A1(new_n874), .A2(new_n869), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n659), .A2(new_n419), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(KEYINPUT123), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n881), .A2(new_n885), .A3(new_n882), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT57), .B1(new_n834), .B2(new_n464), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n785), .B1(new_n860), .B2(new_n816), .ZN(new_n889));
  INV_X1    g688(.A(new_n829), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n870), .B(new_n598), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n888), .A2(new_n659), .A3(new_n869), .A4(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n887), .B1(new_n892), .B2(G148gat), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n887), .A2(G148gat), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n867), .A2(new_n869), .A3(new_n871), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n659), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n884), .A2(new_n886), .B1(new_n893), .B2(new_n896), .ZN(G1345gat));
  INV_X1    g696(.A(G155gat), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n229), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n874), .A2(new_n785), .A3(new_n869), .ZN(new_n900));
  AOI22_X1  g699(.A1(new_n895), .A2(new_n899), .B1(new_n900), .B2(new_n898), .ZN(G1346gat));
  NAND4_X1  g700(.A1(new_n867), .A2(new_n290), .A3(new_n869), .A4(new_n871), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G162gat), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n289), .A2(G162gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n874), .A2(new_n869), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n903), .A2(KEYINPUT124), .A3(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1347gat));
  AND2_X1   g709(.A1(new_n465), .A2(new_n546), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n911), .B(new_n559), .C1(new_n827), .C2(new_n833), .ZN(new_n912));
  OAI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n754), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n545), .B1(new_n557), .B2(new_n558), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n839), .B(new_n914), .C1(new_n827), .C2(new_n833), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n629), .A2(new_n305), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(G1348gat));
  NOR3_X1   g716(.A1(new_n912), .A2(new_n306), .A3(new_n660), .ZN(new_n918));
  INV_X1    g717(.A(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n659), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n918), .B1(new_n306), .B2(new_n920), .ZN(G1349gat));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n313), .A2(new_n314), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n785), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n919), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT125), .B1(new_n915), .B2(new_n924), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G183gat), .B1(new_n912), .B2(new_n229), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT60), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n932), .A3(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1350gat));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n935), .B(G190gat), .C1(new_n912), .C2(new_n289), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n936), .A2(KEYINPUT126), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(KEYINPUT126), .ZN(new_n938));
  OAI21_X1  g737(.A(G190gat), .B1(new_n912), .B2(new_n289), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n919), .A2(new_n322), .A3(new_n290), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1351gat));
  AND2_X1   g742(.A1(new_n888), .A2(new_n891), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n705), .A2(new_n914), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n629), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G197gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n834), .B1(new_n557), .B2(new_n558), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n705), .A2(new_n546), .A3(new_n598), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT127), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n949), .A2(new_n621), .A3(new_n629), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n948), .A2(new_n952), .ZN(G1352gat));
  NOR2_X1   g752(.A1(new_n660), .A2(G204gat), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n835), .A2(new_n559), .A3(new_n951), .A4(new_n954), .ZN(new_n955));
  XOR2_X1   g754(.A(new_n955), .B(KEYINPUT62), .Z(new_n956));
  NAND3_X1  g755(.A1(new_n944), .A2(new_n659), .A3(new_n946), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G204gat), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1353gat));
  NOR2_X1   g758(.A1(new_n229), .A2(new_n428), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n949), .A2(new_n951), .A3(new_n960), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n888), .A2(new_n785), .A3(new_n891), .A4(new_n946), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  AND2_X1   g764(.A1(new_n944), .A2(new_n946), .ZN(new_n966));
  INV_X1    g765(.A(G218gat), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n289), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n949), .A2(new_n290), .A3(new_n951), .ZN(new_n969));
  AOI22_X1  g768(.A1(new_n966), .A2(new_n968), .B1(new_n967), .B2(new_n969), .ZN(G1355gat));
endmodule


