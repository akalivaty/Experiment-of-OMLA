//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G228gat), .A2(G233gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  AND2_X1   g007(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n209));
  NOR2_X1   g008(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT76), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g012(.A(KEYINPUT76), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n214));
  XOR2_X1   g013(.A(G141gat), .B(G148gat), .Z(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(KEYINPUT74), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT74), .ZN(new_n219));
  NOR3_X1   g018(.A1(new_n219), .A2(G155gat), .A3(G162gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n208), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(new_n217), .ZN(new_n225));
  XNOR2_X1  g024(.A(G141gat), .B(G148gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT77), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n217), .A2(new_n224), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n208), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT77), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(new_n215), .A3(new_n230), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n216), .A2(new_n222), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G211gat), .B(G218gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT22), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT70), .B(G211gat), .ZN(new_n235));
  INV_X1    g034(.A(G218gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(G197gat), .B(G204gat), .Z(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n233), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT29), .B1(new_n240), .B2(KEYINPUT79), .ZN(new_n241));
  INV_X1    g040(.A(new_n233), .ZN(new_n242));
  INV_X1    g041(.A(G211gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT70), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G211gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT22), .B1(new_n247), .B2(G218gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n242), .B1(new_n248), .B2(new_n238), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT79), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n237), .A2(new_n233), .A3(new_n239), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n241), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n232), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n249), .A2(new_n251), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n216), .A2(new_n222), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n227), .A2(new_n231), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT29), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n207), .B1(new_n255), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT80), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT80), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n264), .B(new_n207), .C1(new_n255), .C2(new_n261), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n207), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT3), .B1(new_n256), .B2(new_n260), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n267), .B1(new_n268), .B2(new_n232), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n259), .A2(new_n260), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT81), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n256), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT29), .B1(new_n232), .B2(new_n254), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT81), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n269), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n206), .B1(new_n266), .B2(new_n276), .ZN(new_n277));
  AOI211_X1 g076(.A(G22gat), .B(new_n275), .C1(new_n263), .C2(new_n265), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n205), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n265), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT3), .B1(new_n241), .B2(new_n252), .ZN(new_n281));
  OAI22_X1  g080(.A1(new_n281), .A2(new_n232), .B1(new_n273), .B2(new_n256), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n264), .B1(new_n282), .B2(new_n207), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n276), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G22gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n266), .A2(new_n206), .A3(new_n276), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(new_n204), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n288));
  INV_X1    g087(.A(G183gat), .ZN(new_n289));
  INV_X1    g088(.A(G190gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT64), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(G183gat), .A3(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT24), .B1(new_n296), .B2(KEYINPUT64), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n293), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G169gat), .ZN(new_n299));
  INV_X1    g098(.A(G176gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT23), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT23), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n302), .B1(G169gat), .B2(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT25), .B1(new_n298), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT65), .ZN(new_n308));
  OR3_X1    g107(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT65), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n310), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n308), .A2(new_n309), .A3(new_n311), .A4(new_n304), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n289), .A2(KEYINPUT27), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT27), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G183gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n315), .A3(new_n290), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT28), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT27), .B(G183gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT28), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n319), .A3(new_n290), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n312), .A2(new_n317), .A3(new_n320), .A4(new_n296), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n305), .A2(KEYINPUT25), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n293), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n306), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G120gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G113gat), .ZN(new_n328));
  INV_X1    g127(.A(G113gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G120gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n331), .A2(KEYINPUT66), .ZN(new_n332));
  XNOR2_X1  g131(.A(G127gat), .B(G134gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n329), .A2(KEYINPUT66), .A3(G120gat), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n331), .A2(new_n334), .ZN(new_n338));
  INV_X1    g137(.A(new_n333), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n288), .B1(new_n326), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n305), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n297), .A2(new_n295), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(new_n293), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n345), .A2(KEYINPUT25), .B1(new_n324), .B2(new_n322), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n332), .A2(new_n336), .B1(new_n338), .B2(new_n339), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n346), .A2(KEYINPUT67), .A3(new_n347), .A4(new_n321), .ZN(new_n348));
  NAND2_X1  g147(.A1(G227gat), .A2(G233gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n326), .A2(new_n341), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n342), .A2(new_n348), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n351), .B(KEYINPUT34), .Z(new_n352));
  INV_X1    g151(.A(KEYINPUT32), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n342), .A2(new_n348), .A3(new_n350), .ZN(new_n354));
  INV_X1    g153(.A(new_n349), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G15gat), .B(G43gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(KEYINPUT69), .ZN(new_n358));
  XNOR2_X1  g157(.A(G71gat), .B(G99gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT33), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(KEYINPUT68), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n354), .A2(new_n355), .A3(new_n360), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT68), .B1(new_n364), .B2(new_n361), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n352), .B(new_n363), .C1(new_n365), .C2(new_n356), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n363), .B1(new_n365), .B2(new_n356), .ZN(new_n367));
  INV_X1    g166(.A(new_n352), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n279), .A2(new_n287), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT35), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n227), .A2(new_n231), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n226), .B1(new_n211), .B2(new_n212), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n221), .B1(new_n373), .B2(new_n214), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT3), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(new_n259), .A3(new_n341), .ZN(new_n376));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n257), .A2(new_n347), .A3(new_n258), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n232), .A2(KEYINPUT4), .A3(new_n347), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n376), .A2(new_n377), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n341), .B1(new_n372), .B2(new_n374), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n378), .ZN(new_n385));
  INV_X1    g184(.A(new_n377), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n232), .A2(KEYINPUT4), .A3(new_n347), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT4), .B1(new_n232), .B2(new_n347), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n391), .A2(new_n383), .A3(new_n377), .A4(new_n376), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G1gat), .B(G29gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT0), .ZN(new_n395));
  XNOR2_X1  g194(.A(G57gat), .B(G85gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n388), .A2(new_n392), .A3(new_n397), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n393), .A2(KEYINPUT6), .A3(new_n398), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT72), .ZN(new_n405));
  NAND2_X1  g204(.A1(G226gat), .A2(G233gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n406), .B(KEYINPUT71), .Z(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(KEYINPUT29), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n326), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n306), .A2(new_n321), .A3(new_n325), .A4(new_n407), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n256), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n256), .B1(new_n409), .B2(new_n410), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n405), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n409), .A2(new_n410), .ZN(new_n415));
  INV_X1    g214(.A(new_n256), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(KEYINPUT72), .A3(new_n411), .ZN(new_n418));
  XNOR2_X1  g217(.A(G8gat), .B(G36gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(G64gat), .B(G92gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n414), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n417), .A2(new_n411), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(KEYINPUT30), .A3(new_n421), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n412), .A2(new_n413), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n422), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n429), .A2(KEYINPUT30), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n370), .A2(new_n371), .A3(new_n404), .A4(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT78), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n402), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n399), .A2(KEYINPUT78), .A3(new_n400), .A4(new_n401), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n403), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT73), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n426), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n423), .A2(KEYINPUT73), .A3(new_n425), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n440), .A2(new_n441), .A3(new_n430), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n369), .A2(new_n366), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n285), .A2(new_n286), .A3(new_n204), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n204), .B1(new_n285), .B2(new_n286), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT35), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT86), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n279), .A2(new_n287), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n451), .A2(new_n438), .A3(new_n442), .A4(new_n444), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n434), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n384), .A2(new_n378), .A3(new_n377), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n456), .B(KEYINPUT83), .Z(new_n457));
  AOI21_X1  g256(.A(new_n377), .B1(new_n391), .B2(new_n376), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n459), .A3(KEYINPUT39), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT82), .B(KEYINPUT39), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n398), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n455), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT40), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n464), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n465), .A2(new_n466), .A3(new_n399), .A4(new_n431), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n414), .A2(new_n418), .A3(KEYINPUT37), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n422), .B1(new_n428), .B2(KEYINPUT37), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT38), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT85), .ZN(new_n471));
  OR2_X1    g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n404), .ZN(new_n473));
  INV_X1    g272(.A(new_n469), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT38), .B1(new_n428), .B2(KEYINPUT37), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n429), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n470), .A2(new_n471), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n472), .A2(new_n473), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n467), .A2(new_n478), .A3(new_n451), .ZN(new_n479));
  INV_X1    g278(.A(new_n451), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n443), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n444), .B(KEYINPUT36), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n454), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT16), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n485), .B1(new_n486), .B2(G1gat), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(G1gat), .B2(new_n485), .ZN(new_n488));
  INV_X1    g287(.A(G8gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  OR3_X1    g290(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT88), .B(G29gat), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n493), .A2(G36gat), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G43gat), .B(G50gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(KEYINPUT89), .A3(KEYINPUT15), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n499));
  XOR2_X1   g298(.A(KEYINPUT90), .B(G43gat), .Z(new_n500));
  OAI21_X1  g299(.A(new_n499), .B1(new_n500), .B2(G50gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n497), .A2(KEYINPUT15), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT89), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n496), .A2(new_n498), .A3(new_n501), .A4(new_n504), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n492), .A2(KEYINPUT87), .ZN(new_n506));
  INV_X1    g305(.A(new_n495), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n492), .B2(KEYINPUT87), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n506), .A2(new_n508), .B1(G36gat), .B2(new_n493), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n505), .B1(new_n502), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n491), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(KEYINPUT17), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(new_n490), .ZN(new_n513));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT18), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n513), .A2(KEYINPUT18), .A3(new_n514), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n491), .B(new_n510), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n514), .B(KEYINPUT13), .Z(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G113gat), .B(G141gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(G197gat), .ZN(new_n524));
  XOR2_X1   g323(.A(KEYINPUT11), .B(G169gat), .Z(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n526), .B(KEYINPUT12), .Z(new_n527));
  OR2_X1    g326(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n522), .A2(new_n527), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n484), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G57gat), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n533), .A2(G64gat), .ZN(new_n534));
  INV_X1    g333(.A(G64gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(G57gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT91), .ZN(new_n537));
  OAI22_X1  g336(.A1(new_n534), .A2(new_n536), .B1(new_n537), .B2(KEYINPUT9), .ZN(new_n538));
  NOR2_X1   g337(.A1(G71gat), .A2(G78gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(G71gat), .A2(G78gat), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n539), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n538), .B(new_n541), .C1(new_n537), .C2(new_n540), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(KEYINPUT9), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n540), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT92), .B1(new_n533), .B2(G64gat), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(G57gat), .B2(new_n535), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n533), .A2(KEYINPUT92), .A3(G64gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n542), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n549), .A2(KEYINPUT21), .ZN(new_n550));
  NAND2_X1  g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G127gat), .B(G155gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT93), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n552), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G183gat), .B(G211gat), .Z(new_n556));
  XOR2_X1   g355(.A(new_n555), .B(new_n556), .Z(new_n557));
  AOI21_X1  g356(.A(new_n491), .B1(KEYINPUT21), .B2(new_n549), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n557), .B(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G99gat), .ZN(new_n563));
  INV_X1    g362(.A(G106gat), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT8), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT96), .B(G92gat), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n565), .B1(new_n566), .B2(G85gat), .ZN(new_n567));
  XOR2_X1   g366(.A(G99gat), .B(G106gat), .Z(new_n568));
  AOI21_X1  g367(.A(new_n567), .B1(KEYINPUT97), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT7), .ZN(new_n570));
  OAI211_X1 g369(.A(G85gat), .B(G92gat), .C1(new_n570), .C2(KEYINPUT94), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT94), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(KEYINPUT7), .ZN(new_n573));
  OR3_X1    g372(.A1(new_n571), .A2(KEYINPUT95), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT95), .B1(new_n571), .B2(new_n573), .ZN(new_n575));
  INV_X1    g374(.A(G85gat), .ZN(new_n576));
  INV_X1    g375(.A(G92gat), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT7), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n569), .A2(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n568), .A2(KEYINPUT97), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n512), .A2(new_n582), .ZN(new_n583));
  AND3_X1   g382(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n584));
  INV_X1    g383(.A(new_n582), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(new_n510), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G190gat), .B(G218gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n583), .A2(new_n588), .A3(new_n586), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT98), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n593));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n592), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n593), .B1(new_n592), .B2(new_n596), .ZN(new_n598));
  OR3_X1    g397(.A1(new_n590), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n590), .B1(new_n597), .B2(new_n598), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n562), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n585), .A2(new_n549), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n585), .A2(new_n549), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n585), .A2(KEYINPUT10), .A3(new_n549), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n604), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n603), .B1(new_n605), .B2(new_n607), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G120gat), .B(G148gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(G176gat), .B(G204gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n613), .B(new_n614), .Z(new_n615));
  NOR2_X1   g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n615), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT100), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n612), .A2(KEYINPUT100), .A3(new_n615), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n602), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n532), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n438), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g427(.A(new_n489), .B1(new_n625), .B2(new_n431), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT16), .B(G8gat), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n624), .A2(new_n432), .A3(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT42), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n632), .B1(KEYINPUT42), .B2(new_n631), .ZN(G1325gat));
  INV_X1    g432(.A(new_n444), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n624), .A2(G15gat), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n482), .B(KEYINPUT101), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n625), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n635), .B1(G15gat), .B2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT102), .Z(G1326gat));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n451), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT43), .B(G22gat), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(G1327gat));
  NAND2_X1  g442(.A1(new_n621), .A2(new_n561), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n601), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n532), .A2(new_n645), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n646), .A2(new_n438), .A3(new_n493), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n647), .B(KEYINPUT45), .Z(new_n648));
  INV_X1    g447(.A(new_n601), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n649), .A2(KEYINPUT44), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n650), .B1(new_n454), .B2(new_n483), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n644), .A2(new_n531), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n440), .A2(new_n441), .A3(new_n430), .ZN(new_n653));
  INV_X1    g452(.A(new_n403), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n654), .B1(new_n402), .B2(new_n435), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n653), .B1(new_n655), .B2(new_n437), .ZN(new_n656));
  AOI211_X1 g455(.A(new_n449), .B(new_n371), .C1(new_n656), .C2(new_n370), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT86), .B1(new_n452), .B2(KEYINPUT35), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n433), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n481), .A2(KEYINPUT103), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n443), .A2(new_n480), .A3(new_n661), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n660), .A2(new_n482), .A3(new_n479), .A4(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n601), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n651), .B(new_n652), .C1(new_n664), .C2(KEYINPUT44), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n666), .A2(KEYINPUT104), .A3(new_n626), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(new_n665), .B2(new_n438), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n667), .A2(new_n493), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n648), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT105), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n648), .A2(new_n673), .A3(new_n670), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(G1328gat));
  NOR3_X1   g474(.A1(new_n646), .A2(G36gat), .A3(new_n432), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G36gat), .B1(new_n665), .B2(new_n432), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(G1329gat));
  OR3_X1    g479(.A1(new_n665), .A2(KEYINPUT108), .A3(new_n482), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT108), .B1(new_n665), .B2(new_n482), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(new_n500), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n646), .ZN(new_n684));
  INV_X1    g483(.A(new_n500), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(new_n444), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n683), .A2(KEYINPUT47), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(KEYINPUT107), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n685), .B1(new_n666), .B2(new_n637), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n687), .B1(new_n690), .B2(KEYINPUT47), .ZN(G1330gat));
  OR2_X1    g490(.A1(new_n684), .A2(KEYINPUT109), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n684), .A2(KEYINPUT109), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n451), .A2(G50gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(G50gat), .B1(new_n665), .B2(new_n451), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT48), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n697), .B(new_n699), .ZN(G1331gat));
  NAND2_X1  g499(.A1(new_n659), .A2(new_n663), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n602), .A2(new_n530), .A3(new_n621), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n626), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g504(.A(new_n432), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT111), .ZN(new_n708));
  NOR2_X1   g507(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1333gat));
  AND2_X1   g509(.A1(new_n703), .A2(new_n444), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n711), .A2(KEYINPUT112), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(KEYINPUT112), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n712), .A2(new_n713), .A3(G71gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n703), .A2(G71gat), .A3(new_n637), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g516(.A1(new_n703), .A2(new_n480), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g518(.A1(new_n531), .A2(new_n561), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT113), .B1(new_n720), .B2(new_n621), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT113), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n622), .A2(new_n531), .A3(new_n722), .A4(new_n561), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n651), .B(new_n724), .C1(new_n664), .C2(KEYINPUT44), .ZN(new_n725));
  OAI21_X1  g524(.A(G85gat), .B1(new_n725), .B2(new_n438), .ZN(new_n726));
  INV_X1    g525(.A(new_n720), .ZN(new_n727));
  AND4_X1   g526(.A1(KEYINPUT51), .A2(new_n701), .A3(new_n649), .A4(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT51), .B1(new_n664), .B2(new_n727), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n622), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n626), .A2(new_n576), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n726), .B1(new_n731), .B2(new_n732), .ZN(G1336gat));
  OAI21_X1  g532(.A(new_n566), .B1(new_n725), .B2(new_n432), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n431), .A2(new_n577), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n731), .B2(new_n735), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1337gat));
  NOR3_X1   g537(.A1(new_n621), .A2(G99gat), .A3(new_n634), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT115), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n730), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G99gat), .B1(new_n725), .B2(new_n636), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1338gat));
  INV_X1    g542(.A(KEYINPUT119), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n451), .A2(G106gat), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n622), .B(new_n745), .C1(new_n728), .C2(new_n729), .ZN(new_n746));
  OAI21_X1  g545(.A(G106gat), .B1(new_n725), .B2(new_n451), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT116), .B1(new_n748), .B2(KEYINPUT53), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT116), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751));
  AOI211_X1 g550(.A(new_n750), .B(new_n751), .C1(new_n746), .C2(new_n747), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n754));
  NAND3_X1  g553(.A1(new_n746), .A2(new_n747), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT118), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT118), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n746), .A2(new_n747), .A3(new_n757), .A4(new_n754), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n744), .B1(new_n753), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n758), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n761), .B(KEYINPUT119), .C1(new_n749), .C2(new_n752), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(G1339gat));
  NOR2_X1   g562(.A1(new_n513), .A2(new_n514), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n519), .A2(new_n520), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n526), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n528), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n649), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n601), .A2(new_n531), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n619), .A2(new_n620), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT54), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n610), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n608), .A2(new_n609), .A3(new_n604), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n615), .B1(new_n610), .B2(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT55), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n768), .A2(new_n769), .A3(new_n770), .A4(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n622), .A2(new_n528), .A3(new_n601), .A4(new_n766), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n562), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n602), .A2(new_n622), .A3(new_n530), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n438), .A2(new_n431), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n370), .A3(new_n784), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n785), .A2(new_n329), .A3(new_n531), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n782), .A2(new_n438), .A3(new_n431), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n370), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n530), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n786), .B1(new_n790), .B2(new_n329), .ZN(G1340gat));
  NOR3_X1   g590(.A1(new_n785), .A2(new_n327), .A3(new_n621), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n622), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n793), .B2(new_n327), .ZN(G1341gat));
  OAI21_X1  g593(.A(G127gat), .B1(new_n785), .B2(new_n561), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n561), .A2(G127gat), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(new_n788), .B2(new_n796), .ZN(G1342gat));
  OR4_X1    g596(.A1(KEYINPUT56), .A2(new_n788), .A3(G134gat), .A4(new_n601), .ZN(new_n798));
  OAI21_X1  g597(.A(G134gat), .B1(new_n785), .B2(new_n601), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n601), .A2(G134gat), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT56), .B1(new_n788), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(G1343gat));
  NOR2_X1   g601(.A1(new_n637), .A2(new_n451), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n783), .A2(new_n784), .A3(new_n803), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n531), .A2(G141gat), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n782), .B2(new_n451), .ZN(new_n808));
  OAI211_X1 g607(.A(KEYINPUT57), .B(new_n480), .C1(new_n780), .C2(new_n781), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n482), .A2(new_n784), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n530), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n806), .B1(new_n813), .B2(G141gat), .ZN(new_n814));
  XOR2_X1   g613(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n815));
  XNOR2_X1  g614(.A(new_n814), .B(new_n815), .ZN(G1344gat));
  NOR3_X1   g615(.A1(new_n804), .A2(G148gat), .A3(new_n621), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT121), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n810), .A2(new_n622), .A3(new_n812), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(G148gat), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(new_n822), .A3(new_n823), .ZN(G1345gat));
  INV_X1    g623(.A(new_n804), .ZN(new_n825));
  INV_X1    g624(.A(G155gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n826), .A3(new_n562), .ZN(new_n827));
  INV_X1    g626(.A(new_n810), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n828), .A2(new_n561), .A3(new_n811), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n829), .B2(new_n826), .ZN(G1346gat));
  AOI21_X1  g629(.A(G162gat), .B1(new_n825), .B2(new_n649), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n828), .A2(new_n811), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n649), .A2(G162gat), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(G1347gat));
  NOR2_X1   g633(.A1(new_n626), .A2(new_n432), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n783), .A2(new_n370), .A3(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n836), .A2(new_n299), .A3(new_n531), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n782), .A2(new_n626), .A3(new_n432), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n370), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n530), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n837), .B1(new_n841), .B2(new_n299), .ZN(G1348gat));
  NOR3_X1   g641(.A1(new_n836), .A2(new_n300), .A3(new_n621), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n300), .B1(new_n839), .B2(new_n621), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n843), .B1(new_n846), .B2(new_n847), .ZN(G1349gat));
  OAI21_X1  g647(.A(G183gat), .B1(new_n836), .B2(new_n561), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n838), .A2(new_n318), .A3(new_n370), .A4(new_n562), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT60), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n849), .A2(new_n850), .B1(KEYINPUT123), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n851), .A2(KEYINPUT123), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n852), .B(new_n853), .ZN(G1350gat));
  OAI21_X1  g653(.A(G190gat), .B1(new_n836), .B2(new_n601), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT61), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n840), .A2(new_n290), .A3(new_n649), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1351gat));
  NAND3_X1  g657(.A1(new_n783), .A2(new_n803), .A3(new_n835), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(G197gat), .B1(new_n860), .B2(new_n530), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n636), .A2(new_n835), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n862), .B1(new_n808), .B2(new_n809), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n530), .A2(G197gat), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(G1352gat));
  INV_X1    g664(.A(G204gat), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n863), .A2(new_n622), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(KEYINPUT125), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(KEYINPUT125), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n621), .A2(G204gat), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT124), .B1(new_n859), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n838), .A2(new_n873), .A3(new_n803), .A4(new_n870), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n872), .A2(new_n874), .A3(KEYINPUT62), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT62), .B1(new_n872), .B2(new_n874), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n869), .A2(new_n877), .ZN(G1353gat));
  NAND3_X1  g677(.A1(new_n860), .A2(new_n235), .A3(new_n562), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n562), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(KEYINPUT126), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n243), .B1(KEYINPUT126), .B2(new_n881), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n882), .B1(new_n880), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(G1354gat));
  INV_X1    g685(.A(KEYINPUT127), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n863), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n649), .B1(new_n863), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g688(.A(G218gat), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n860), .A2(new_n236), .A3(new_n649), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1355gat));
endmodule


