//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1243,
    new_n1244, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0002(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT66), .ZN(new_n204));
  AOI22_X1  g0004(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n207));
  AND3_X1   g0007(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(new_n204), .A2(new_n208), .B1(G1), .B2(G20), .ZN(new_n209));
  INV_X1    g0009(.A(KEYINPUT1), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G20), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT65), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n209), .A2(new_n210), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT64), .Z(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT0), .ZN(new_n221));
  AOI211_X1 g0021(.A(new_n216), .B(new_n221), .C1(new_n210), .C2(new_n209), .ZN(G361));
  XNOR2_X1  g0022(.A(G238), .B(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT2), .B(G226), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G250), .B(G257), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G264), .B(G270), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n227), .B(new_n230), .ZN(G358));
  XNOR2_X1  g0031(.A(G68), .B(G77), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT67), .ZN(new_n233));
  XOR2_X1   g0033(.A(G50), .B(G58), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G97), .B(G107), .Z(new_n236));
  XNOR2_X1  g0036(.A(G87), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G351));
  NOR2_X1   g0039(.A1(G20), .A2(G33), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G150), .ZN(new_n241));
  INV_X1    g0041(.A(G50), .ZN(new_n242));
  INV_X1    g0042(.A(G58), .ZN(new_n243));
  INV_X1    g0043(.A(G68), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G20), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT8), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n247), .B1(new_n243), .B2(KEYINPUT69), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT69), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(KEYINPUT8), .A3(G58), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n241), .B(new_n246), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT68), .B1(new_n217), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT68), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n257), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(new_n211), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n254), .A2(KEYINPUT70), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n242), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n254), .A2(new_n259), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT70), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n259), .A2(new_n263), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n261), .A2(G20), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(G50), .A3(new_n269), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n260), .A2(new_n264), .A3(new_n267), .A4(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT9), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n212), .B1(new_n255), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G226), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  NOR3_X1   g0079(.A1(new_n278), .A2(new_n279), .A3(new_n275), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G222), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n285), .B1(new_n286), .B2(new_n283), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n282), .B1(new_n289), .B2(new_n278), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G190), .ZN(new_n291));
  INV_X1    g0091(.A(G200), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n272), .B(new_n291), .C1(new_n292), .C2(new_n290), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT10), .ZN(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g0096(.A(new_n296), .B(KEYINPUT71), .Z(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(new_n271), .C1(G169), .C2(new_n290), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n240), .A2(G50), .B1(G20), .B2(new_n244), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n286), .B2(new_n253), .ZN(new_n301));
  AOI21_X1  g0101(.A(KEYINPUT11), .B1(new_n301), .B2(new_n259), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n262), .A2(G68), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT12), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n301), .A2(KEYINPUT11), .A3(new_n259), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n268), .A2(G68), .A3(new_n269), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT14), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n283), .A2(G232), .A3(G1698), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n283), .A2(G226), .A3(new_n284), .ZN(new_n311));
  INV_X1    g0111(.A(G97), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n310), .B(new_n311), .C1(new_n255), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n278), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT13), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n280), .B1(new_n276), .B2(G238), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n315), .B1(new_n314), .B2(new_n316), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n309), .B(G169), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n318), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n319), .B1(new_n322), .B2(new_n295), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n309), .B1(new_n322), .B2(G169), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n308), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G20), .A2(G77), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT15), .B(G87), .ZN(new_n328));
  INV_X1    g0128(.A(new_n240), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT8), .B(G58), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n327), .B1(new_n328), .B2(new_n253), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n331), .A2(new_n259), .B1(new_n286), .B2(new_n263), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n268), .A2(G77), .A3(new_n269), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G238), .ZN(new_n335));
  INV_X1    g0135(.A(G107), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n287), .A2(new_n335), .B1(new_n336), .B2(new_n283), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT3), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G33), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n341), .A2(new_n224), .A3(G1698), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n278), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n280), .B1(new_n276), .B2(G244), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n334), .B1(G200), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G190), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(new_n345), .ZN(new_n348));
  INV_X1    g0148(.A(G169), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n343), .A2(new_n295), .A3(new_n344), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(new_n334), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT72), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n317), .A2(new_n318), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n308), .B1(new_n355), .B2(G190), .ZN(new_n356));
  OAI21_X1  g0156(.A(G200), .B1(new_n317), .B2(new_n318), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n320), .A2(G190), .A3(new_n321), .ZN(new_n359));
  INV_X1    g0159(.A(new_n308), .ZN(new_n360));
  AND4_X1   g0160(.A1(new_n354), .A2(new_n359), .A3(new_n360), .A4(new_n357), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NOR4_X1   g0162(.A1(new_n299), .A2(new_n326), .A3(new_n353), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n276), .A2(G232), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n281), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n338), .A2(new_n340), .A3(G223), .A4(new_n284), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G33), .A2(G87), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(G226), .A2(G1698), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n338), .A2(new_n340), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT74), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n283), .A2(KEYINPUT74), .A3(new_n370), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n369), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n278), .B1(new_n375), .B2(KEYINPUT75), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT74), .B1(new_n283), .B2(new_n370), .ZN(new_n377));
  AND4_X1   g0177(.A1(KEYINPUT74), .A2(new_n338), .A3(new_n340), .A4(new_n370), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n368), .B(new_n367), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT75), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n347), .B(new_n366), .C1(new_n376), .C2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n274), .B1(new_n379), .B2(new_n380), .ZN(new_n383));
  INV_X1    g0183(.A(new_n369), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n384), .B(KEYINPUT75), .C1(new_n377), .C2(new_n378), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n365), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n382), .B(KEYINPUT77), .C1(G200), .C2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n251), .B1(new_n261), .B2(G20), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n268), .A2(new_n388), .B1(new_n263), .B2(new_n251), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT16), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n283), .B2(G20), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n341), .A2(KEYINPUT7), .A3(new_n252), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT73), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT73), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n396), .B(new_n392), .C1(new_n283), .C2(G20), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n395), .A2(G68), .A3(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n243), .A2(new_n244), .ZN(new_n399));
  NOR2_X1   g0199(.A1(G58), .A2(G68), .ZN(new_n400));
  OAI21_X1  g0200(.A(G20), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n240), .A2(G159), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n391), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n259), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n244), .B1(new_n393), .B2(new_n394), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(new_n403), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n405), .B1(new_n407), .B2(KEYINPUT16), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n390), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n377), .A2(new_n378), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n380), .B1(new_n410), .B2(new_n369), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n411), .A2(new_n385), .A3(new_n278), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT77), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(new_n347), .A4(new_n366), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n387), .A2(new_n409), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT17), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n404), .A2(new_n408), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n418), .A2(new_n414), .A3(new_n389), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(KEYINPUT17), .A3(new_n387), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  AOI211_X1 g0222(.A(G179), .B(new_n365), .C1(new_n383), .C2(new_n385), .ZN(new_n423));
  AOI21_X1  g0223(.A(G169), .B1(new_n412), .B2(new_n366), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT76), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n412), .A2(new_n295), .A3(new_n366), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT76), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n426), .B(new_n427), .C1(G169), .C2(new_n386), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n409), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n422), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI211_X1 g0231(.A(KEYINPUT18), .B(new_n409), .C1(new_n425), .C2(new_n428), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n421), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n363), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n338), .A2(new_n340), .A3(G244), .A4(new_n284), .ZN(new_n436));
  XOR2_X1   g0236(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G250), .A2(G1698), .ZN(new_n439));
  NAND2_X1  g0239(.A1(KEYINPUT4), .A2(G244), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(new_n440), .B2(G1698), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n283), .A2(new_n441), .B1(G33), .B2(G283), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT80), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n438), .A2(new_n442), .A3(KEYINPUT80), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n274), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G45), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G1), .ZN(new_n449));
  XNOR2_X1  g0249(.A(KEYINPUT5), .B(G41), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n278), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G257), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n274), .A2(G274), .A3(new_n449), .A4(new_n450), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(G200), .B1(new_n447), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n263), .A2(new_n312), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT78), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n261), .A2(G33), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n268), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n459), .B2(new_n312), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n395), .A2(G107), .A3(new_n397), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n336), .A2(KEYINPUT6), .A3(G97), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n312), .A2(new_n336), .ZN(new_n463));
  NOR2_X1   g0263(.A1(G97), .A2(G107), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n462), .B1(new_n465), .B2(KEYINPUT6), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n466), .A2(G20), .B1(G77), .B2(new_n240), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n460), .B1(new_n468), .B2(new_n259), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n438), .A2(new_n442), .A3(KEYINPUT80), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT80), .B1(new_n438), .B2(new_n442), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n278), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n454), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(G190), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n455), .A2(new_n469), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT81), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n455), .A2(new_n469), .A3(KEYINPUT81), .A4(new_n474), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n452), .A2(new_n295), .A3(new_n453), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT82), .B1(new_n447), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n479), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT82), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n472), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n472), .A2(new_n473), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n468), .A2(new_n259), .ZN(new_n486));
  INV_X1    g0286(.A(new_n460), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n349), .A2(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n477), .A2(new_n478), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n338), .A2(new_n340), .A3(G257), .A4(new_n284), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT85), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT85), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n283), .A2(new_n492), .A3(G257), .A4(new_n284), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n341), .A2(G303), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n283), .A2(G264), .A3(G1698), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n491), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n278), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n450), .A2(new_n449), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(G270), .A3(new_n274), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n453), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n405), .A2(G116), .A3(new_n262), .A4(new_n458), .ZN(new_n503));
  INV_X1    g0303(.A(G116), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n263), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(G20), .B1(G33), .B2(G283), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n255), .A2(G97), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n506), .A2(new_n507), .B1(G20), .B2(new_n504), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n259), .A2(KEYINPUT20), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT20), .B1(new_n259), .B2(new_n508), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n503), .B(new_n505), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n502), .A2(new_n511), .A3(G169), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n512), .B(KEYINPUT21), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT86), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n500), .B1(new_n278), .B2(new_n496), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G179), .ZN(new_n516));
  INV_X1    g0316(.A(new_n511), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n515), .A2(new_n511), .A3(KEYINPUT86), .A4(G179), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n511), .B1(new_n502), .B2(G200), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n347), .B2(new_n502), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n513), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n338), .A2(new_n340), .A3(new_n252), .A4(G87), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT22), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT22), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n283), .A2(new_n526), .A3(new_n252), .A4(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G116), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(G20), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT23), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n252), .B2(G107), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n336), .A2(KEYINPUT23), .A3(G20), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  XOR2_X1   g0334(.A(KEYINPUT87), .B(KEYINPUT24), .Z(new_n535));
  AND3_X1   g0335(.A1(new_n528), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n535), .B1(new_n528), .B2(new_n534), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n259), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n263), .A2(new_n336), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n539), .B(KEYINPUT25), .ZN(new_n540));
  INV_X1    g0340(.A(new_n459), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n283), .A2(G250), .A3(new_n284), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n283), .A2(G257), .A3(G1698), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G294), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n278), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n451), .A2(G264), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n547), .A2(new_n347), .A3(new_n453), .A4(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n453), .A3(new_n548), .ZN(new_n550));
  AOI22_X1  g0350(.A1(KEYINPUT88), .A2(new_n549), .B1(new_n550), .B2(new_n292), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n550), .A2(KEYINPUT88), .A3(new_n292), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n538), .B(new_n542), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n550), .A2(G179), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n546), .A2(new_n278), .B1(G264), .B2(new_n451), .ZN(new_n556));
  AOI21_X1  g0356(.A(G169), .B1(new_n556), .B2(new_n453), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n538), .A2(new_n542), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT84), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n338), .A2(new_n340), .A3(new_n252), .A4(G68), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT19), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n253), .B2(new_n312), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g0366(.A(KEYINPUT83), .B(G87), .ZN(new_n567));
  NAND3_X1  g0367(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n567), .A2(new_n464), .B1(new_n252), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n562), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(G87), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT83), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT83), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G87), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n574), .A3(new_n464), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n568), .A2(new_n252), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n577), .A2(KEYINPUT84), .A3(new_n563), .A4(new_n565), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n570), .A2(new_n259), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n328), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n268), .A2(new_n580), .A3(new_n458), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n328), .A2(new_n263), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n338), .A2(new_n340), .A3(G244), .A4(G1698), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n338), .A2(new_n340), .A3(G238), .A4(new_n284), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n585), .A3(new_n529), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n278), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n278), .A2(new_n279), .ZN(new_n588));
  INV_X1    g0388(.A(G250), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n449), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n588), .A2(new_n449), .B1(new_n274), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n587), .A2(new_n591), .A3(new_n295), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n587), .A2(new_n591), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n593), .B2(G169), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n587), .A2(new_n591), .A3(new_n347), .ZN(new_n595));
  AOI21_X1  g0395(.A(G200), .B1(new_n587), .B2(new_n591), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n268), .A2(G87), .A3(new_n458), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n579), .A2(new_n582), .A3(new_n598), .ZN(new_n599));
  OAI22_X1  g0399(.A1(new_n583), .A2(new_n594), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n554), .A2(new_n561), .A3(new_n600), .ZN(new_n601));
  AND4_X1   g0401(.A1(new_n435), .A2(new_n489), .A3(new_n523), .A4(new_n601), .ZN(G372));
  NOR2_X1   g0402(.A1(new_n431), .A2(new_n432), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n352), .A2(KEYINPUT91), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT91), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n350), .A2(new_n605), .A3(new_n351), .A4(new_n334), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n357), .B2(new_n356), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n608), .A2(new_n326), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n603), .B1(new_n609), .B2(new_n421), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n294), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n298), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n583), .A2(new_n594), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT26), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n485), .A2(new_n349), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n486), .A2(new_n487), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n447), .A2(KEYINPUT82), .A3(new_n479), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n482), .B1(new_n472), .B2(new_n481), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n615), .B1(new_n620), .B2(new_n600), .ZN(new_n621));
  INV_X1    g0421(.A(new_n597), .ZN(new_n622));
  INV_X1    g0422(.A(new_n599), .ZN(new_n623));
  AOI21_X1  g0423(.A(G169), .B1(new_n587), .B2(new_n591), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n295), .B2(new_n593), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n622), .A2(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n627), .A2(new_n488), .A3(KEYINPUT26), .A4(new_n484), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n614), .B1(new_n621), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n477), .A2(new_n478), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n553), .A2(new_n620), .A3(new_n627), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT89), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n477), .A2(new_n478), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n600), .B1(new_n484), .B2(new_n488), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT89), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .A4(new_n553), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT21), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n512), .A2(new_n638), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n512), .A2(new_n638), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n520), .A2(new_n560), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n633), .A2(new_n637), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT90), .ZN(new_n643));
  INV_X1    g0443(.A(new_n641), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n634), .A2(new_n553), .A3(new_n635), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(KEYINPUT89), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT90), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(new_n637), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n630), .B1(new_n643), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n613), .B1(new_n434), .B2(new_n649), .ZN(G369));
  NAND2_X1  g0450(.A1(new_n513), .A2(new_n520), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n261), .A2(new_n252), .A3(G13), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(G213), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n511), .A2(new_n657), .ZN(new_n658));
  MUX2_X1   g0458(.A(new_n651), .B(new_n523), .S(new_n658), .Z(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n560), .A2(new_n657), .ZN(new_n661));
  INV_X1    g0461(.A(new_n559), .ZN(new_n662));
  INV_X1    g0462(.A(new_n657), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n553), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n661), .B1(new_n664), .B2(new_n560), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n651), .A2(new_n663), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n661), .B1(new_n668), .B2(new_n665), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(G399));
  INV_X1    g0470(.A(new_n218), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n575), .A2(G116), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G1), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n215), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n649), .A2(KEYINPUT29), .A3(new_n657), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n620), .A2(new_n615), .A3(new_n600), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n614), .B1(new_n680), .B2(KEYINPUT94), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n634), .A2(new_n641), .A3(new_n635), .A4(new_n553), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT94), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n621), .A2(new_n683), .A3(new_n628), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n679), .B1(new_n685), .B2(new_n663), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n678), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n472), .A2(new_n473), .A3(new_n556), .A4(new_n593), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n689), .B2(new_n516), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n593), .A2(G179), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n485), .A2(new_n691), .A3(new_n502), .A4(new_n550), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT92), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n447), .A2(new_n454), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n502), .A2(new_n295), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n593), .A2(new_n556), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n696), .A2(new_n697), .A3(KEYINPUT30), .A4(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n693), .B2(new_n694), .ZN(new_n700));
  OAI211_X1 g0500(.A(KEYINPUT31), .B(new_n657), .C1(new_n695), .C2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n690), .A3(new_n692), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT93), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n699), .A2(new_n690), .A3(KEYINPUT93), .A4(new_n692), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n657), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n601), .A2(new_n489), .A3(new_n523), .A4(new_n663), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n701), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n687), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n677), .B1(new_n713), .B2(G1), .ZN(G364));
  AND2_X1   g0514(.A1(new_n252), .A2(G13), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n261), .B1(new_n715), .B2(G45), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n672), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n660), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(G330), .B2(new_n659), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G13), .A2(G33), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n211), .B1(G20), .B2(new_n349), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n725), .B(KEYINPUT96), .Z(new_n726));
  NAND2_X1  g0526(.A1(new_n283), .A2(new_n218), .ZN(new_n727));
  INV_X1    g0527(.A(G355), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n727), .A2(new_n728), .B1(G116), .B2(new_n218), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n235), .A2(G45), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n671), .A2(new_n283), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n215), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n732), .B1(new_n448), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n729), .B1(new_n730), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n726), .B1(new_n735), .B2(KEYINPUT95), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(KEYINPUT95), .B2(new_n735), .ZN(new_n737));
  INV_X1    g0537(.A(new_n718), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n252), .A2(G179), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(new_n347), .A3(G200), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n336), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n252), .A2(new_n295), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G190), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n742), .A2(G190), .A3(new_n292), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n283), .B1(new_n744), .B2(new_n286), .C1(new_n243), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n742), .A2(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n347), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n741), .B(new_n746), .C1(G50), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n739), .A2(new_n743), .ZN(new_n750));
  INV_X1    g0550(.A(G159), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g0552(.A(KEYINPUT97), .B(KEYINPUT32), .Z(new_n753));
  XNOR2_X1  g0553(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n347), .A2(G179), .A3(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n252), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n747), .A2(G190), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G97), .A2(new_n757), .B1(new_n758), .B2(G68), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n749), .A2(new_n754), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n739), .A2(G190), .A3(G200), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n761), .A2(KEYINPUT98), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(KEYINPUT98), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n567), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT99), .ZN(new_n767));
  INV_X1    g0567(.A(G311), .ZN(new_n768));
  INV_X1    g0568(.A(G329), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n744), .A2(new_n768), .B1(new_n750), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n745), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n283), .B(new_n770), .C1(G322), .C2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n764), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G303), .ZN(new_n774));
  INV_X1    g0574(.A(new_n740), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n748), .A2(G326), .B1(new_n775), .B2(G283), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G294), .A2(new_n757), .B1(new_n758), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n772), .A2(new_n774), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n766), .B1(new_n767), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n767), .B2(new_n779), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n738), .B1(new_n781), .B2(new_n724), .ZN(new_n782));
  INV_X1    g0582(.A(new_n723), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n737), .B(new_n782), .C1(new_n659), .C2(new_n783), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n720), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G396));
  AOI21_X1  g0586(.A(new_n663), .B1(new_n332), .B2(new_n333), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n348), .A2(new_n352), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n604), .A2(new_n606), .A3(new_n787), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(new_n649), .B2(new_n657), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n642), .A2(KEYINPUT90), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n647), .B1(new_n646), .B2(new_n637), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n629), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n353), .A2(new_n657), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n738), .B1(new_n799), .B2(new_n711), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT101), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n799), .A2(new_n711), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n724), .A2(new_n721), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n718), .B1(G77), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G294), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n745), .A2(new_n808), .B1(new_n750), .B2(new_n768), .ZN(new_n809));
  INV_X1    g0609(.A(new_n744), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n283), .B(new_n809), .C1(G116), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n773), .A2(G107), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G97), .A2(new_n757), .B1(new_n748), .B2(G303), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n740), .A2(new_n571), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G283), .B2(new_n758), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n811), .A2(new_n812), .A3(new_n813), .A4(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G132), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n283), .B1(new_n750), .B2(new_n817), .C1(new_n244), .C2(new_n740), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G58), .B2(new_n757), .ZN(new_n819));
  XNOR2_X1  g0619(.A(KEYINPUT100), .B(G143), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n771), .A2(new_n821), .B1(new_n810), .B2(G159), .ZN(new_n822));
  INV_X1    g0622(.A(new_n748), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  INV_X1    g0624(.A(G150), .ZN(new_n825));
  INV_X1    g0625(.A(new_n758), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n822), .B1(new_n823), .B2(new_n824), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT34), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n819), .B1(new_n242), .B2(new_n764), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n827), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(KEYINPUT34), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n816), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n807), .B1(new_n832), .B2(new_n724), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n791), .B2(new_n722), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n805), .A2(new_n834), .ZN(G384));
  AND2_X1   g0635(.A1(new_n466), .A2(KEYINPUT35), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n466), .A2(KEYINPUT35), .ZN(new_n837));
  NOR4_X1   g0637(.A1(new_n836), .A2(new_n837), .A3(new_n504), .A4(new_n214), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT36), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n733), .B(G77), .C1(new_n243), .C2(new_n244), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n242), .A2(G68), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n261), .B(G13), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT38), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT102), .ZN(new_n845));
  INV_X1    g0645(.A(new_n403), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n393), .A2(new_n394), .ZN(new_n847));
  OAI211_X1 g0647(.A(KEYINPUT16), .B(new_n846), .C1(new_n847), .C2(new_n244), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n391), .B1(new_n406), .B2(new_n403), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n849), .A3(new_n259), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n845), .B1(new_n850), .B2(new_n389), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n655), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n850), .A2(new_n845), .A3(new_n389), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AND4_X1   g0655(.A1(KEYINPUT17), .A2(new_n387), .A3(new_n409), .A4(new_n414), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT17), .B1(new_n419), .B2(new_n387), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n855), .B1(new_n603), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n850), .A2(new_n845), .A3(new_n389), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n861), .A2(new_n851), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n853), .A2(new_n862), .B1(new_n419), .B2(new_n387), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n429), .A2(new_n862), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n430), .A2(new_n853), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n415), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n409), .B1(new_n425), .B2(new_n428), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n867), .A2(new_n868), .A3(KEYINPUT37), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n844), .B1(new_n859), .B2(new_n870), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n861), .B(new_n851), .C1(new_n425), .C2(new_n428), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n855), .A2(new_n415), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT37), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n428), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n366), .B1(new_n376), .B2(new_n381), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n349), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n427), .B1(new_n877), .B2(new_n426), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n430), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n879), .A2(new_n860), .A3(new_n415), .A4(new_n866), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n881), .B(KEYINPUT38), .C1(new_n433), .C2(new_n855), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n871), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n704), .A2(KEYINPUT31), .A3(new_n657), .A4(new_n705), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n708), .A2(new_n709), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n323), .A2(new_n324), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n358), .B2(new_n361), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n360), .A2(new_n663), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n888), .B1(new_n356), .B2(new_n357), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n325), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n792), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n883), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT40), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n893), .A2(new_n896), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT103), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n866), .B1(new_n603), .B2(new_n858), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT37), .B1(new_n867), .B2(new_n868), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n880), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n899), .B(new_n844), .C1(new_n900), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n882), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n880), .A2(new_n901), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n433), .B2(new_n866), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n899), .B1(new_n906), .B2(new_n844), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n898), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n897), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n435), .A2(new_n885), .ZN(new_n910));
  OAI21_X1  g0710(.A(G330), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT104), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n909), .A2(new_n910), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n889), .A2(new_n891), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n352), .A2(new_n657), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n918), .B1(new_n798), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n883), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n904), .B2(new_n907), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n871), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n326), .A2(new_n663), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n924), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n603), .A2(new_n853), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n922), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n678), .A2(new_n686), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n612), .B1(new_n933), .B2(new_n435), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n932), .B(new_n934), .Z(new_n935));
  NAND2_X1  g0735(.A1(new_n916), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n261), .B2(new_n715), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n916), .A2(new_n935), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n843), .B1(new_n937), .B2(new_n938), .ZN(G367));
  OAI21_X1  g0739(.A(new_n489), .B1(new_n469), .B2(new_n663), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n620), .B2(new_n663), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n660), .A2(new_n665), .A3(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(KEYINPUT105), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n599), .A2(new_n657), .ZN(new_n944));
  MUX2_X1   g0744(.A(new_n614), .B(new_n627), .S(new_n944), .Z(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n942), .A2(KEYINPUT105), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n943), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n941), .A2(new_n665), .A3(new_n668), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n620), .B1(new_n940), .B2(new_n560), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n951), .A2(KEYINPUT42), .B1(new_n663), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(KEYINPUT42), .B2(new_n951), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n947), .B1(new_n943), .B2(new_n948), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n950), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n956), .B1(new_n950), .B2(new_n957), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n941), .A2(new_n669), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT45), .Z(new_n962));
  NOR2_X1   g0762(.A1(new_n941), .A2(new_n669), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT44), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(new_n660), .A3(new_n665), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n962), .A2(new_n666), .A3(new_n964), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n668), .B(new_n665), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n660), .B(new_n969), .Z(new_n970));
  OAI21_X1  g0770(.A(new_n713), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n672), .B(KEYINPUT41), .Z(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n960), .B1(new_n974), .B2(new_n716), .ZN(new_n975));
  INV_X1    g0775(.A(new_n750), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n341), .B1(new_n976), .B2(G137), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n977), .B1(new_n242), .B2(new_n744), .C1(new_n825), .C2(new_n745), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n823), .A2(new_n820), .B1(new_n286), .B2(new_n740), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n826), .A2(new_n751), .B1(new_n244), .B2(new_n756), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n243), .B2(new_n764), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT106), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT46), .B1(new_n773), .B2(G116), .ZN(new_n984));
  AOI22_X1  g0784(.A1(G107), .A2(new_n757), .B1(new_n748), .B2(G311), .ZN(new_n985));
  INV_X1    g0785(.A(G303), .ZN(new_n986));
  INV_X1    g0786(.A(G283), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n745), .A2(new_n986), .B1(new_n744), .B2(new_n987), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n283), .B(new_n988), .C1(G317), .C2(new_n976), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n773), .A2(KEYINPUT46), .A3(G116), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n758), .A2(G294), .B1(new_n775), .B2(G97), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n985), .A2(new_n989), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n983), .B1(new_n984), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT47), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n724), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n230), .A2(new_n731), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n724), .B(new_n723), .C1(new_n671), .C2(new_n580), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n738), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n995), .B(new_n998), .C1(new_n783), .C2(new_n945), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT107), .Z(new_n1000));
  NOR2_X1   g0800(.A1(new_n975), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(G387));
  AOI22_X1  g0802(.A1(new_n771), .A2(G317), .B1(new_n810), .B2(G303), .ZN(new_n1003));
  INV_X1    g0803(.A(G322), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1003), .B1(new_n823), .B2(new_n1004), .C1(new_n768), .C2(new_n826), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT48), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n773), .A2(G294), .B1(G283), .B2(new_n757), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT49), .Z(new_n1011));
  AOI21_X1  g0811(.A(new_n283), .B1(new_n976), .B2(G326), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n504), .B2(new_n740), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n251), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n758), .A2(new_n1015), .B1(new_n810), .B2(G68), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT110), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n764), .A2(new_n286), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n283), .B1(new_n750), .B2(new_n825), .C1(new_n745), .C2(new_n242), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n757), .A2(new_n580), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n312), .B2(new_n740), .C1(new_n823), .C2(new_n751), .ZN(new_n1021));
  NOR4_X1   g0821(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n724), .B1(new_n1014), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n227), .A2(G45), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT108), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n330), .A2(G50), .ZN(new_n1026));
  XOR2_X1   g0826(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1027));
  XNOR2_X1  g0827(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n674), .B(new_n448), .C1(new_n244), .C2(new_n286), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1025), .B(new_n731), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(G107), .B2(new_n218), .C1(new_n674), .C2(new_n727), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n726), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n738), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1023), .B(new_n1033), .C1(new_n665), .C2(new_n783), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT111), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n712), .A2(new_n970), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n672), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n970), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n713), .A2(new_n1039), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1035), .B1(new_n716), .B2(new_n970), .C1(new_n1038), .C2(new_n1040), .ZN(G393));
  AOI21_X1  g0841(.A(KEYINPUT114), .B1(new_n1037), .B2(new_n968), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n968), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT114), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1043), .A2(new_n1036), .A3(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n672), .B1(new_n1037), .B2(new_n968), .C1(new_n1042), .C2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n941), .A2(new_n783), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G317), .A2(new_n748), .B1(new_n771), .B2(G311), .ZN(new_n1048));
  XOR2_X1   g0848(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n1049));
  XNOR2_X1  g0849(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n764), .A2(new_n987), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n341), .B1(new_n750), .B2(new_n1004), .C1(new_n744), .C2(new_n808), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n741), .B1(G116), .B2(new_n757), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n986), .B2(new_n826), .ZN(new_n1054));
  NOR4_X1   g0854(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1056), .A2(KEYINPUT113), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n823), .A2(new_n825), .B1(new_n751), .B2(new_n745), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT51), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n756), .A2(new_n286), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n814), .B(new_n1060), .C1(G50), .C2(new_n758), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n773), .A2(G68), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n283), .B1(new_n744), .B2(new_n330), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n976), .B2(new_n821), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .A4(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT113), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n1055), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n724), .B1(new_n1057), .B2(new_n1067), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n725), .B1(new_n312), .B2(new_n218), .C1(new_n238), .C2(new_n732), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n718), .A3(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1047), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n1043), .B2(new_n717), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1046), .A2(new_n1072), .ZN(G390));
  AND2_X1   g0873(.A1(new_n885), .A2(G330), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n435), .A2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1075), .B(new_n613), .C1(new_n687), .C2(new_n434), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n892), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n711), .A2(new_n792), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(new_n917), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n797), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n920), .B1(new_n649), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n685), .A2(new_n663), .A3(new_n791), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n920), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1078), .B2(new_n917), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1074), .A2(new_n791), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n918), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1079), .A2(new_n1081), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1076), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n928), .B1(new_n1083), .B2(new_n917), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n904), .B2(new_n907), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1078), .A2(new_n917), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n879), .A2(KEYINPUT18), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n868), .A2(new_n422), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n858), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n866), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1094), .A2(new_n1095), .B1(new_n880), .B2(new_n901), .ZN(new_n1096));
  OAI21_X1  g0896(.A(KEYINPUT103), .B1(new_n1096), .B2(KEYINPUT38), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(new_n882), .A3(new_n903), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n925), .B1(new_n1098), .B2(new_n923), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n928), .B1(new_n1081), .B2(new_n917), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1090), .B(new_n1091), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1090), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n924), .A2(new_n926), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n919), .B1(new_n796), .B2(new_n797), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n927), .B1(new_n1104), .B2(new_n918), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1102), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1088), .B(new_n1101), .C1(new_n1106), .C2(new_n1077), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1076), .A2(new_n1087), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1101), .B1(new_n1106), .B2(new_n1077), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1110), .A3(new_n672), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1101), .B(new_n717), .C1(new_n1106), .C2(new_n1077), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n718), .B1(new_n1015), .B2(new_n806), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n748), .A2(G283), .B1(new_n810), .B2(G97), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n336), .B2(new_n826), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT116), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n740), .A2(new_n244), .B1(new_n750), .B2(new_n808), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT117), .Z(new_n1118));
  OAI21_X1  g0918(.A(new_n341), .B1(new_n745), .B2(new_n504), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1060), .B(new_n1119), .C1(new_n773), .C2(G87), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1116), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n764), .A2(new_n825), .ZN(new_n1122));
  XOR2_X1   g0922(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1123));
  XNOR2_X1  g0923(.A(new_n1122), .B(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G128), .A2(new_n748), .B1(new_n758), .B2(G137), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n341), .B1(new_n771), .B2(G132), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n810), .A2(new_n1128), .B1(new_n976), .B2(G125), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n757), .A2(G159), .B1(new_n775), .B2(G50), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1125), .A2(new_n1126), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1121), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1113), .B1(new_n1132), .B2(new_n724), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n1099), .B2(new_n722), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1112), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1111), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1136), .A2(KEYINPUT118), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT118), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n1111), .B2(new_n1135), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1137), .A2(new_n1139), .ZN(G378));
  INV_X1    g0940(.A(KEYINPUT120), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n299), .A2(new_n271), .A3(new_n853), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n271), .A2(new_n853), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n294), .A2(new_n298), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1142), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n894), .A2(KEYINPUT40), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT38), .B1(new_n1152), .B2(new_n905), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n855), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1094), .A2(new_n1154), .B1(new_n874), .B2(new_n880), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1153), .A2(new_n899), .B1(KEYINPUT38), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1151), .B1(new_n1156), .B2(new_n1097), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n893), .B1(new_n871), .B2(new_n882), .ZN(new_n1158));
  OAI21_X1  g0958(.A(G330), .B1(new_n1158), .B2(KEYINPUT40), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1150), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n930), .B1(new_n921), .B2(new_n883), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n897), .A2(new_n908), .A3(G330), .A4(new_n1162), .ZN(new_n1163));
  AND4_X1   g0963(.A1(new_n929), .A2(new_n1160), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1163), .A2(new_n1160), .B1(new_n1161), .B2(new_n929), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1141), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n932), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .A4(new_n929), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(KEYINPUT120), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1166), .A2(new_n717), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1150), .A2(new_n721), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n718), .B1(G50), .B2(new_n806), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n740), .A2(new_n243), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n826), .A2(new_n312), .B1(new_n823), .B2(new_n504), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(G68), .C2(new_n757), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1018), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n341), .A2(new_n273), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G283), .B2(new_n976), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n771), .A2(G107), .B1(new_n810), .B2(new_n580), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(KEYINPUT58), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1178), .B(new_n242), .C1(G33), .C2(G41), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT119), .Z(new_n1185));
  AND2_X1   g0985(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(G128), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n745), .A2(new_n1187), .B1(new_n744), .B2(new_n824), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G132), .B2(new_n758), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G150), .A2(new_n757), .B1(new_n748), .B2(G125), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n764), .C2(new_n1127), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n775), .A2(G159), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G33), .B(G41), .C1(new_n976), .C2(G124), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1186), .B1(KEYINPUT58), .B2(new_n1182), .C1(new_n1192), .C2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1173), .B1(new_n1197), .B2(new_n724), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1172), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1171), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1076), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n1109), .B2(new_n1087), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT57), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n672), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1166), .A2(new_n1202), .A3(new_n1170), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n1203), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1206), .B1(new_n1208), .B2(KEYINPUT121), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT121), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1207), .A2(new_n1210), .A3(new_n1203), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1200), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(G375));
  NOR2_X1   g1013(.A1(new_n1087), .A2(new_n716), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n918), .A2(new_n721), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n718), .B1(G68), .B2(new_n806), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n826), .A2(new_n504), .B1(new_n744), .B2(new_n336), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(KEYINPUT122), .A2(new_n1217), .B1(new_n773), .B2(G97), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(KEYINPUT122), .B2(new_n1217), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1020), .B1(new_n286), .B2(new_n740), .C1(new_n823), .C2(new_n808), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n341), .B1(new_n750), .B2(new_n986), .C1(new_n745), .C2(new_n987), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1174), .B1(G50), .B2(new_n757), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n341), .B1(new_n771), .B2(G137), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G150), .A2(new_n810), .B1(new_n976), .B2(G128), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n758), .A2(new_n1128), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n748), .A2(G132), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT123), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n751), .B2(new_n764), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n1219), .A2(new_n1222), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1216), .B1(new_n1231), .B2(new_n724), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1214), .B1(new_n1215), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1088), .A2(new_n972), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1076), .A2(new_n1087), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1234), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(G381));
  OR3_X1    g1038(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1239), .A2(G390), .A3(G381), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1136), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1240), .A2(new_n1212), .A3(new_n1001), .A4(new_n1241), .ZN(G407));
  INV_X1    g1042(.A(G213), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(G343), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1212), .A2(new_n1241), .A3(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(G407), .A2(G213), .A3(new_n1245), .ZN(G409));
  NAND3_X1  g1046(.A1(G387), .A2(new_n1046), .A3(new_n1072), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(G393), .B(new_n785), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(G390), .A2(new_n1001), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1248), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT60), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1236), .B1(new_n1088), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1076), .A2(KEYINPUT60), .A3(new_n1087), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n672), .A3(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(G384), .A3(new_n1233), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(G384), .B1(new_n1257), .B2(new_n1233), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1244), .ZN(new_n1262));
  INV_X1    g1062(.A(G2897), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1261), .A2(KEYINPUT125), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1257), .A2(new_n1233), .ZN(new_n1266));
  INV_X1    g1066(.A(G384), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1258), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT125), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1268), .A2(KEYINPUT125), .A3(new_n1258), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1264), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1265), .B1(new_n1272), .B2(new_n1275), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1207), .A2(new_n972), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1278), .A2(KEYINPUT124), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n716), .B1(new_n1278), .B2(KEYINPUT124), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1279), .A2(new_n1280), .B1(new_n1172), .B2(new_n1198), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1136), .B1(new_n1277), .B2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(new_n1212), .B2(G378), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1276), .B1(new_n1283), .B2(new_n1244), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1208), .A2(KEYINPUT121), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1206), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(new_n1211), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1200), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(G378), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1282), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n1244), .B(new_n1269), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1284), .B(new_n1285), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1244), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1261), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1296), .A2(KEYINPUT62), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1253), .B1(new_n1294), .B2(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1264), .B1(new_n1261), .B2(KEYINPUT125), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1299), .B1(new_n1300), .B2(new_n1271), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1285), .B(new_n1252), .C1(new_n1295), .C2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1296), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1306), .A2(KEYINPUT63), .A3(new_n1262), .A4(new_n1261), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(KEYINPUT126), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT126), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1292), .A2(new_n1309), .A3(KEYINPUT63), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1303), .A2(new_n1305), .A3(new_n1308), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1298), .A2(new_n1311), .ZN(G405));
  NAND2_X1  g1112(.A1(G375), .A2(new_n1241), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1290), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT127), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1261), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1269), .A2(KEYINPUT127), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1314), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1313), .A2(new_n1315), .A3(new_n1290), .A4(new_n1261), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1318), .A2(new_n1319), .A3(new_n1252), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1252), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(G402));
endmodule


