//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1210, new_n1211, new_n1212, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  XOR2_X1   g0009(.A(KEYINPUT66), .B(G244), .Z(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  OR3_X1    g0019(.A1(new_n209), .A2(KEYINPUT64), .A3(G13), .ZN(new_n220));
  OAI21_X1  g0020(.A(KEYINPUT64), .B1(new_n209), .B2(G13), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT0), .Z(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT65), .Z(new_n230));
  AOI211_X1 g0030(.A(new_n219), .B(new_n224), .C1(new_n227), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n225), .ZN(new_n248));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G13), .A3(G20), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n249), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n226), .A2(G1), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(G50), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n252), .A2(new_n253), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n226), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n259), .A2(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(G20), .B2(new_n203), .ZN(new_n265));
  INV_X1    g0065(.A(new_n248), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n257), .B1(G50), .B2(new_n258), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT9), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  INV_X1    g0069(.A(new_n225), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n271), .A2(G1), .A3(G13), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G226), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OR2_X1    g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1698), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n284), .A2(G222), .B1(new_n287), .B2(G77), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n282), .A2(new_n283), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G1698), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT67), .B(G223), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n281), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n267), .A2(new_n268), .B1(G190), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G200), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n295), .B1(new_n268), .B2(new_n267), .C1(new_n296), .C2(new_n294), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT10), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT15), .B(G87), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT70), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(new_n260), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n259), .A2(new_n263), .B1(new_n226), .B2(new_n211), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n248), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OR3_X1    g0104(.A1(new_n258), .A2(KEYINPUT71), .A3(G77), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT71), .B1(new_n258), .B2(G77), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n255), .A2(new_n211), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n305), .A2(new_n306), .B1(new_n254), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n284), .A2(G232), .B1(new_n287), .B2(G107), .ZN(new_n310));
  INV_X1    g0110(.A(G238), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(new_n290), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n293), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n293), .A2(new_n269), .A3(new_n278), .ZN(new_n314));
  INV_X1    g0114(.A(new_n210), .ZN(new_n315));
  INV_X1    g0115(.A(new_n279), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n309), .B1(G200), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT72), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n320), .ZN(new_n322));
  INV_X1    g0122(.A(new_n318), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G190), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n298), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n316), .A2(KEYINPUT78), .A3(G232), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT78), .ZN(new_n328));
  INV_X1    g0128(.A(G232), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n328), .B1(new_n279), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n280), .A2(G1698), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(G223), .B2(G1698), .ZN(new_n333));
  INV_X1    g0133(.A(G33), .ZN(new_n334));
  INV_X1    g0134(.A(G87), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n333), .A2(new_n287), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n314), .B1(new_n336), .B2(new_n293), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT79), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT79), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n331), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(G169), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n338), .A2(G179), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G58), .ZN(new_n345));
  INV_X1    g0145(.A(G68), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n347), .A2(new_n201), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(G20), .B1(G159), .B2(new_n262), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n289), .A2(new_n350), .A3(G20), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT75), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n289), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n287), .A2(KEYINPUT75), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(new_n354), .A3(new_n226), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n351), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(KEYINPUT16), .B(new_n349), .C1(new_n357), .C2(new_n346), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT16), .ZN(new_n359));
  INV_X1    g0159(.A(new_n349), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n350), .B1(new_n289), .B2(G20), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n287), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n346), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n359), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n358), .A2(new_n364), .A3(new_n248), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n259), .A2(new_n255), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT77), .ZN(new_n367));
  INV_X1    g0167(.A(new_n258), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n367), .A2(new_n254), .B1(new_n368), .B2(new_n259), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n344), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT18), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT17), .ZN(new_n373));
  INV_X1    g0173(.A(G190), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n374), .A2(KEYINPUT80), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(KEYINPUT80), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n338), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n339), .A2(new_n341), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n378), .B1(new_n379), .B2(new_n296), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n373), .B1(new_n380), .B2(new_n370), .ZN(new_n381));
  INV_X1    g0181(.A(new_n370), .ZN(new_n382));
  INV_X1    g0182(.A(new_n341), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n340), .B1(new_n331), .B2(new_n337), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n385), .A2(G200), .B1(new_n338), .B2(new_n377), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n382), .A2(new_n386), .A3(KEYINPUT17), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT18), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n344), .A2(new_n388), .A3(new_n370), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n372), .A2(new_n381), .A3(new_n387), .A4(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n254), .A2(G68), .A3(new_n256), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n346), .A2(G20), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n393), .B1(new_n260), .B2(new_n211), .C1(new_n263), .C2(new_n202), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n248), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n395), .A2(KEYINPUT11), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(KEYINPUT11), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n392), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n258), .A2(G68), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n399), .B(KEYINPUT12), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n329), .A2(G1698), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n289), .B(new_n403), .C1(G226), .C2(G1698), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G97), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n293), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n276), .B1(new_n279), .B2(new_n311), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT13), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n277), .B1(new_n404), .B2(new_n405), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT13), .B1(new_n412), .B2(new_n408), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G169), .ZN(new_n415));
  INV_X1    g0215(.A(G179), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n415), .A2(KEYINPUT14), .B1(new_n416), .B2(new_n414), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n415), .A2(KEYINPUT14), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n402), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n296), .B1(new_n411), .B2(new_n413), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT73), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n414), .A2(new_n374), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n402), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT74), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n422), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n422), .B2(new_n424), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n419), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n294), .A2(new_n416), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n267), .C1(G169), .C2(new_n294), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n431), .B(KEYINPUT69), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n323), .A2(new_n416), .ZN(new_n433));
  INV_X1    g0233(.A(G169), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n318), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n309), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n326), .A2(new_n391), .A3(new_n429), .A4(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT21), .ZN(new_n441));
  OAI211_X1 g0241(.A(G264), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n442));
  INV_X1    g0242(.A(G1698), .ZN(new_n443));
  OAI211_X1 g0243(.A(G257), .B(new_n443), .C1(new_n285), .C2(new_n286), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n282), .A2(G303), .A3(new_n283), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n446), .A2(new_n293), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT5), .B(G41), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n249), .A2(G45), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(G270), .A3(new_n277), .ZN(new_n452));
  NOR2_X1   g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(KEYINPUT5), .A2(G41), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n449), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n272), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(G169), .B1(new_n447), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n249), .A2(G33), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n258), .A2(G116), .A3(new_n266), .A4(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G116), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n252), .A2(new_n462), .A3(new_n253), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n247), .A2(new_n225), .B1(G20), .B2(new_n462), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n466), .B(new_n226), .C1(G33), .C2(new_n205), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n465), .A2(KEYINPUT20), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT20), .B1(new_n465), .B2(new_n467), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n441), .B1(new_n459), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(G200), .B1(new_n447), .B2(new_n458), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n448), .A2(new_n450), .B1(new_n270), .B2(new_n271), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n474), .A2(G270), .B1(new_n272), .B2(new_n456), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n446), .A2(new_n293), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(new_n377), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n473), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n461), .B(new_n463), .C1(new_n469), .C2(new_n468), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n479), .A2(G179), .A3(new_n476), .A4(new_n475), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n475), .A2(new_n476), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT21), .A4(G169), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n472), .A2(new_n478), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT83), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n482), .A2(new_n480), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT83), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n485), .A2(new_n486), .A3(new_n472), .A4(new_n478), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n289), .A2(G238), .A3(new_n443), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G116), .ZN(new_n490));
  OAI211_X1 g0290(.A(G244), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n293), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n450), .A2(new_n277), .A3(G274), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n277), .A2(G250), .A3(new_n449), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G200), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n289), .A2(new_n226), .A3(G68), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT19), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n226), .B1(new_n405), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(G87), .B2(new_n207), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n501), .B1(new_n260), .B2(new_n205), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n500), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n248), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n301), .A2(new_n368), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n254), .A2(G87), .A3(new_n460), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n496), .B1(new_n492), .B2(new_n293), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G190), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n499), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  XNOR2_X1  g0313(.A(new_n299), .B(KEYINPUT70), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(new_n254), .A3(new_n460), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n506), .A3(new_n507), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT82), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n515), .A2(new_n506), .A3(new_n507), .A4(KEYINPUT82), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n510), .A2(KEYINPUT81), .A3(new_n416), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n510), .A2(new_n416), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT81), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n522), .A2(new_n523), .B1(new_n498), .B2(new_n434), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n513), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(G257), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n526));
  OAI211_X1 g0326(.A(G250), .B(new_n443), .C1(new_n285), .C2(new_n286), .ZN(new_n527));
  INV_X1    g0327(.A(G294), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n527), .C1(new_n334), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n293), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n474), .A2(G264), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n457), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n434), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n529), .A2(new_n293), .B1(G264), .B2(new_n474), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(new_n416), .A3(new_n457), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g0336(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT87), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT23), .B1(new_n226), .B2(G107), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT23), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(new_n206), .A3(G20), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n226), .A2(G33), .A3(G116), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT86), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n540), .A2(new_n542), .A3(new_n543), .A4(KEYINPUT86), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n539), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n226), .B(G87), .C1(new_n285), .C2(new_n286), .ZN(new_n549));
  AND2_X1   g0349(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n537), .A2(new_n538), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n548), .A2(new_n551), .A3(new_n538), .A4(new_n537), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n266), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n254), .A2(new_n460), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n368), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT25), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n258), .B2(G107), .ZN(new_n561));
  AOI22_X1  g0361(.A1(G107), .A2(new_n558), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n536), .B1(new_n556), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n555), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n548), .A2(new_n551), .B1(new_n538), .B2(new_n537), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n248), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n532), .A2(new_n296), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(G190), .B2(new_n532), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n569), .A3(new_n562), .ZN(new_n570));
  OAI211_X1 g0370(.A(G250), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n571));
  OAI211_X1 g0371(.A(G244), .B(new_n443), .C1(new_n285), .C2(new_n286), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT4), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n466), .B(new_n571), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT4), .B1(new_n284), .B2(G244), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n293), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n474), .A2(G257), .B1(new_n272), .B2(new_n456), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n416), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n258), .A2(G97), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n558), .B2(G97), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT6), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n582), .A2(new_n205), .A3(G107), .ZN(new_n583));
  XNOR2_X1  g0383(.A(G97), .B(G107), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n583), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n585), .A2(new_n226), .B1(new_n211), .B2(new_n263), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n206), .B1(new_n361), .B2(new_n362), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n248), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n581), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n576), .A2(new_n577), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n434), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n579), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n578), .A2(G190), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(G200), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n593), .A2(new_n588), .A3(new_n581), .A4(new_n594), .ZN(new_n595));
  AND4_X1   g0395(.A1(new_n564), .A2(new_n570), .A3(new_n592), .A4(new_n595), .ZN(new_n596));
  AND4_X1   g0396(.A1(new_n440), .A2(new_n488), .A3(new_n525), .A4(new_n596), .ZN(G372));
  NAND2_X1  g0397(.A1(new_n387), .A2(new_n381), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n437), .B1(new_n426), .B2(new_n427), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n598), .B1(new_n599), .B2(new_n419), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n372), .A2(new_n389), .ZN(new_n601));
  OR2_X1    g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n432), .B1(new_n602), .B2(new_n298), .ZN(new_n603));
  INV_X1    g0403(.A(new_n592), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n524), .A2(new_n519), .A3(new_n520), .A4(new_n518), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT26), .A4(new_n512), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT26), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n522), .B(new_n516), .C1(G169), .C2(new_n510), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n512), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n607), .B1(new_n609), .B2(new_n592), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n606), .A2(KEYINPUT88), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT88), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n525), .A2(new_n612), .A3(KEYINPUT26), .A4(new_n604), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n512), .A2(new_n608), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n615), .A2(new_n570), .A3(new_n592), .A4(new_n595), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n472), .A2(new_n480), .A3(new_n482), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n567), .A2(new_n562), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n536), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n608), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  OR2_X1    g0420(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n440), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n603), .A2(new_n622), .ZN(G369));
  NAND3_X1  g0423(.A1(new_n249), .A2(new_n226), .A3(G13), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(G213), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(G343), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n479), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n488), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT89), .ZN(new_n632));
  INV_X1    g0432(.A(new_n630), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n617), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n633), .B1(new_n484), .B2(new_n487), .ZN(new_n636));
  INV_X1    g0436(.A(new_n634), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT89), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n618), .A2(new_n629), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(new_n564), .A3(new_n570), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n618), .A2(new_n536), .A3(new_n629), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n640), .A2(G330), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n629), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n617), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n618), .A2(new_n536), .A3(new_n646), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n645), .A2(new_n651), .ZN(G399));
  NAND2_X1  g0452(.A1(new_n222), .A2(new_n273), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT90), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n655), .A2(new_n249), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n229), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(new_n655), .ZN(new_n660));
  XOR2_X1   g0460(.A(new_n660), .B(KEYINPUT28), .Z(new_n661));
  NAND3_X1  g0461(.A1(new_n475), .A2(new_n476), .A3(G179), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n578), .A2(new_n663), .A3(new_n510), .A4(new_n534), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT30), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n510), .A2(new_n534), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n662), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(KEYINPUT30), .A3(new_n578), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(G179), .B1(new_n493), .B2(new_n497), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n671), .A2(new_n590), .A3(new_n481), .A4(new_n532), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT91), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n457), .A2(new_n534), .B1(new_n576), .B2(new_n577), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n675), .A2(KEYINPUT91), .A3(new_n481), .A4(new_n671), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n629), .B1(new_n670), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT31), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT92), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n596), .A2(new_n488), .A3(new_n525), .A4(new_n646), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT92), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n678), .A2(new_n683), .A3(new_n679), .ZN(new_n684));
  INV_X1    g0484(.A(new_n672), .ZN(new_n685));
  OAI211_X1 g0485(.A(KEYINPUT31), .B(new_n629), .C1(new_n670), .C2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n681), .A2(new_n682), .A3(new_n684), .A4(new_n686), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n687), .A2(KEYINPUT93), .A3(G330), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT93), .B1(new_n687), .B2(G330), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n604), .A2(new_n605), .A3(new_n607), .A4(new_n512), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT26), .B1(new_n609), .B2(new_n592), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n646), .B1(new_n620), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT29), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT29), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n695), .B(new_n646), .C1(new_n614), .C2(new_n620), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n688), .A2(new_n689), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n661), .B1(new_n698), .B2(G1), .ZN(G364));
  NAND3_X1  g0499(.A1(new_n635), .A2(G330), .A3(new_n638), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n226), .A2(G13), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n249), .B1(new_n701), .B2(G45), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n655), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT94), .B1(new_n640), .B2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n640), .A2(KEYINPUT94), .A3(G330), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n700), .B(new_n705), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n225), .B1(G20), .B2(new_n434), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n374), .A2(G179), .A3(G200), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n226), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n205), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n226), .A2(G179), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(new_n374), .A3(new_n296), .ZN(new_n716));
  INV_X1    g0516(.A(G159), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT32), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n377), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n226), .A2(new_n416), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G200), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n718), .B1(new_n723), .B2(new_n202), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n720), .A2(new_n296), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  AOI211_X1 g0526(.A(new_n714), .B(new_n724), .C1(G58), .C2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n720), .A2(new_n374), .A3(G200), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT97), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n728), .A2(KEYINPUT97), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n715), .A2(new_n374), .A3(G200), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n734), .B(KEYINPUT96), .Z(new_n735));
  AOI22_X1  g0535(.A1(new_n733), .A2(G68), .B1(G107), .B2(new_n735), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n716), .A2(KEYINPUT32), .A3(new_n717), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n725), .A2(G190), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n737), .B1(G77), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n715), .A2(G190), .A3(G200), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n335), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n287), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT95), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n727), .A2(new_n736), .A3(new_n739), .A4(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n726), .ZN(new_n745));
  INV_X1    g0545(.A(G322), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n745), .A2(new_n746), .B1(new_n528), .B2(new_n713), .ZN(new_n747));
  XOR2_X1   g0547(.A(KEYINPUT98), .B(G326), .Z(new_n748));
  INV_X1    g0548(.A(G311), .ZN(new_n749));
  INV_X1    g0549(.A(new_n738), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n723), .A2(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n716), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n289), .B1(new_n752), .B2(G329), .ZN(new_n753));
  INV_X1    g0553(.A(G303), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n753), .B1(new_n754), .B2(new_n740), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n747), .A2(new_n751), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n735), .A2(G283), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT33), .B(G317), .Z(new_n758));
  OAI211_X1 g0558(.A(new_n756), .B(new_n757), .C1(new_n732), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n711), .B1(new_n744), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n222), .A2(G355), .A3(new_n289), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(G116), .B2(new_n222), .ZN(new_n762));
  INV_X1    g0562(.A(new_n222), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n353), .A2(new_n354), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n274), .B2(new_n230), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n242), .A2(new_n274), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n762), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n710), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n704), .B1(new_n770), .B2(new_n775), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n760), .B(new_n776), .C1(new_n639), .C2(new_n773), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n709), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT99), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n779), .B(new_n780), .ZN(G396));
  NOR2_X1   g0581(.A1(new_n688), .A2(new_n689), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n621), .A2(new_n646), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n309), .A2(new_n629), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n437), .B1(new_n325), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n436), .A2(new_n629), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n621), .A2(new_n787), .A3(new_n646), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n704), .B1(new_n782), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(new_n782), .B2(new_n791), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n711), .A2(new_n772), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n704), .B1(G77), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n726), .A2(G294), .B1(G116), .B2(new_n738), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n797), .B1(new_n206), .B2(new_n740), .C1(new_n754), .C2(new_n723), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n735), .A2(G87), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT100), .B(G283), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n732), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n287), .B1(new_n716), .B2(new_n749), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n798), .A2(new_n801), .A3(new_n714), .A4(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n722), .A2(G137), .B1(G159), .B2(new_n738), .ZN(new_n804));
  INV_X1    g0604(.A(G143), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n804), .B1(new_n805), .B2(new_n745), .C1(new_n732), .C2(new_n261), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT34), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n764), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G132), .B2(new_n752), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n735), .A2(G68), .ZN(new_n811));
  INV_X1    g0611(.A(new_n713), .ZN(new_n812));
  INV_X1    g0612(.A(new_n740), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n812), .A2(G58), .B1(new_n813), .B2(G50), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n810), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(new_n806), .B2(new_n807), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n803), .B1(new_n808), .B2(new_n816), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n796), .B1(new_n711), .B2(new_n817), .C1(new_n787), .C2(new_n772), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n793), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G384));
  OAI21_X1  g0620(.A(new_n349), .B1(new_n357), .B2(new_n346), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n359), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n822), .A2(new_n248), .A3(new_n358), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n627), .B1(new_n823), .B2(new_n369), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n390), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT101), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n434), .B1(new_n383), .B2(new_n384), .ZN(new_n827));
  INV_X1    g0627(.A(new_n343), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n829), .A2(new_n627), .B1(new_n823), .B2(new_n369), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n380), .A2(new_n370), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n826), .B(KEYINPUT37), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n382), .A2(new_n386), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT37), .ZN(new_n834));
  INV_X1    g0634(.A(new_n627), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n370), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n833), .A2(new_n371), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n823), .A2(new_n369), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n627), .B1(new_n342), .B2(new_n343), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n833), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n826), .B1(new_n842), .B2(KEYINPUT37), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n825), .B(KEYINPUT38), .C1(new_n838), .C2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n839), .A2(new_n840), .B1(new_n382), .B2(new_n386), .ZN(new_n846));
  OAI21_X1  g0646(.A(KEYINPUT101), .B1(new_n846), .B2(new_n834), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(new_n837), .A3(new_n832), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT38), .B1(new_n848), .B2(new_n825), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT39), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n390), .A2(new_n370), .A3(new_n835), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n833), .A2(new_n371), .A3(new_n836), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n837), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT38), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT39), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(new_n844), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n850), .A2(KEYINPUT102), .A3(new_n859), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n419), .A2(new_n629), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n825), .B1(new_n838), .B2(new_n843), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n856), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n844), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT102), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT39), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n860), .A2(new_n862), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n401), .A2(new_n646), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n428), .A2(new_n869), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n419), .B1(new_n401), .B2(new_n646), .C1(new_n426), .C2(new_n427), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n786), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n873), .B1(new_n790), .B2(new_n874), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n875), .A2(new_n865), .B1(new_n601), .B2(new_n627), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n868), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n440), .A2(new_n697), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n603), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n877), .B(new_n879), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n678), .A2(new_n679), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n682), .A3(new_n680), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n872), .A2(new_n882), .A3(new_n787), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n857), .A2(new_n844), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT40), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT40), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n883), .A2(new_n865), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(new_n440), .A3(new_n882), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n440), .A2(new_n882), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n886), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n890), .A2(G330), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n880), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n894), .A2(KEYINPUT103), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(KEYINPUT103), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n880), .A2(new_n893), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n701), .A2(new_n249), .ZN(new_n898));
  NOR4_X1   g0698(.A1(new_n895), .A2(new_n896), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n585), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n900), .A2(KEYINPUT35), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(KEYINPUT35), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n901), .A2(G116), .A3(new_n227), .A4(new_n902), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(KEYINPUT36), .Z(new_n904));
  OR3_X1    g0704(.A1(new_n229), .A2(new_n211), .A3(new_n347), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n202), .A2(G68), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n249), .B(G13), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  OR3_X1    g0707(.A1(new_n899), .A2(new_n904), .A3(new_n907), .ZN(G367));
  NAND2_X1  g0708(.A1(new_n604), .A2(new_n629), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n589), .A2(new_n629), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n595), .A2(new_n592), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n648), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n913), .A2(KEYINPUT42), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT104), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n911), .A2(new_n564), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n629), .B1(new_n916), .B2(new_n592), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n913), .B2(KEYINPUT42), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n509), .A2(new_n646), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n615), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n608), .B2(new_n920), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n915), .A2(new_n918), .B1(KEYINPUT43), .B2(new_n922), .ZN(new_n923));
  OR3_X1    g0723(.A1(new_n923), .A2(KEYINPUT43), .A3(new_n922), .ZN(new_n924));
  INV_X1    g0724(.A(new_n912), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n645), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n923), .B1(KEYINPUT43), .B2(new_n922), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n926), .B1(new_n924), .B2(new_n927), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n655), .B(new_n931), .Z(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT109), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT107), .B1(new_n642), .B2(new_n647), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n700), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n644), .B1(new_n617), .B2(new_n646), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n635), .A2(new_n638), .A3(G330), .A4(new_n935), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n938), .B1(new_n937), .B2(new_n939), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT108), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n687), .A2(G330), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT93), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n687), .A2(KEYINPUT93), .A3(G330), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n694), .A2(new_n696), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n942), .A2(new_n943), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n937), .A2(new_n939), .ZN(new_n951));
  INV_X1    g0751(.A(new_n938), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT108), .B1(new_n955), .B2(new_n698), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n934), .B1(new_n950), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n943), .B1(new_n942), .B2(new_n949), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n955), .A2(new_n698), .A3(KEYINPUT108), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n958), .A2(KEYINPUT109), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n651), .A2(new_n912), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT45), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n961), .B(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n925), .B1(new_n648), .B2(new_n650), .ZN(new_n964));
  XNOR2_X1  g0764(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n963), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(new_n645), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n957), .A2(new_n960), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n933), .B1(new_n970), .B2(new_n698), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n930), .B1(new_n971), .B2(new_n703), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n766), .A2(new_n238), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n775), .B1(new_n514), .B2(new_n763), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n705), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n773), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n722), .A2(G143), .B1(G68), .B2(new_n812), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n261), .B2(new_n745), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT110), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(KEYINPUT110), .ZN(new_n980));
  INV_X1    g0780(.A(G137), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n289), .B1(new_n716), .B2(new_n981), .C1(new_n345), .C2(new_n740), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n750), .A2(new_n202), .B1(new_n734), .B2(new_n211), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(new_n733), .C2(G159), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n979), .A2(new_n980), .A3(new_n984), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n745), .A2(new_n754), .B1(new_n206), .B2(new_n713), .ZN(new_n986));
  INV_X1    g0786(.A(new_n800), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n986), .B1(new_n738), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n764), .B1(G317), .B2(new_n752), .ZN(new_n989));
  INV_X1    g0789(.A(new_n734), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n722), .A2(G311), .B1(G97), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT46), .B1(new_n740), .B2(new_n462), .ZN(new_n992));
  OR3_X1    g0792(.A1(new_n740), .A2(KEYINPUT46), .A3(new_n462), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n733), .A2(G294), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n988), .A2(new_n989), .A3(new_n991), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n985), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n975), .B1(new_n976), .B2(new_n922), .C1(new_n998), .C2(new_n711), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n972), .A2(new_n999), .ZN(G387));
  NAND3_X1  g0800(.A1(new_n642), .A2(new_n643), .A3(new_n773), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n765), .B1(new_n235), .B2(new_n274), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n222), .A2(new_n657), .A3(new_n289), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OR3_X1    g0804(.A1(new_n259), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT50), .B1(new_n259), .B2(G50), .ZN(new_n1006));
  AOI21_X1  g0806(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1005), .A2(new_n656), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1004), .A2(new_n1008), .B1(new_n206), .B2(new_n763), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n704), .B1(new_n1009), .B2(new_n775), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n740), .A2(new_n211), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n745), .A2(new_n202), .B1(new_n346), .B2(new_n750), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(G159), .C2(new_n722), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n514), .A2(new_n812), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n809), .B1(G150), .B2(new_n752), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n259), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n733), .A2(new_n1016), .B1(G97), .B2(new_n735), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n748), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n764), .B1(new_n752), .B2(new_n1019), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n713), .A2(new_n800), .B1(new_n740), .B2(new_n528), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT112), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n726), .A2(G317), .B1(G303), .B2(new_n738), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n746), .B2(new_n723), .C1(new_n732), .C2(new_n749), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT48), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n1025), .B2(new_n1024), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT49), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1020), .B1(new_n462), .B2(new_n734), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1018), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1010), .B1(new_n1031), .B2(new_n710), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n955), .A2(new_n703), .B1(new_n1001), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n958), .A2(new_n959), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n655), .B(KEYINPUT113), .Z(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n955), .B2(new_n698), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1033), .B1(new_n1035), .B2(new_n1037), .ZN(G393));
  OAI211_X1 g0838(.A(new_n970), .B(new_n1036), .C1(new_n1035), .C2(new_n969), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n925), .A2(new_n773), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT114), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n774), .B1(new_n205), .B2(new_n222), .C1(new_n766), .C2(new_n245), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n704), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G150), .A2(new_n722), .B1(new_n726), .B2(G159), .ZN(new_n1044));
  XOR2_X1   g0844(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1045));
  XNOR2_X1  g0845(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1046), .B(new_n799), .C1(new_n202), .C2(new_n732), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n764), .B1(new_n805), .B2(new_n716), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G77), .A2(new_n812), .B1(new_n738), .B2(new_n1016), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n346), .B2(new_n740), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(KEYINPUT116), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G311), .A2(new_n726), .B1(new_n722), .B2(G317), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT52), .Z(new_n1055));
  OAI221_X1 g0855(.A(new_n287), .B1(new_n716), .B2(new_n746), .C1(new_n740), .C2(new_n800), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n750), .A2(new_n528), .B1(new_n713), .B2(new_n462), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(G107), .C2(new_n735), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1055), .B(new_n1058), .C1(new_n754), .C2(new_n732), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1052), .A2(KEYINPUT116), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1053), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1043), .B1(new_n1061), .B2(new_n710), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n969), .A2(new_n703), .B1(new_n1041), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1039), .A2(new_n1063), .ZN(G390));
  OR2_X1    g0864(.A1(new_n693), .A2(new_n785), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n874), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n872), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(new_n861), .A3(new_n884), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n788), .B1(new_n946), .B2(new_n947), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n872), .ZN(new_n1070));
  AOI211_X1 g0870(.A(KEYINPUT102), .B(new_n858), .C1(new_n864), .C2(new_n844), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n866), .B1(new_n865), .B2(KEYINPUT39), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1071), .B1(new_n1072), .B2(new_n859), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n790), .A2(new_n874), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n862), .B1(new_n1074), .B2(new_n872), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1068), .B(new_n1070), .C1(new_n1073), .C2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n872), .A2(new_n787), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n882), .A2(G330), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1075), .B1(new_n860), .B2(new_n867), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1068), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1076), .A2(new_n1082), .A3(new_n703), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n704), .B1(new_n1016), .B2(new_n794), .ZN(new_n1084));
  XOR2_X1   g0884(.A(KEYINPUT54), .B(G143), .Z(new_n1085));
  AOI22_X1  g0885(.A1(new_n726), .A2(G132), .B1(new_n738), .B2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n812), .A2(G159), .B1(new_n752), .B2(G125), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n722), .A2(G128), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n289), .B1(new_n734), .B2(new_n202), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT118), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n740), .A2(new_n261), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT53), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1091), .B(new_n1093), .C1(new_n981), .C2(new_n732), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n726), .A2(G116), .B1(G77), .B2(new_n812), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n722), .A2(G283), .B1(G97), .B2(new_n738), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n289), .B(new_n741), .C1(G294), .C2(new_n752), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n811), .B1(new_n732), .B2(new_n206), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n1089), .A2(new_n1094), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1084), .B1(new_n1100), .B2(new_n710), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1073), .B2(new_n772), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1083), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1036), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1076), .A2(new_n1082), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1066), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n882), .A2(KEYINPUT117), .A3(G330), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n787), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT117), .B1(new_n882), .B2(G330), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n873), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1070), .A2(new_n1106), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1074), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n787), .B1(new_n688), .B2(new_n689), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1079), .B1(new_n1113), .B2(new_n873), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1111), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  OR2_X1    g0915(.A1(new_n439), .A2(new_n1078), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n603), .A2(new_n878), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1104), .B1(new_n1105), .B2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1076), .A2(new_n1082), .A3(new_n1115), .A4(new_n1118), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1103), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(G378));
  NAND2_X1  g0923(.A1(new_n267), .A2(new_n835), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n298), .A2(new_n431), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1124), .B1(new_n298), .B2(new_n431), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OR3_X1    g0928(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1128), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n889), .B2(G330), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n887), .B1(new_n883), .B2(new_n884), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n872), .A2(new_n882), .A3(new_n887), .A4(new_n787), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n844), .B2(new_n864), .ZN(new_n1135));
  OAI211_X1 g0935(.A(G330), .B(new_n1131), .C1(new_n1133), .C2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n877), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n868), .A2(new_n876), .ZN(new_n1139));
  OAI21_X1  g0939(.A(G330), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1140), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1139), .A2(new_n1141), .A3(new_n1136), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n703), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n704), .B1(G50), .B2(new_n794), .ZN(new_n1145));
  INV_X1    g0945(.A(G283), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n273), .B1(new_n716), .B2(new_n1146), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1147), .B(new_n764), .C1(new_n514), .C2(new_n738), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1011), .B1(G68), .B2(new_n812), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n734), .A2(new_n345), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n722), .B2(G116), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1148), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n726), .A2(G107), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT120), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(G97), .C2(new_n733), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT58), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n764), .A2(G33), .ZN(new_n1157));
  AOI21_X1  g0957(.A(G50), .B1(new_n1157), .B2(new_n273), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT119), .Z(new_n1159));
  AND2_X1   g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n713), .A2(new_n261), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n726), .A2(G128), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1161), .B(new_n1162), .C1(G125), .C2(new_n722), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n738), .A2(G137), .B1(new_n813), .B2(new_n1085), .ZN(new_n1164));
  INV_X1    g0964(.A(G132), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1163), .B(new_n1164), .C1(new_n1165), .C2(new_n732), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n990), .A2(G159), .ZN(new_n1169));
  AOI211_X1 g0969(.A(G33), .B(G41), .C1(new_n752), .C2(G124), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1160), .B1(KEYINPUT58), .B2(new_n1155), .C1(new_n1167), .C2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1145), .B1(new_n1172), .B2(new_n710), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n1131), .B2(new_n772), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1144), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1121), .A2(new_n1118), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1139), .A2(new_n1141), .A3(KEYINPUT121), .A4(new_n1136), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT121), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1138), .A2(new_n1142), .A3(new_n1178), .ZN(new_n1179));
  AND4_X1   g0979(.A1(KEYINPUT57), .A2(new_n1176), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1121), .A2(new_n1118), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1036), .B1(new_n1181), .B2(KEYINPUT57), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1175), .B1(new_n1180), .B2(new_n1182), .ZN(G375));
  OAI211_X1 g0983(.A(new_n1111), .B(new_n1117), .C1(new_n1112), .C2(new_n1114), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1119), .A2(new_n932), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n873), .A2(new_n771), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n704), .B1(G68), .B2(new_n794), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n723), .A2(new_n528), .B1(new_n205), .B2(new_n740), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G107), .B2(new_n738), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n287), .B1(new_n716), .B2(new_n754), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n726), .B2(G283), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n733), .A2(G116), .B1(G77), .B2(new_n735), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1189), .A2(new_n1014), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1193), .A2(KEYINPUT122), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n723), .A2(new_n1165), .B1(new_n717), .B2(new_n740), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1150), .B(new_n1195), .C1(G137), .C2(new_n726), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G50), .A2(new_n812), .B1(new_n738), .B2(G150), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT123), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n733), .A2(new_n1085), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n809), .B1(G128), .B2(new_n752), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1196), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1193), .A2(KEYINPUT122), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1194), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1187), .B1(new_n1203), .B2(new_n710), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1115), .A2(new_n703), .B1(new_n1186), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1185), .A2(new_n1205), .ZN(G381));
  OR4_X1    g1006(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1207), .A2(G387), .A3(G378), .A4(G390), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n1175), .C1(new_n1180), .C2(new_n1182), .ZN(G407));
  NAND2_X1  g1009(.A1(new_n628), .A2(G213), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1122), .A2(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(G407), .B(G213), .C1(G375), .C2(new_n1212), .ZN(G409));
  INV_X1    g1013(.A(KEYINPUT63), .ZN(new_n1214));
  OAI211_X1 g1014(.A(G378), .B(new_n1175), .C1(new_n1180), .C2(new_n1182), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1181), .A2(new_n932), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1179), .A2(new_n703), .A3(new_n1177), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1174), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1122), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1215), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1210), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1104), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT60), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1184), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT124), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1184), .B2(new_n1223), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1114), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1110), .A2(new_n1106), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1228), .A2(new_n1074), .B1(new_n1070), .B2(new_n1229), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1230), .A2(KEYINPUT124), .A3(KEYINPUT60), .A4(new_n1117), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1225), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1205), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n819), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1227), .A2(new_n1231), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1237), .A2(G384), .A3(new_n1205), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1214), .B1(new_n1221), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1211), .A2(G2897), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G384), .B1(new_n1237), .B2(new_n1205), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n819), .B(new_n1233), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1234), .A2(new_n1238), .A3(new_n1241), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT61), .B1(new_n1221), .B2(new_n1247), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n972), .A2(new_n999), .A3(G390), .ZN(new_n1249));
  AOI21_X1  g1049(.A(G390), .B1(new_n972), .B2(new_n999), .ZN(new_n1250));
  XOR2_X1   g1050(.A(G393), .B(G396), .Z(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1249), .A2(new_n1250), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(G390), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G387), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n972), .A2(new_n999), .A3(G390), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1251), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1253), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1211), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1239), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(KEYINPUT63), .A3(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1240), .A2(new_n1248), .A3(new_n1258), .A4(new_n1261), .ZN(new_n1262));
  XOR2_X1   g1062(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n1263));
  AND3_X1   g1063(.A1(new_n1259), .A2(new_n1260), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT61), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1265), .B1(new_n1259), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1264), .A2(new_n1267), .A3(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT126), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n1253), .B2(new_n1257), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1252), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1255), .A2(new_n1251), .A3(new_n1256), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(KEYINPUT126), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1262), .B1(new_n1270), .B2(new_n1276), .ZN(G405));
  NAND2_X1  g1077(.A1(G375), .A2(new_n1122), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1278), .A2(new_n1239), .A3(new_n1215), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1239), .B1(new_n1278), .B2(new_n1215), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1273), .A2(new_n1274), .A3(KEYINPUT126), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT126), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT127), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT127), .B1(new_n1272), .B2(new_n1275), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1281), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1284), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1272), .A2(KEYINPUT127), .A3(new_n1275), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1288), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1287), .A2(new_n1291), .ZN(G402));
endmodule


