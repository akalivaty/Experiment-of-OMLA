

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U561 ( .A1(n531), .A2(n528), .ZN(n914) );
  NOR2_X1 U562 ( .A1(KEYINPUT33), .A2(n794), .ZN(n796) );
  XNOR2_X1 U563 ( .A(n782), .B(KEYINPUT32), .ZN(n548) );
  OR2_X1 U564 ( .A1(n742), .A2(n743), .ZN(n534) );
  AND2_X1 U565 ( .A1(n575), .A2(G2105), .ZN(n918) );
  XNOR2_X1 U566 ( .A(n535), .B(KEYINPUT65), .ZN(n742) );
  NOR2_X1 U567 ( .A1(n737), .A2(n1004), .ZN(n535) );
  AND2_X1 U568 ( .A1(n542), .A2(n540), .ZN(n539) );
  NAND2_X1 U569 ( .A1(n543), .A2(KEYINPUT29), .ZN(n542) );
  AND2_X1 U570 ( .A1(n754), .A2(n755), .ZN(n541) );
  AND2_X1 U571 ( .A1(n537), .A2(n760), .ZN(n536) );
  NAND2_X1 U572 ( .A1(n538), .A2(KEYINPUT29), .ZN(n537) );
  AND2_X1 U573 ( .A1(n1002), .A2(n792), .ZN(n793) );
  XNOR2_X1 U574 ( .A(n727), .B(n726), .ZN(n828) );
  AND2_X1 U575 ( .A1(n725), .A2(n724), .ZN(n727) );
  NOR2_X1 U576 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n533) );
  INV_X1 U577 ( .A(G2105), .ZN(n532) );
  NAND2_X1 U578 ( .A1(G2105), .A2(KEYINPUT17), .ZN(n529) );
  NAND2_X1 U579 ( .A1(n552), .A2(n526), .ZN(n551) );
  XNOR2_X1 U580 ( .A(n769), .B(KEYINPUT31), .ZN(n770) );
  NOR2_X1 U581 ( .A1(n728), .A2(G1384), .ZN(n729) );
  NAND2_X1 U582 ( .A1(n548), .A2(n525), .ZN(n547) );
  NAND2_X1 U583 ( .A1(n793), .A2(n546), .ZN(n545) );
  INV_X1 U584 ( .A(n1011), .ZN(n546) );
  INV_X1 U585 ( .A(KEYINPUT97), .ZN(n587) );
  AND2_X1 U586 ( .A1(n530), .A2(n529), .ZN(n528) );
  NAND2_X1 U587 ( .A1(n533), .A2(n532), .ZN(n531) );
  NAND2_X1 U588 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n530) );
  AND2_X1 U589 ( .A1(G2104), .A2(G2105), .ZN(n920) );
  XNOR2_X1 U590 ( .A(KEYINPUT68), .B(KEYINPUT23), .ZN(n576) );
  XNOR2_X1 U591 ( .A(n550), .B(n549), .ZN(G329) );
  INV_X1 U592 ( .A(KEYINPUT40), .ZN(n549) );
  NAND2_X1 U593 ( .A1(n551), .A2(n527), .ZN(n550) );
  AND2_X1 U594 ( .A1(n789), .A2(n793), .ZN(n525) );
  BUF_X1 U595 ( .A(n732), .Z(n774) );
  NAND2_X1 U596 ( .A1(n773), .A2(n772), .ZN(n784) );
  AND2_X1 U597 ( .A1(n851), .A2(n553), .ZN(n526) );
  NAND2_X1 U598 ( .A1(n860), .A2(n859), .ZN(n527) );
  INV_X1 U599 ( .A(KEYINPUT29), .ZN(n755) );
  NAND2_X1 U600 ( .A1(n534), .A2(n741), .ZN(n745) );
  NAND2_X1 U601 ( .A1(n539), .A2(n536), .ZN(n773) );
  INV_X1 U602 ( .A(n754), .ZN(n538) );
  NAND2_X1 U603 ( .A1(n544), .A2(n541), .ZN(n540) );
  INV_X1 U604 ( .A(n544), .ZN(n543) );
  NAND2_X1 U605 ( .A1(n751), .A2(n750), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n548), .A2(n789), .ZN(n803) );
  NAND2_X1 U607 ( .A1(n547), .A2(n545), .ZN(n794) );
  NAND2_X1 U608 ( .A1(n802), .A2(n801), .ZN(n552) );
  NOR2_X1 U609 ( .A1(G2105), .A2(n575), .ZN(n599) );
  XNOR2_X1 U610 ( .A(n588), .B(n587), .ZN(n594) );
  NAND2_X1 U611 ( .A1(n914), .A2(G138), .ZN(n588) );
  NOR2_X1 U612 ( .A1(n850), .A2(n849), .ZN(n553) );
  INV_X1 U613 ( .A(KEYINPUT110), .ZN(n769) );
  XNOR2_X1 U614 ( .A(n771), .B(n770), .ZN(n772) );
  INV_X1 U615 ( .A(n809), .ZN(n792) );
  XNOR2_X1 U616 ( .A(n577), .B(n576), .ZN(n722) );
  XOR2_X1 U617 ( .A(KEYINPUT0), .B(G543), .Z(n674) );
  INV_X1 U618 ( .A(G651), .ZN(n559) );
  NOR2_X1 U619 ( .A1(n674), .A2(n559), .ZN(n687) );
  NAND2_X1 U620 ( .A1(n687), .A2(G76), .ZN(n554) );
  XNOR2_X1 U621 ( .A(KEYINPUT82), .B(n554), .ZN(n557) );
  NOR2_X1 U622 ( .A1(G651), .A2(G543), .ZN(n686) );
  NAND2_X1 U623 ( .A1(n686), .A2(G89), .ZN(n555) );
  XNOR2_X1 U624 ( .A(KEYINPUT4), .B(n555), .ZN(n556) );
  NAND2_X1 U625 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(KEYINPUT5), .B(n558), .ZN(n568) );
  XNOR2_X1 U627 ( .A(KEYINPUT6), .B(KEYINPUT84), .ZN(n566) );
  NOR2_X1 U628 ( .A1(G543), .A2(n559), .ZN(n560) );
  XOR2_X1 U629 ( .A(KEYINPUT1), .B(n560), .Z(n690) );
  NAND2_X1 U630 ( .A1(n690), .A2(G63), .ZN(n564) );
  NOR2_X1 U631 ( .A1(G651), .A2(n674), .ZN(n561) );
  XNOR2_X1 U632 ( .A(KEYINPUT66), .B(n561), .ZN(n691) );
  NAND2_X1 U633 ( .A1(G51), .A2(n691), .ZN(n562) );
  XOR2_X1 U634 ( .A(KEYINPUT83), .B(n562), .Z(n563) );
  NAND2_X1 U635 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U636 ( .A(n566), .B(n565), .Z(n567) );
  NAND2_X1 U637 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U638 ( .A(KEYINPUT7), .B(n569), .ZN(G168) );
  XOR2_X1 U639 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U640 ( .A1(G137), .A2(n914), .ZN(n571) );
  NAND2_X1 U641 ( .A1(G113), .A2(n920), .ZN(n570) );
  NAND2_X1 U642 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U643 ( .A(n572), .B(KEYINPUT69), .ZN(n574) );
  XNOR2_X1 U644 ( .A(G2104), .B(KEYINPUT67), .ZN(n575) );
  NAND2_X1 U645 ( .A1(G125), .A2(n918), .ZN(n573) );
  AND2_X1 U646 ( .A1(n574), .A2(n573), .ZN(n724) );
  NAND2_X1 U647 ( .A1(G101), .A2(n599), .ZN(n577) );
  INV_X1 U648 ( .A(n722), .ZN(n578) );
  AND2_X1 U649 ( .A1(n724), .A2(n578), .ZN(G160) );
  NAND2_X1 U650 ( .A1(G90), .A2(n686), .ZN(n580) );
  NAND2_X1 U651 ( .A1(G77), .A2(n687), .ZN(n579) );
  NAND2_X1 U652 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U653 ( .A(KEYINPUT9), .B(n581), .ZN(n586) );
  NAND2_X1 U654 ( .A1(G64), .A2(n690), .ZN(n583) );
  NAND2_X1 U655 ( .A1(G52), .A2(n691), .ZN(n582) );
  NAND2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U657 ( .A(KEYINPUT73), .B(n584), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(G301) );
  INV_X1 U659 ( .A(G301), .ZN(G171) );
  AND2_X1 U660 ( .A1(n920), .A2(G114), .ZN(n592) );
  NAND2_X1 U661 ( .A1(G102), .A2(n599), .ZN(n590) );
  NAND2_X1 U662 ( .A1(G126), .A2(n918), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n594), .A2(n593), .ZN(n596) );
  INV_X1 U666 ( .A(KEYINPUT98), .ZN(n595) );
  XNOR2_X1 U667 ( .A(n596), .B(n595), .ZN(n728) );
  BUF_X1 U668 ( .A(n728), .Z(G164) );
  AND2_X1 U669 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U670 ( .A1(G111), .A2(n920), .ZN(n606) );
  NAND2_X1 U671 ( .A1(G123), .A2(n918), .ZN(n597) );
  XNOR2_X1 U672 ( .A(n597), .B(KEYINPUT86), .ZN(n598) );
  XNOR2_X1 U673 ( .A(n598), .B(KEYINPUT18), .ZN(n601) );
  BUF_X1 U674 ( .A(n599), .Z(n915) );
  NAND2_X1 U675 ( .A1(G99), .A2(n915), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U677 ( .A1(G135), .A2(n914), .ZN(n602) );
  XNOR2_X1 U678 ( .A(KEYINPUT87), .B(n602), .ZN(n603) );
  NOR2_X1 U679 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U681 ( .A(n607), .B(KEYINPUT88), .ZN(n952) );
  XNOR2_X1 U682 ( .A(n952), .B(G2096), .ZN(n608) );
  OR2_X1 U683 ( .A1(G2100), .A2(n608), .ZN(G156) );
  INV_X1 U684 ( .A(G132), .ZN(G219) );
  INV_X1 U685 ( .A(G82), .ZN(G220) );
  NAND2_X1 U686 ( .A1(G7), .A2(G661), .ZN(n609) );
  XNOR2_X1 U687 ( .A(n609), .B(KEYINPUT76), .ZN(n610) );
  XNOR2_X1 U688 ( .A(KEYINPUT10), .B(n610), .ZN(G223) );
  INV_X1 U689 ( .A(G223), .ZN(n861) );
  NAND2_X1 U690 ( .A1(n861), .A2(G567), .ZN(n611) );
  XOR2_X1 U691 ( .A(KEYINPUT11), .B(n611), .Z(G234) );
  NAND2_X1 U692 ( .A1(n690), .A2(G56), .ZN(n612) );
  XNOR2_X1 U693 ( .A(KEYINPUT14), .B(n612), .ZN(n623) );
  XNOR2_X1 U694 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n686), .A2(G81), .ZN(n613) );
  XNOR2_X1 U696 ( .A(n613), .B(KEYINPUT12), .ZN(n615) );
  NAND2_X1 U697 ( .A1(G68), .A2(n687), .ZN(n614) );
  NAND2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U699 ( .A(n616), .B(KEYINPUT13), .ZN(n617) );
  XNOR2_X1 U700 ( .A(n618), .B(n617), .ZN(n621) );
  NAND2_X1 U701 ( .A1(G43), .A2(n691), .ZN(n619) );
  XNOR2_X1 U702 ( .A(KEYINPUT79), .B(n619), .ZN(n620) );
  NOR2_X1 U703 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n1004) );
  INV_X1 U705 ( .A(G860), .ZN(n644) );
  OR2_X1 U706 ( .A1(n1004), .A2(n644), .ZN(G153) );
  INV_X1 U707 ( .A(G868), .ZN(n705) );
  NOR2_X1 U708 ( .A1(G171), .A2(n705), .ZN(n624) );
  XOR2_X1 U709 ( .A(KEYINPUT80), .B(n624), .Z(n634) );
  NAND2_X1 U710 ( .A1(G92), .A2(n686), .ZN(n626) );
  NAND2_X1 U711 ( .A1(G66), .A2(n690), .ZN(n625) );
  NAND2_X1 U712 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U713 ( .A1(G79), .A2(n687), .ZN(n628) );
  NAND2_X1 U714 ( .A1(G54), .A2(n691), .ZN(n627) );
  NAND2_X1 U715 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U716 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U717 ( .A(KEYINPUT15), .B(n631), .Z(n1010) );
  NOR2_X1 U718 ( .A1(n1010), .A2(G868), .ZN(n632) );
  XNOR2_X1 U719 ( .A(KEYINPUT81), .B(n632), .ZN(n633) );
  NAND2_X1 U720 ( .A1(n634), .A2(n633), .ZN(G284) );
  NAND2_X1 U721 ( .A1(G91), .A2(n686), .ZN(n636) );
  NAND2_X1 U722 ( .A1(G65), .A2(n690), .ZN(n635) );
  NAND2_X1 U723 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U724 ( .A1(n687), .A2(G78), .ZN(n637) );
  XOR2_X1 U725 ( .A(KEYINPUT74), .B(n637), .Z(n638) );
  NOR2_X1 U726 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U727 ( .A1(G53), .A2(n691), .ZN(n640) );
  NAND2_X1 U728 ( .A1(n641), .A2(n640), .ZN(G299) );
  NOR2_X1 U729 ( .A1(G286), .A2(n705), .ZN(n643) );
  NOR2_X1 U730 ( .A1(G868), .A2(G299), .ZN(n642) );
  NOR2_X1 U731 ( .A1(n643), .A2(n642), .ZN(G297) );
  NAND2_X1 U732 ( .A1(n644), .A2(G559), .ZN(n645) );
  NAND2_X1 U733 ( .A1(n645), .A2(n1010), .ZN(n646) );
  XNOR2_X1 U734 ( .A(n646), .B(KEYINPUT85), .ZN(n647) );
  XOR2_X1 U735 ( .A(KEYINPUT16), .B(n647), .Z(G148) );
  NOR2_X1 U736 ( .A1(G868), .A2(n1004), .ZN(n650) );
  NAND2_X1 U737 ( .A1(G868), .A2(n1010), .ZN(n648) );
  NOR2_X1 U738 ( .A1(G559), .A2(n648), .ZN(n649) );
  NOR2_X1 U739 ( .A1(n650), .A2(n649), .ZN(G282) );
  NAND2_X1 U740 ( .A1(G559), .A2(n1010), .ZN(n651) );
  XNOR2_X1 U741 ( .A(n651), .B(n1004), .ZN(n702) );
  NOR2_X1 U742 ( .A1(n702), .A2(G860), .ZN(n660) );
  NAND2_X1 U743 ( .A1(G93), .A2(n686), .ZN(n653) );
  NAND2_X1 U744 ( .A1(G67), .A2(n690), .ZN(n652) );
  NAND2_X1 U745 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U746 ( .A1(G80), .A2(n687), .ZN(n654) );
  XNOR2_X1 U747 ( .A(KEYINPUT89), .B(n654), .ZN(n655) );
  NOR2_X1 U748 ( .A1(n656), .A2(n655), .ZN(n658) );
  NAND2_X1 U749 ( .A1(G55), .A2(n691), .ZN(n657) );
  NAND2_X1 U750 ( .A1(n658), .A2(n657), .ZN(n704) );
  XOR2_X1 U751 ( .A(n704), .B(KEYINPUT90), .Z(n659) );
  XNOR2_X1 U752 ( .A(n660), .B(n659), .ZN(G145) );
  NAND2_X1 U753 ( .A1(G73), .A2(n687), .ZN(n661) );
  XNOR2_X1 U754 ( .A(n661), .B(KEYINPUT2), .ZN(n669) );
  NAND2_X1 U755 ( .A1(G61), .A2(n690), .ZN(n662) );
  XNOR2_X1 U756 ( .A(n662), .B(KEYINPUT92), .ZN(n664) );
  NAND2_X1 U757 ( .A1(n686), .A2(G86), .ZN(n663) );
  NAND2_X1 U758 ( .A1(n664), .A2(n663), .ZN(n667) );
  NAND2_X1 U759 ( .A1(G48), .A2(n691), .ZN(n665) );
  XNOR2_X1 U760 ( .A(KEYINPUT93), .B(n665), .ZN(n666) );
  NOR2_X1 U761 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U762 ( .A1(n669), .A2(n668), .ZN(G305) );
  NAND2_X1 U763 ( .A1(G651), .A2(G74), .ZN(n671) );
  NAND2_X1 U764 ( .A1(G49), .A2(n691), .ZN(n670) );
  NAND2_X1 U765 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U766 ( .A1(n690), .A2(n672), .ZN(n673) );
  XOR2_X1 U767 ( .A(KEYINPUT91), .B(n673), .Z(n676) );
  NAND2_X1 U768 ( .A1(n674), .A2(G87), .ZN(n675) );
  NAND2_X1 U769 ( .A1(n676), .A2(n675), .ZN(G288) );
  NAND2_X1 U770 ( .A1(n687), .A2(G72), .ZN(n677) );
  XNOR2_X1 U771 ( .A(KEYINPUT71), .B(n677), .ZN(n680) );
  NAND2_X1 U772 ( .A1(n686), .A2(G85), .ZN(n678) );
  XOR2_X1 U773 ( .A(KEYINPUT70), .B(n678), .Z(n679) );
  NOR2_X1 U774 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U775 ( .A(KEYINPUT72), .B(n681), .ZN(n685) );
  NAND2_X1 U776 ( .A1(n691), .A2(G47), .ZN(n683) );
  NAND2_X1 U777 ( .A1(G60), .A2(n690), .ZN(n682) );
  AND2_X1 U778 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U779 ( .A1(n685), .A2(n684), .ZN(G290) );
  NAND2_X1 U780 ( .A1(G88), .A2(n686), .ZN(n689) );
  NAND2_X1 U781 ( .A1(G75), .A2(n687), .ZN(n688) );
  NAND2_X1 U782 ( .A1(n689), .A2(n688), .ZN(n695) );
  NAND2_X1 U783 ( .A1(G62), .A2(n690), .ZN(n693) );
  NAND2_X1 U784 ( .A1(G50), .A2(n691), .ZN(n692) );
  NAND2_X1 U785 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U786 ( .A1(n695), .A2(n694), .ZN(G166) );
  XOR2_X1 U787 ( .A(KEYINPUT19), .B(KEYINPUT94), .Z(n696) );
  XNOR2_X1 U788 ( .A(G305), .B(n696), .ZN(n699) );
  INV_X1 U789 ( .A(G299), .ZN(n1007) );
  XNOR2_X1 U790 ( .A(n1007), .B(G288), .ZN(n697) );
  XNOR2_X1 U791 ( .A(n697), .B(n704), .ZN(n698) );
  XNOR2_X1 U792 ( .A(n699), .B(n698), .ZN(n701) );
  XNOR2_X1 U793 ( .A(G290), .B(G166), .ZN(n700) );
  XNOR2_X1 U794 ( .A(n701), .B(n700), .ZN(n930) );
  XNOR2_X1 U795 ( .A(n702), .B(n930), .ZN(n703) );
  NAND2_X1 U796 ( .A1(n703), .A2(G868), .ZN(n707) );
  NAND2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U798 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U799 ( .A(KEYINPUT95), .B(n708), .Z(G295) );
  NAND2_X1 U800 ( .A1(G2084), .A2(G2078), .ZN(n709) );
  XOR2_X1 U801 ( .A(KEYINPUT20), .B(n709), .Z(n710) );
  NAND2_X1 U802 ( .A1(G2090), .A2(n710), .ZN(n711) );
  XNOR2_X1 U803 ( .A(KEYINPUT21), .B(n711), .ZN(n712) );
  NAND2_X1 U804 ( .A1(n712), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U805 ( .A(KEYINPUT75), .B(G57), .ZN(G237) );
  XNOR2_X1 U806 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U807 ( .A1(G108), .A2(G120), .ZN(n713) );
  NOR2_X1 U808 ( .A1(G237), .A2(n713), .ZN(n714) );
  NAND2_X1 U809 ( .A1(G69), .A2(n714), .ZN(n867) );
  NAND2_X1 U810 ( .A1(n867), .A2(G567), .ZN(n720) );
  NOR2_X1 U811 ( .A1(G220), .A2(G219), .ZN(n715) );
  XNOR2_X1 U812 ( .A(KEYINPUT22), .B(n715), .ZN(n716) );
  NAND2_X1 U813 ( .A1(n716), .A2(G96), .ZN(n717) );
  NOR2_X1 U814 ( .A1(G218), .A2(n717), .ZN(n718) );
  XOR2_X1 U815 ( .A(KEYINPUT96), .B(n718), .Z(n868) );
  NAND2_X1 U816 ( .A1(n868), .A2(G2106), .ZN(n719) );
  NAND2_X1 U817 ( .A1(n720), .A2(n719), .ZN(n869) );
  NAND2_X1 U818 ( .A1(G661), .A2(G483), .ZN(n721) );
  NOR2_X1 U819 ( .A1(n869), .A2(n721), .ZN(n865) );
  NAND2_X1 U820 ( .A1(n865), .A2(G36), .ZN(G176) );
  INV_X1 U821 ( .A(G166), .ZN(G303) );
  INV_X1 U822 ( .A(KEYINPUT107), .ZN(n736) );
  INV_X1 U823 ( .A(G40), .ZN(n723) );
  NOR2_X1 U824 ( .A1(n723), .A2(n722), .ZN(n725) );
  INV_X1 U825 ( .A(KEYINPUT99), .ZN(n726) );
  XNOR2_X1 U826 ( .A(n729), .B(KEYINPUT64), .ZN(n827) );
  NAND2_X1 U827 ( .A1(n828), .A2(n827), .ZN(n732) );
  INV_X1 U828 ( .A(n732), .ZN(n730) );
  NAND2_X1 U829 ( .A1(n730), .A2(G1996), .ZN(n731) );
  XNOR2_X1 U830 ( .A(n731), .B(KEYINPUT26), .ZN(n734) );
  NAND2_X1 U831 ( .A1(G1341), .A2(n774), .ZN(n733) );
  NAND2_X1 U832 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U833 ( .A(n736), .B(n735), .ZN(n737) );
  INV_X1 U834 ( .A(n1010), .ZN(n743) );
  NAND2_X1 U835 ( .A1(n774), .A2(G1348), .ZN(n738) );
  XNOR2_X1 U836 ( .A(n738), .B(KEYINPUT108), .ZN(n740) );
  NAND2_X1 U837 ( .A1(n730), .A2(G2067), .ZN(n739) );
  NAND2_X1 U838 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U839 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U840 ( .A1(n745), .A2(n744), .ZN(n751) );
  NAND2_X1 U841 ( .A1(G2072), .A2(n730), .ZN(n747) );
  XNOR2_X1 U842 ( .A(KEYINPUT106), .B(KEYINPUT27), .ZN(n746) );
  XNOR2_X1 U843 ( .A(n747), .B(n746), .ZN(n749) );
  INV_X1 U844 ( .A(G1956), .ZN(n1024) );
  NOR2_X1 U845 ( .A1(n730), .A2(n1024), .ZN(n748) );
  NOR2_X1 U846 ( .A1(n749), .A2(n748), .ZN(n752) );
  NAND2_X1 U847 ( .A1(n1007), .A2(n752), .ZN(n750) );
  NOR2_X1 U848 ( .A1(n1007), .A2(n752), .ZN(n753) );
  XOR2_X1 U849 ( .A(n753), .B(KEYINPUT28), .Z(n754) );
  XOR2_X1 U850 ( .A(G2078), .B(KEYINPUT25), .Z(n756) );
  XNOR2_X1 U851 ( .A(KEYINPUT104), .B(n756), .ZN(n979) );
  NOR2_X1 U852 ( .A1(n774), .A2(n979), .ZN(n757) );
  XNOR2_X1 U853 ( .A(n757), .B(KEYINPUT105), .ZN(n759) );
  INV_X1 U854 ( .A(G1961), .ZN(n1023) );
  NAND2_X1 U855 ( .A1(n1023), .A2(n774), .ZN(n758) );
  NAND2_X1 U856 ( .A1(n759), .A2(n758), .ZN(n761) );
  NAND2_X1 U857 ( .A1(n761), .A2(G171), .ZN(n760) );
  OR2_X1 U858 ( .A1(n761), .A2(G171), .ZN(n762) );
  XNOR2_X1 U859 ( .A(n762), .B(KEYINPUT109), .ZN(n768) );
  NAND2_X1 U860 ( .A1(G8), .A2(n774), .ZN(n809) );
  NOR2_X1 U861 ( .A1(G1966), .A2(n809), .ZN(n786) );
  NOR2_X1 U862 ( .A1(G2084), .A2(n774), .ZN(n763) );
  XOR2_X1 U863 ( .A(KEYINPUT103), .B(n763), .Z(n783) );
  NOR2_X1 U864 ( .A1(n786), .A2(n783), .ZN(n764) );
  NAND2_X1 U865 ( .A1(G8), .A2(n764), .ZN(n765) );
  XNOR2_X1 U866 ( .A(n765), .B(KEYINPUT30), .ZN(n766) );
  NOR2_X1 U867 ( .A1(n766), .A2(G168), .ZN(n767) );
  NOR2_X1 U868 ( .A1(n768), .A2(n767), .ZN(n771) );
  NAND2_X1 U869 ( .A1(n784), .A2(G286), .ZN(n779) );
  NOR2_X1 U870 ( .A1(G2090), .A2(n774), .ZN(n776) );
  NOR2_X1 U871 ( .A1(G1971), .A2(n809), .ZN(n775) );
  NOR2_X1 U872 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U873 ( .A1(n777), .A2(G303), .ZN(n778) );
  NAND2_X1 U874 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U875 ( .A(n780), .B(KEYINPUT112), .ZN(n781) );
  NAND2_X1 U876 ( .A1(n781), .A2(G8), .ZN(n782) );
  NAND2_X1 U877 ( .A1(G8), .A2(n783), .ZN(n788) );
  XNOR2_X1 U878 ( .A(KEYINPUT111), .B(n784), .ZN(n785) );
  NOR2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U881 ( .A1(G1976), .A2(G288), .ZN(n797) );
  NOR2_X1 U882 ( .A1(G1971), .A2(G303), .ZN(n790) );
  NOR2_X1 U883 ( .A1(n797), .A2(n790), .ZN(n1011) );
  NAND2_X1 U884 ( .A1(G288), .A2(G1976), .ZN(n791) );
  XOR2_X1 U885 ( .A(KEYINPUT113), .B(n791), .Z(n1002) );
  INV_X1 U886 ( .A(KEYINPUT114), .ZN(n795) );
  XNOR2_X1 U887 ( .A(n796), .B(n795), .ZN(n802) );
  NAND2_X1 U888 ( .A1(n797), .A2(KEYINPUT33), .ZN(n798) );
  NOR2_X1 U889 ( .A1(n809), .A2(n798), .ZN(n800) );
  XOR2_X1 U890 ( .A(G1981), .B(G305), .Z(n999) );
  INV_X1 U891 ( .A(n999), .ZN(n799) );
  NOR2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U893 ( .A1(G2090), .A2(G303), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G8), .A2(n804), .ZN(n805) );
  NAND2_X1 U895 ( .A1(n803), .A2(n805), .ZN(n806) );
  NAND2_X1 U896 ( .A1(n806), .A2(n809), .ZN(n851) );
  NOR2_X1 U897 ( .A1(G1981), .A2(G305), .ZN(n807) );
  XOR2_X1 U898 ( .A(n807), .B(KEYINPUT24), .Z(n808) );
  NOR2_X1 U899 ( .A1(n809), .A2(n808), .ZN(n850) );
  NAND2_X1 U900 ( .A1(G141), .A2(n914), .ZN(n811) );
  NAND2_X1 U901 ( .A1(G117), .A2(n920), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n811), .A2(n810), .ZN(n814) );
  NAND2_X1 U903 ( .A1(n915), .A2(G105), .ZN(n812) );
  XOR2_X1 U904 ( .A(KEYINPUT38), .B(n812), .Z(n813) );
  NOR2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U906 ( .A1(n918), .A2(G129), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n900) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n900), .ZN(n960) );
  NAND2_X1 U909 ( .A1(G107), .A2(n920), .ZN(n817) );
  XNOR2_X1 U910 ( .A(n817), .B(KEYINPUT100), .ZN(n820) );
  NAND2_X1 U911 ( .A1(G95), .A2(n915), .ZN(n818) );
  XOR2_X1 U912 ( .A(KEYINPUT101), .B(n818), .Z(n819) );
  NAND2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n824) );
  NAND2_X1 U914 ( .A1(G131), .A2(n914), .ZN(n822) );
  NAND2_X1 U915 ( .A1(G119), .A2(n918), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n823) );
  OR2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n896) );
  AND2_X1 U918 ( .A1(n896), .A2(G1991), .ZN(n826) );
  AND2_X1 U919 ( .A1(G1996), .A2(n900), .ZN(n825) );
  NOR2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n958) );
  INV_X1 U921 ( .A(n828), .ZN(n829) );
  NOR2_X1 U922 ( .A1(n827), .A2(n829), .ZN(n847) );
  INV_X1 U923 ( .A(n847), .ZN(n852) );
  NOR2_X1 U924 ( .A1(n958), .A2(n852), .ZN(n853) );
  NOR2_X1 U925 ( .A1(G1991), .A2(n896), .ZN(n955) );
  NOR2_X1 U926 ( .A1(G1986), .A2(G290), .ZN(n830) );
  NOR2_X1 U927 ( .A1(n955), .A2(n830), .ZN(n831) );
  NOR2_X1 U928 ( .A1(n853), .A2(n831), .ZN(n832) );
  XOR2_X1 U929 ( .A(KEYINPUT115), .B(n832), .Z(n833) );
  NOR2_X1 U930 ( .A1(n960), .A2(n833), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n834), .B(KEYINPUT39), .ZN(n844) );
  XNOR2_X1 U932 ( .A(G2067), .B(KEYINPUT37), .ZN(n845) );
  NAND2_X1 U933 ( .A1(G140), .A2(n914), .ZN(n836) );
  NAND2_X1 U934 ( .A1(G104), .A2(n915), .ZN(n835) );
  NAND2_X1 U935 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U936 ( .A(KEYINPUT34), .B(n837), .ZN(n842) );
  NAND2_X1 U937 ( .A1(G128), .A2(n918), .ZN(n839) );
  NAND2_X1 U938 ( .A1(G116), .A2(n920), .ZN(n838) );
  NAND2_X1 U939 ( .A1(n839), .A2(n838), .ZN(n840) );
  XOR2_X1 U940 ( .A(KEYINPUT35), .B(n840), .Z(n841) );
  NOR2_X1 U941 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U942 ( .A(KEYINPUT36), .B(n843), .ZN(n910) );
  NOR2_X1 U943 ( .A1(n845), .A2(n910), .ZN(n956) );
  NAND2_X1 U944 ( .A1(n847), .A2(n956), .ZN(n855) );
  NAND2_X1 U945 ( .A1(n844), .A2(n855), .ZN(n846) );
  NAND2_X1 U946 ( .A1(n845), .A2(n910), .ZN(n951) );
  NAND2_X1 U947 ( .A1(n846), .A2(n951), .ZN(n848) );
  NAND2_X1 U948 ( .A1(n848), .A2(n847), .ZN(n860) );
  INV_X1 U949 ( .A(n860), .ZN(n849) );
  XOR2_X1 U950 ( .A(G1986), .B(G290), .Z(n1003) );
  NOR2_X1 U951 ( .A1(n1003), .A2(n852), .ZN(n858) );
  INV_X1 U952 ( .A(n853), .ZN(n854) );
  NAND2_X1 U953 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n856), .B(KEYINPUT102), .ZN(n857) );
  OR2_X1 U955 ( .A1(n858), .A2(n857), .ZN(n859) );
  NAND2_X1 U956 ( .A1(n861), .A2(G2106), .ZN(n862) );
  XOR2_X1 U957 ( .A(KEYINPUT117), .B(n862), .Z(G217) );
  AND2_X1 U958 ( .A1(G15), .A2(G2), .ZN(n863) );
  NAND2_X1 U959 ( .A1(G661), .A2(n863), .ZN(G259) );
  NAND2_X1 U960 ( .A1(G3), .A2(G1), .ZN(n864) );
  XNOR2_X1 U961 ( .A(KEYINPUT118), .B(n864), .ZN(n866) );
  NAND2_X1 U962 ( .A1(n866), .A2(n865), .ZN(G188) );
  XNOR2_X1 U963 ( .A(G96), .B(KEYINPUT119), .ZN(G221) );
  NOR2_X1 U964 ( .A1(n868), .A2(n867), .ZN(G325) );
  XOR2_X1 U965 ( .A(KEYINPUT120), .B(G325), .Z(G261) );
  INV_X1 U967 ( .A(G120), .ZN(G236) );
  INV_X1 U968 ( .A(G108), .ZN(G238) );
  INV_X1 U969 ( .A(G69), .ZN(G235) );
  INV_X1 U970 ( .A(n869), .ZN(G319) );
  XOR2_X1 U971 ( .A(KEYINPUT121), .B(G2090), .Z(n871) );
  XNOR2_X1 U972 ( .A(G2067), .B(G2084), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(n872), .B(G2100), .Z(n874) );
  XNOR2_X1 U975 ( .A(G2078), .B(G2072), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U977 ( .A(G2096), .B(KEYINPUT43), .Z(n876) );
  XNOR2_X1 U978 ( .A(G2678), .B(KEYINPUT42), .ZN(n875) );
  XNOR2_X1 U979 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U980 ( .A(n878), .B(n877), .Z(G227) );
  XNOR2_X1 U981 ( .A(G1961), .B(G2474), .ZN(n888) );
  XOR2_X1 U982 ( .A(G1976), .B(G1971), .Z(n880) );
  XNOR2_X1 U983 ( .A(G1986), .B(G1956), .ZN(n879) );
  XNOR2_X1 U984 ( .A(n880), .B(n879), .ZN(n884) );
  XOR2_X1 U985 ( .A(G1981), .B(G1966), .Z(n882) );
  XNOR2_X1 U986 ( .A(G1996), .B(G1991), .ZN(n881) );
  XNOR2_X1 U987 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U988 ( .A(n884), .B(n883), .Z(n886) );
  XNOR2_X1 U989 ( .A(KEYINPUT122), .B(KEYINPUT41), .ZN(n885) );
  XNOR2_X1 U990 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U991 ( .A(n888), .B(n887), .ZN(G229) );
  NAND2_X1 U992 ( .A1(G136), .A2(n914), .ZN(n890) );
  NAND2_X1 U993 ( .A1(G112), .A2(n920), .ZN(n889) );
  NAND2_X1 U994 ( .A1(n890), .A2(n889), .ZN(n895) );
  NAND2_X1 U995 ( .A1(G124), .A2(n918), .ZN(n891) );
  XNOR2_X1 U996 ( .A(n891), .B(KEYINPUT44), .ZN(n893) );
  NAND2_X1 U997 ( .A1(n915), .A2(G100), .ZN(n892) );
  NAND2_X1 U998 ( .A1(n893), .A2(n892), .ZN(n894) );
  NOR2_X1 U999 ( .A1(n895), .A2(n894), .ZN(G162) );
  XNOR2_X1 U1000 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n898) );
  XOR2_X1 U1001 ( .A(G164), .B(n896), .Z(n897) );
  XNOR2_X1 U1002 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U1003 ( .A(n899), .B(n952), .Z(n902) );
  XOR2_X1 U1004 ( .A(n900), .B(G162), .Z(n901) );
  XNOR2_X1 U1005 ( .A(n902), .B(n901), .ZN(n913) );
  NAND2_X1 U1006 ( .A1(G130), .A2(n918), .ZN(n904) );
  NAND2_X1 U1007 ( .A1(G118), .A2(n920), .ZN(n903) );
  NAND2_X1 U1008 ( .A1(n904), .A2(n903), .ZN(n909) );
  NAND2_X1 U1009 ( .A1(G142), .A2(n914), .ZN(n906) );
  NAND2_X1 U1010 ( .A1(G106), .A2(n915), .ZN(n905) );
  NAND2_X1 U1011 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1012 ( .A(n907), .B(KEYINPUT45), .Z(n908) );
  NOR2_X1 U1013 ( .A1(n909), .A2(n908), .ZN(n911) );
  XNOR2_X1 U1014 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1015 ( .A(n913), .B(n912), .Z(n928) );
  NAND2_X1 U1016 ( .A1(G139), .A2(n914), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(G103), .A2(n915), .ZN(n916) );
  NAND2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n925) );
  NAND2_X1 U1019 ( .A1(n918), .A2(G127), .ZN(n919) );
  XOR2_X1 U1020 ( .A(KEYINPUT123), .B(n919), .Z(n922) );
  NAND2_X1 U1021 ( .A1(n920), .A2(G115), .ZN(n921) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1023 ( .A(KEYINPUT47), .B(n923), .Z(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1025 ( .A(KEYINPUT124), .B(n926), .Z(n966) );
  XNOR2_X1 U1026 ( .A(G160), .B(n966), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(n928), .B(n927), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(G37), .A2(n929), .ZN(G395) );
  XNOR2_X1 U1029 ( .A(n1004), .B(n930), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(G171), .B(n1010), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(n932), .B(n931), .ZN(n933) );
  XOR2_X1 U1032 ( .A(G286), .B(n933), .Z(n934) );
  NOR2_X1 U1033 ( .A1(G37), .A2(n934), .ZN(G397) );
  XOR2_X1 U1034 ( .A(KEYINPUT116), .B(G2446), .Z(n936) );
  XNOR2_X1 U1035 ( .A(G2443), .B(G2454), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(n936), .B(n935), .ZN(n937) );
  XOR2_X1 U1037 ( .A(n937), .B(G2451), .Z(n939) );
  XNOR2_X1 U1038 ( .A(G1348), .B(G1341), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(n939), .B(n938), .ZN(n943) );
  XOR2_X1 U1040 ( .A(G2435), .B(G2427), .Z(n941) );
  XNOR2_X1 U1041 ( .A(G2430), .B(G2438), .ZN(n940) );
  XNOR2_X1 U1042 ( .A(n941), .B(n940), .ZN(n942) );
  XOR2_X1 U1043 ( .A(n943), .B(n942), .Z(n944) );
  NAND2_X1 U1044 ( .A1(G14), .A2(n944), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(G319), .A2(n950), .ZN(n947) );
  NOR2_X1 U1046 ( .A1(G227), .A2(G229), .ZN(n945) );
  XNOR2_X1 U1047 ( .A(KEYINPUT49), .B(n945), .ZN(n946) );
  NOR2_X1 U1048 ( .A1(n947), .A2(n946), .ZN(n949) );
  NOR2_X1 U1049 ( .A1(G395), .A2(G397), .ZN(n948) );
  NAND2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(G225) );
  INV_X1 U1051 ( .A(G225), .ZN(G308) );
  INV_X1 U1052 ( .A(n950), .ZN(G401) );
  NAND2_X1 U1053 ( .A1(n952), .A2(n951), .ZN(n954) );
  XOR2_X1 U1054 ( .A(G160), .B(G2084), .Z(n953) );
  NOR2_X1 U1055 ( .A1(n954), .A2(n953), .ZN(n965) );
  NOR2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n963) );
  XOR2_X1 U1058 ( .A(G2090), .B(G162), .Z(n959) );
  NOR2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1060 ( .A(n961), .B(KEYINPUT51), .ZN(n962) );
  NOR2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n972) );
  XOR2_X1 U1063 ( .A(G164), .B(G2078), .Z(n968) );
  XNOR2_X1 U1064 ( .A(G2072), .B(n966), .ZN(n967) );
  NOR2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(KEYINPUT125), .B(n969), .ZN(n970) );
  XNOR2_X1 U1067 ( .A(KEYINPUT50), .B(n970), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(KEYINPUT52), .B(n973), .ZN(n974) );
  INV_X1 U1070 ( .A(KEYINPUT55), .ZN(n994) );
  NAND2_X1 U1071 ( .A1(n974), .A2(n994), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n975), .A2(G29), .ZN(n1052) );
  XNOR2_X1 U1073 ( .A(G2090), .B(G35), .ZN(n988) );
  XOR2_X1 U1074 ( .A(G2067), .B(G26), .Z(n976) );
  NAND2_X1 U1075 ( .A1(n976), .A2(G28), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(G1991), .B(G25), .ZN(n978) );
  XNOR2_X1 U1077 ( .A(G2072), .B(G33), .ZN(n977) );
  NOR2_X1 U1078 ( .A1(n978), .A2(n977), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(n979), .B(G27), .ZN(n981) );
  XNOR2_X1 U1080 ( .A(G1996), .B(G32), .ZN(n980) );
  NOR2_X1 U1081 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1082 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1083 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1084 ( .A(KEYINPUT53), .B(n986), .ZN(n987) );
  NOR2_X1 U1085 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1086 ( .A(n989), .B(KEYINPUT126), .ZN(n992) );
  XOR2_X1 U1087 ( .A(G2084), .B(G34), .Z(n990) );
  XNOR2_X1 U1088 ( .A(KEYINPUT54), .B(n990), .ZN(n991) );
  NAND2_X1 U1089 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1090 ( .A(n994), .B(n993), .ZN(n996) );
  INV_X1 U1091 ( .A(G29), .ZN(n995) );
  NAND2_X1 U1092 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1093 ( .A1(G11), .A2(n997), .ZN(n1050) );
  INV_X1 U1094 ( .A(G16), .ZN(n1046) );
  XNOR2_X1 U1095 ( .A(KEYINPUT56), .B(KEYINPUT127), .ZN(n998) );
  XNOR2_X1 U1096 ( .A(n1046), .B(n998), .ZN(n1022) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G168), .ZN(n1000) );
  NAND2_X1 U1098 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1099 ( .A(n1001), .B(KEYINPUT57), .ZN(n1020) );
  NAND2_X1 U1100 ( .A1(n1003), .A2(n1002), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(G301), .B(G1961), .ZN(n1006) );
  XNOR2_X1 U1102 ( .A(n1004), .B(G1341), .ZN(n1005) );
  NOR2_X1 U1103 ( .A1(n1006), .A2(n1005), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(n1007), .B(G1956), .ZN(n1009) );
  NAND2_X1 U1105 ( .A1(G1971), .A2(G303), .ZN(n1008) );
  NAND2_X1 U1106 ( .A1(n1009), .A2(n1008), .ZN(n1014) );
  XNOR2_X1 U1107 ( .A(G1348), .B(n1010), .ZN(n1012) );
  NAND2_X1 U1108 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1109 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1110 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1111 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1112 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1113 ( .A1(n1022), .A2(n1021), .ZN(n1048) );
  XNOR2_X1 U1114 ( .A(G5), .B(n1023), .ZN(n1036) );
  XNOR2_X1 U1115 ( .A(G20), .B(n1024), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(G1341), .B(G19), .ZN(n1026) );
  XNOR2_X1 U1117 ( .A(G1981), .B(G6), .ZN(n1025) );
  NOR2_X1 U1118 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1119 ( .A1(n1028), .A2(n1027), .ZN(n1031) );
  XOR2_X1 U1120 ( .A(KEYINPUT59), .B(G1348), .Z(n1029) );
  XNOR2_X1 U1121 ( .A(G4), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1122 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1123 ( .A(KEYINPUT60), .B(n1032), .Z(n1034) );
  XNOR2_X1 U1124 ( .A(G1966), .B(G21), .ZN(n1033) );
  NOR2_X1 U1125 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1126 ( .A1(n1036), .A2(n1035), .ZN(n1043) );
  XNOR2_X1 U1127 ( .A(G1971), .B(G22), .ZN(n1038) );
  XNOR2_X1 U1128 ( .A(G23), .B(G1976), .ZN(n1037) );
  NOR2_X1 U1129 ( .A1(n1038), .A2(n1037), .ZN(n1040) );
  XOR2_X1 U1130 ( .A(G1986), .B(G24), .Z(n1039) );
  NAND2_X1 U1131 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1132 ( .A(KEYINPUT58), .B(n1041), .ZN(n1042) );
  NOR2_X1 U1133 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  XNOR2_X1 U1134 ( .A(KEYINPUT61), .B(n1044), .ZN(n1045) );
  NAND2_X1 U1135 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  NAND2_X1 U1136 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
  NOR2_X1 U1137 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  NAND2_X1 U1138 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
  XOR2_X1 U1139 ( .A(KEYINPUT62), .B(n1053), .Z(G311) );
  INV_X1 U1140 ( .A(G311), .ZN(G150) );
endmodule

