//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934;
  XOR2_X1   g000(.A(KEYINPUT91), .B(G29gat), .Z(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G36gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT92), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT92), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n202), .A2(new_n205), .A3(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(KEYINPUT93), .B(G43gat), .Z(new_n208));
  INV_X1    g007(.A(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n209), .A2(G43gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT15), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n207), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT89), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT15), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n217), .B1(new_n214), .B2(new_n215), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT14), .ZN(new_n220));
  INV_X1    g019(.A(G29gat), .ZN(new_n221));
  INV_X1    g020(.A(G36gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n216), .A2(new_n218), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n219), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT90), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(new_n206), .A3(new_n204), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n216), .A2(new_n218), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n213), .A2(new_n224), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(G1gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G1gat), .B2(new_n230), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(G8gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT94), .B1(new_n229), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n227), .A2(new_n228), .ZN(new_n237));
  INV_X1    g036(.A(new_n212), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n238), .A2(new_n224), .A3(new_n206), .A4(new_n204), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT94), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(new_n234), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT17), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n229), .A2(KEYINPUT17), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(new_n235), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G229gat), .A2(G233gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT18), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n229), .A2(new_n235), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n229), .A2(new_n235), .A3(KEYINPUT94), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n241), .B1(new_n240), .B2(new_n234), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n249), .B(KEYINPUT13), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n243), .A2(new_n247), .A3(KEYINPUT18), .A4(new_n249), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n261));
  XNOR2_X1  g060(.A(G113gat), .B(G141gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(G169gat), .B(G197gat), .Z(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT12), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n252), .A2(new_n259), .A3(new_n260), .A4(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n259), .A2(new_n260), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT95), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT95), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n252), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n266), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n272), .A2(KEYINPUT96), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT96), .B1(new_n272), .B2(new_n273), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n267), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT36), .ZN(new_n278));
  XOR2_X1   g077(.A(KEYINPUT27), .B(G183gat), .Z(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G190gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G183gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(KEYINPUT70), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT27), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n286), .B(new_n287), .C1(KEYINPUT27), .C2(new_n284), .ZN(new_n288));
  NOR2_X1   g087(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n289));
  AOI22_X1  g088(.A1(KEYINPUT28), .A2(new_n282), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n290), .A2(KEYINPUT71), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(KEYINPUT71), .ZN(new_n293));
  INV_X1    g092(.A(G169gat), .ZN(new_n294));
  INV_X1    g093(.A(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n297));
  OR3_X1    g096(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT26), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT26), .B1(new_n296), .B2(new_n297), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n298), .B(new_n299), .C1(new_n294), .C2(new_n295), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n291), .A2(new_n292), .A3(new_n293), .A4(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT25), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n292), .B(KEYINPUT24), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  OR3_X1    g103(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT23), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT65), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n307), .A2(new_n308), .B1(G169gat), .B2(G176gat), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n306), .B(new_n309), .C1(new_n308), .C2(new_n307), .ZN(new_n310));
  AND2_X1   g109(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n311));
  NOR2_X1   g110(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n296), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(new_n313), .B(KEYINPUT67), .Z(new_n314));
  OAI21_X1  g113(.A(new_n302), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT68), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n285), .A2(G183gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n287), .A2(new_n317), .A3(new_n281), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n303), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n307), .B(KEYINPUT25), .C1(new_n294), .C2(new_n295), .ZN(new_n320));
  OR3_X1    g119(.A1(new_n314), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n315), .A2(KEYINPUT68), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n301), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT1), .ZN(new_n325));
  XOR2_X1   g124(.A(G113gat), .B(G120gat), .Z(new_n326));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n327));
  OAI211_X1 g126(.A(KEYINPUT74), .B(new_n325), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G127gat), .B(G134gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT74), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT73), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(new_n325), .A3(new_n326), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n324), .B(new_n334), .ZN(new_n335));
  AND2_X1   g134(.A1(G227gat), .A2(G233gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT32), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT33), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n335), .B2(new_n337), .ZN(new_n340));
  XNOR2_X1  g139(.A(G15gat), .B(G43gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G71gat), .B(G99gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  NAND3_X1  g142(.A1(new_n338), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n343), .ZN(new_n345));
  OAI221_X1 g144(.A(KEYINPUT32), .B1(new_n339), .B2(new_n345), .C1(new_n335), .C2(new_n337), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n335), .A2(new_n337), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT34), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n347), .B1(new_n350), .B2(KEYINPUT75), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n348), .B(KEYINPUT34), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n352), .A2(new_n344), .A3(new_n353), .A4(new_n346), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n278), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT77), .B1(new_n347), .B2(new_n352), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n347), .A2(new_n352), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n350), .A2(new_n344), .A3(new_n358), .A4(new_n346), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n361));
  AOI21_X1  g160(.A(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G197gat), .B(G204gat), .ZN(new_n363));
  INV_X1    g162(.A(G211gat), .ZN(new_n364));
  INV_X1    g163(.A(G218gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n363), .B1(KEYINPUT22), .B2(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(G211gat), .B(G218gat), .Z(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(G155gat), .B(G162gat), .Z(new_n371));
  XOR2_X1   g170(.A(G141gat), .B(G148gat), .Z(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(KEYINPUT79), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G155gat), .ZN(new_n374));
  INV_X1    g173(.A(G162gat), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT2), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n376), .B(new_n372), .C1(new_n371), .C2(KEYINPUT79), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n370), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n384), .B1(G228gat), .B2(G233gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n380), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n367), .A2(new_n368), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n383), .B1(new_n387), .B2(KEYINPUT83), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n388), .B1(new_n369), .B2(KEYINPUT83), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n386), .B1(new_n389), .B2(KEYINPUT3), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n370), .A2(new_n383), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n380), .B1(new_n392), .B2(new_n381), .ZN(new_n393));
  OAI211_X1 g192(.A(G228gat), .B(G233gat), .C1(new_n393), .C2(new_n384), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(G22gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(G78gat), .B(G106gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT31), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(G50gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n396), .B(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n324), .A2(G226gat), .A3(G233gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n324), .A2(new_n383), .B1(G226gat), .B2(G233gat), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT78), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n403), .A2(KEYINPUT78), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n369), .ZN(new_n407));
  XNOR2_X1  g206(.A(G8gat), .B(G36gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(G64gat), .B(G92gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n402), .A2(new_n403), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n370), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n407), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n370), .B1(new_n404), .B2(new_n405), .ZN(new_n415));
  INV_X1    g214(.A(new_n403), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n401), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(new_n369), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n410), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n414), .A2(KEYINPUT30), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n415), .A2(new_n418), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n422), .A3(new_n411), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT5), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n334), .B(KEYINPUT80), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n386), .A2(KEYINPUT3), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n382), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n380), .A2(new_n334), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT4), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G225gat), .A2(G233gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n427), .A2(new_n386), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n430), .ZN(new_n436));
  INV_X1    g235(.A(new_n433), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n426), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT5), .B1(new_n432), .B2(new_n433), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(KEYINPUT81), .B(KEYINPUT0), .Z(new_n442));
  XNOR2_X1  g241(.A(G1gat), .B(G29gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G57gat), .B(G85gat), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n444), .B(new_n445), .Z(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n425), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n446), .B1(new_n439), .B2(new_n440), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n441), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(new_n447), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n400), .B1(new_n424), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n362), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n454), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n414), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT38), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(new_n412), .B2(new_n370), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n417), .A2(KEYINPUT85), .A3(new_n369), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n461), .B(new_n462), .C1(new_n406), .C2(new_n369), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n463), .A2(KEYINPUT86), .A3(KEYINPUT37), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT86), .B1(new_n463), .B2(KEYINPUT37), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(new_n421), .B2(new_n468), .ZN(new_n469));
  NOR4_X1   g268(.A1(new_n415), .A2(new_n418), .A3(KEYINPUT87), .A4(KEYINPUT37), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n410), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n459), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n469), .A2(new_n470), .ZN(new_n473));
  OAI211_X1 g272(.A(KEYINPUT38), .B(new_n410), .C1(new_n421), .C2(new_n468), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n458), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n424), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n420), .A2(KEYINPUT84), .A3(new_n423), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n432), .A2(new_n433), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT39), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n437), .B2(new_n436), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n447), .B1(new_n481), .B2(new_n482), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n486), .A2(KEYINPUT40), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(KEYINPUT40), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n487), .A2(new_n448), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n479), .A2(new_n480), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n400), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n456), .B1(new_n477), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n479), .A2(new_n480), .ZN(new_n493));
  INV_X1    g292(.A(new_n400), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n360), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n457), .A2(KEYINPUT35), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n494), .B1(new_n351), .B2(new_n354), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(new_n424), .A3(new_n454), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n277), .B1(new_n492), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G230gat), .A2(G233gat), .ZN(new_n503));
  INV_X1    g302(.A(G57gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G64gat), .ZN(new_n505));
  INV_X1    g304(.A(G64gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(G57gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT9), .ZN(new_n508));
  NAND2_X1  g307(.A1(G71gat), .A2(G78gat), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n505), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT98), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g311(.A1(G71gat), .A2(G78gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n509), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(KEYINPUT97), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT97), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n510), .B2(new_n511), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n505), .A2(new_n507), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n509), .A2(new_n508), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n520), .A2(new_n509), .A3(new_n513), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n515), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G99gat), .A2(G106gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT101), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT101), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(G99gat), .A3(G106gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n526), .A3(KEYINPUT8), .ZN(new_n527));
  NOR2_X1   g326(.A1(G85gat), .A2(G92gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G99gat), .B(G106gat), .ZN(new_n532));
  NAND4_X1  g331(.A1(KEYINPUT100), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n527), .A2(new_n531), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT102), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n529), .A2(new_n530), .ZN(new_n536));
  INV_X1    g335(.A(G85gat), .ZN(new_n537));
  INV_X1    g336(.A(G92gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n536), .A2(new_n533), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT102), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n540), .A2(new_n541), .A3(new_n532), .A4(new_n527), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n532), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n524), .A2(new_n526), .A3(KEYINPUT8), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n536), .A2(new_n533), .A3(new_n539), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT103), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n527), .A2(new_n533), .A3(new_n531), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(KEYINPUT103), .A3(new_n544), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n522), .B1(new_n543), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n547), .A2(new_n534), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n522), .A2(new_n554), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n553), .A2(new_n555), .A3(KEYINPUT10), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n522), .A2(KEYINPUT10), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT104), .ZN(new_n558));
  AOI211_X1 g357(.A(new_n548), .B(new_n532), .C1(new_n540), .C2(new_n527), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT103), .B1(new_n550), .B2(new_n544), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n535), .A2(new_n542), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n543), .A2(new_n552), .A3(KEYINPUT104), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n557), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n503), .B1(new_n556), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT105), .ZN(new_n567));
  INV_X1    g366(.A(new_n503), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n568), .B1(new_n553), .B2(new_n555), .ZN(new_n569));
  INV_X1    g368(.A(new_n557), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n561), .A2(new_n558), .A3(new_n562), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT104), .B1(new_n543), .B2(new_n552), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n522), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(new_n561), .B2(new_n562), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT10), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n522), .A2(new_n554), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT105), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n503), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n567), .A2(new_n569), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G120gat), .B(G148gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n586), .A2(KEYINPUT106), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT106), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n588), .B1(new_n582), .B2(new_n585), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n585), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n566), .A2(new_n591), .A3(new_n569), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT107), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(KEYINPUT107), .B(new_n592), .C1(new_n587), .C2(new_n589), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT21), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n235), .B1(new_n598), .B2(new_n574), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT99), .ZN(new_n600));
  AND2_X1   g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n574), .A2(new_n598), .ZN(new_n603));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n602), .B(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G183gat), .B(G211gat), .Z(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n606), .B(new_n609), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n245), .A2(new_n246), .A3(new_n563), .A4(new_n564), .ZN(new_n611));
  NAND3_X1  g410(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n240), .B1(new_n571), .B2(new_n572), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G134gat), .B(G162gat), .Z(new_n615));
  AND2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  XNOR2_X1  g416(.A(G190gat), .B(G218gat), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n616), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n614), .A2(new_n615), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n614), .A2(new_n615), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n620), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n597), .A2(new_n610), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n502), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n457), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G1gat), .ZN(G1324gat));
  INV_X1    g430(.A(new_n493), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT16), .B(G8gat), .Z(new_n633));
  NAND3_X1  g432(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n634), .A2(KEYINPUT42), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT42), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n629), .A2(new_n632), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n637), .B2(G8gat), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n635), .B1(new_n634), .B2(new_n638), .ZN(G1325gat));
  INV_X1    g438(.A(G15gat), .ZN(new_n640));
  INV_X1    g439(.A(new_n362), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n628), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n360), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n629), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n642), .B1(new_n640), .B2(new_n644), .ZN(G1326gat));
  NOR2_X1   g444(.A1(new_n628), .A2(new_n400), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT43), .B(G22gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1327gat));
  NAND2_X1  g447(.A1(new_n501), .A2(KEYINPUT109), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT109), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n497), .A2(new_n650), .A3(new_n500), .ZN(new_n651));
  OAI221_X1 g450(.A(new_n410), .B1(new_n469), .B2(new_n470), .C1(new_n464), .C2(new_n465), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n475), .B1(new_n652), .B2(new_n459), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n400), .B(new_n490), .C1(new_n653), .C2(new_n458), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n649), .A2(new_n651), .B1(new_n654), .B2(new_n456), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT110), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(new_n622), .B2(new_n625), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n624), .A2(new_n620), .A3(new_n623), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n621), .B1(new_n616), .B2(new_n617), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT110), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n626), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n665), .B1(new_n492), .B2(new_n501), .ZN(new_n666));
  OAI22_X1  g465(.A1(new_n655), .A2(new_n664), .B1(new_n666), .B2(new_n663), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n667), .A2(new_n610), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n597), .A2(new_n277), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n202), .B1(new_n670), .B2(new_n454), .ZN(new_n671));
  INV_X1    g470(.A(new_n610), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n665), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT107), .B1(new_n590), .B2(new_n592), .ZN(new_n674));
  INV_X1    g473(.A(new_n596), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT108), .Z(new_n678));
  NAND2_X1  g477(.A1(new_n502), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n679), .A2(new_n454), .A3(new_n202), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT45), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n671), .A2(new_n681), .ZN(G1328gat));
  OAI21_X1  g481(.A(G36gat), .B1(new_n670), .B2(new_n493), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n632), .A2(new_n222), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT46), .B1(new_n679), .B2(new_n684), .ZN(new_n685));
  OR3_X1    g484(.A1(new_n679), .A2(KEYINPUT46), .A3(new_n684), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(G1329gat));
  NOR3_X1   g486(.A1(new_n679), .A2(new_n360), .A3(new_n208), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n667), .A2(new_n362), .A3(new_n610), .A4(new_n669), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n689), .B2(new_n208), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n690), .B(new_n692), .ZN(G1330gat));
  NAND4_X1  g492(.A1(new_n667), .A2(new_n494), .A3(new_n610), .A4(new_n669), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G50gat), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n502), .A2(new_n209), .A3(new_n494), .A4(new_n678), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n695), .A2(KEYINPUT48), .A3(new_n696), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1331gat));
  NAND2_X1  g500(.A1(new_n649), .A2(new_n651), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n492), .ZN(new_n703));
  NOR4_X1   g502(.A1(new_n676), .A2(new_n276), .A3(new_n610), .A4(new_n626), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n454), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(new_n504), .ZN(G1332gat));
  AND2_X1   g506(.A1(new_n703), .A2(new_n704), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n493), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT112), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n711), .B(new_n712), .Z(G1333gat));
  NAND3_X1  g512(.A1(new_n708), .A2(G71gat), .A3(new_n362), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n705), .A2(new_n360), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(G71gat), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g516(.A1(new_n708), .A2(new_n494), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g518(.A1(new_n676), .A2(new_n276), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n668), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G85gat), .B1(new_n721), .B2(new_n454), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n703), .A2(KEYINPUT51), .A3(new_n277), .A4(new_n673), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT51), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n673), .A2(new_n277), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n655), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT113), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(KEYINPUT113), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n597), .A2(new_n457), .A3(new_n537), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n722), .B1(new_n731), .B2(new_n732), .ZN(G1336gat));
  NAND3_X1  g532(.A1(new_n632), .A2(new_n538), .A3(new_n597), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n729), .B2(new_n730), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n667), .A2(new_n632), .A3(new_n610), .A4(new_n720), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G92gat), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n734), .B1(new_n723), .B2(new_n726), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(G92gat), .B2(new_n736), .ZN(new_n741));
  OAI22_X1  g540(.A1(new_n735), .A2(new_n739), .B1(new_n741), .B2(new_n738), .ZN(G1337gat));
  OAI21_X1  g541(.A(G99gat), .B1(new_n721), .B2(new_n641), .ZN(new_n743));
  OR3_X1    g542(.A1(new_n676), .A2(new_n360), .A3(G99gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n731), .B2(new_n744), .ZN(G1338gat));
  OR3_X1    g544(.A1(new_n676), .A2(G106gat), .A3(new_n400), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(new_n729), .B2(new_n730), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n667), .A2(new_n494), .A3(new_n610), .A4(new_n720), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G106gat), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n746), .B1(new_n723), .B2(new_n726), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(G106gat), .B2(new_n748), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n747), .A2(new_n751), .B1(new_n753), .B2(new_n750), .ZN(G1339gat));
  NAND2_X1  g553(.A1(new_n627), .A2(new_n277), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n573), .A2(new_n568), .A3(new_n578), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n566), .A2(KEYINPUT54), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT54), .B1(new_n567), .B2(new_n581), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT114), .B1(new_n759), .B2(new_n591), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n580), .B1(new_n579), .B2(new_n503), .ZN(new_n762));
  AOI211_X1 g561(.A(KEYINPUT105), .B(new_n568), .C1(new_n573), .C2(new_n578), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n764), .A2(new_n765), .A3(new_n585), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n756), .B(new_n758), .C1(new_n760), .C2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n592), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT115), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n256), .A2(new_n258), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(KEYINPUT116), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n243), .A2(KEYINPUT116), .A3(new_n253), .A4(new_n257), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n248), .B2(new_n249), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n265), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n267), .A2(new_n774), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n775), .A2(new_n660), .A3(new_n657), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n766), .ZN(new_n777));
  INV_X1    g576(.A(new_n758), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(KEYINPUT55), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(new_n780), .A3(new_n592), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n777), .A2(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n756), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n769), .A2(new_n776), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT117), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n779), .A2(new_n592), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n787), .A2(KEYINPUT115), .B1(new_n756), .B2(new_n782), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n788), .A2(KEYINPUT117), .A3(new_n781), .A4(new_n776), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n769), .A2(new_n276), .A3(new_n781), .A4(new_n783), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n775), .B1(new_n674), .B2(new_n675), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n786), .A2(new_n789), .B1(new_n792), .B2(new_n661), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n755), .B1(new_n793), .B2(new_n672), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(new_n498), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n632), .A2(new_n454), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OR3_X1    g596(.A1(new_n797), .A2(G113gat), .A3(new_n277), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n493), .A2(new_n495), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n786), .A2(new_n789), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n792), .A2(new_n661), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n672), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n755), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n457), .B(new_n799), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n794), .A2(KEYINPUT118), .A3(new_n457), .A4(new_n799), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n276), .A3(new_n807), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n808), .A2(KEYINPUT119), .A3(G113gat), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT119), .B1(new_n808), .B2(G113gat), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n798), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT120), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT120), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n813), .B(new_n798), .C1(new_n809), .C2(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1340gat));
  NAND2_X1  g614(.A1(new_n806), .A2(new_n807), .ZN(new_n816));
  OAI21_X1  g615(.A(G120gat), .B1(new_n816), .B2(new_n676), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n676), .A2(G120gat), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n797), .B2(new_n818), .ZN(G1341gat));
  NAND4_X1  g618(.A1(new_n806), .A2(G127gat), .A3(new_n672), .A4(new_n807), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n797), .ZN(new_n823));
  AOI21_X1  g622(.A(G127gat), .B1(new_n823), .B2(new_n672), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n820), .A2(new_n821), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(G1342gat));
  NOR3_X1   g625(.A1(new_n797), .A2(G134gat), .A3(new_n665), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT56), .ZN(new_n828));
  OAI21_X1  g627(.A(G134gat), .B1(new_n816), .B2(new_n665), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1343gat));
  NOR2_X1   g629(.A1(new_n802), .A2(new_n803), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n400), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n791), .ZN(new_n835));
  AND4_X1   g634(.A1(new_n276), .A2(new_n592), .A3(new_n779), .A4(new_n783), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n665), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n672), .B1(new_n800), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n494), .B1(new_n838), .B2(new_n803), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT57), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n641), .A2(new_n493), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n454), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n834), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G141gat), .B1(new_n843), .B2(new_n277), .ZN(new_n844));
  XNOR2_X1  g643(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n831), .B2(new_n454), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n794), .A2(KEYINPUT122), .A3(new_n457), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n841), .A2(new_n400), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(G141gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n852), .A3(new_n276), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n844), .A2(new_n845), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n845), .B1(new_n844), .B2(new_n853), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(G1344gat));
  NOR2_X1   g655(.A1(new_n676), .A2(G148gat), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n850), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT124), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n859), .B(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT57), .B1(new_n831), .B2(new_n400), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n788), .A2(new_n626), .A3(new_n781), .A4(new_n775), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n672), .B1(new_n837), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n833), .B(new_n494), .C1(new_n865), .C2(new_n803), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n863), .A2(new_n866), .A3(new_n597), .A4(new_n842), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(KEYINPUT125), .ZN(new_n868));
  INV_X1    g667(.A(G148gat), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n867), .B2(KEYINPUT125), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n862), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n862), .A2(G148gat), .ZN(new_n872));
  INV_X1    g671(.A(new_n843), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n597), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n861), .B1(new_n871), .B2(new_n874), .ZN(G1345gat));
  NOR3_X1   g674(.A1(new_n843), .A2(new_n374), .A3(new_n610), .ZN(new_n876));
  AOI21_X1  g675(.A(G155gat), .B1(new_n851), .B2(new_n672), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(G1346gat));
  NOR3_X1   g677(.A1(new_n843), .A2(new_n375), .A3(new_n661), .ZN(new_n879));
  AOI21_X1  g678(.A(G162gat), .B1(new_n851), .B2(new_n626), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(G1347gat));
  NOR2_X1   g680(.A1(new_n493), .A2(new_n457), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n795), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n294), .A3(new_n276), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n882), .A2(new_n643), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n494), .B1(new_n886), .B2(KEYINPUT126), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n882), .A2(new_n888), .A3(new_n643), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n887), .A2(new_n794), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n276), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n885), .B1(new_n294), .B2(new_n892), .ZN(G1348gat));
  AOI21_X1  g692(.A(G176gat), .B1(new_n884), .B2(new_n597), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n676), .A2(new_n295), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n890), .B2(new_n895), .ZN(G1349gat));
  NAND2_X1  g695(.A1(new_n890), .A2(new_n672), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n287), .A2(new_n317), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n672), .A2(new_n280), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n883), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n281), .A3(new_n662), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n890), .A2(new_n626), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(G190gat), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT61), .B(new_n281), .C1(new_n890), .C2(new_n626), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT127), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n910), .B(new_n903), .C1(new_n906), .C2(new_n907), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1351gat));
  AND2_X1   g711(.A1(new_n863), .A2(new_n866), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n882), .A2(new_n641), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n276), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G197gat), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n832), .A2(new_n915), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n277), .A2(G197gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(G1352gat));
  NOR3_X1   g720(.A1(new_n919), .A2(G204gat), .A3(new_n676), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT62), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n913), .A2(new_n597), .A3(new_n915), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G204gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1353gat));
  INV_X1    g725(.A(new_n919), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n364), .A3(new_n672), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n913), .A2(new_n672), .A3(new_n915), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT63), .B1(new_n929), .B2(G211gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1354gat));
  AOI21_X1  g731(.A(G218gat), .B1(new_n927), .B2(new_n662), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n665), .A2(new_n365), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n916), .B2(new_n934), .ZN(G1355gat));
endmodule


