

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594;

  INV_X1 U324 ( .A(KEYINPUT107), .ZN(n495) );
  INV_X1 U325 ( .A(n395), .ZN(n396) );
  XOR2_X1 U326 ( .A(G211GAT), .B(KEYINPUT21), .Z(n292) );
  XOR2_X1 U327 ( .A(KEYINPUT40), .B(n512), .Z(n293) );
  XNOR2_X1 U328 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U329 ( .A(n461), .B(KEYINPUT27), .ZN(n462) );
  XNOR2_X1 U330 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n388) );
  XNOR2_X1 U331 ( .A(n418), .B(n417), .ZN(n421) );
  XNOR2_X1 U332 ( .A(n463), .B(n462), .ZN(n474) );
  XNOR2_X1 U333 ( .A(n419), .B(n388), .ZN(n392) );
  XNOR2_X1 U334 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U335 ( .A(n399), .B(n398), .ZN(n401) );
  INV_X1 U336 ( .A(G190GAT), .ZN(n456) );
  XOR2_X1 U337 ( .A(KEYINPUT78), .B(n562), .Z(n546) );
  XNOR2_X1 U338 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U339 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(G176GAT), .B(G183GAT), .Z(n295) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n294) );
  XNOR2_X1 U342 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U343 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n297) );
  XNOR2_X1 U344 ( .A(KEYINPUT85), .B(KEYINPUT17), .ZN(n296) );
  XNOR2_X1 U345 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n461) );
  XOR2_X1 U347 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n301) );
  XNOR2_X1 U348 ( .A(KEYINPUT86), .B(KEYINPUT20), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U350 ( .A(n461), .B(n302), .Z(n312) );
  XNOR2_X1 U351 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n303), .B(KEYINPUT81), .ZN(n437) );
  XOR2_X1 U353 ( .A(KEYINPUT64), .B(n437), .Z(n305) );
  NAND2_X1 U354 ( .A1(G227GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U356 ( .A(G43GAT), .B(G134GAT), .Z(n389) );
  XNOR2_X1 U357 ( .A(n306), .B(n389), .ZN(n310) );
  XOR2_X1 U358 ( .A(G99GAT), .B(G190GAT), .Z(n308) );
  XOR2_X1 U359 ( .A(G120GAT), .B(G71GAT), .Z(n379) );
  XOR2_X1 U360 ( .A(G15GAT), .B(G127GAT), .Z(n329) );
  XNOR2_X1 U361 ( .A(n379), .B(n329), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U364 ( .A(n312), .B(n311), .Z(n537) );
  INV_X1 U365 ( .A(n537), .ZN(n511) );
  XOR2_X1 U366 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n314) );
  XNOR2_X1 U367 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U369 ( .A(KEYINPUT3), .B(n315), .Z(n450) );
  XOR2_X1 U370 ( .A(G106GAT), .B(G218GAT), .Z(n317) );
  XOR2_X1 U371 ( .A(G50GAT), .B(G162GAT), .Z(n395) );
  XOR2_X1 U372 ( .A(G148GAT), .B(G78GAT), .Z(n371) );
  XNOR2_X1 U373 ( .A(n395), .B(n371), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n322) );
  XNOR2_X1 U375 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n292), .B(n318), .ZN(n413) );
  XOR2_X1 U377 ( .A(G204GAT), .B(n413), .Z(n320) );
  NAND2_X1 U378 ( .A1(G228GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U380 ( .A(n322), .B(n321), .Z(n327) );
  XOR2_X1 U381 ( .A(G141GAT), .B(G22GAT), .Z(n352) );
  XOR2_X1 U382 ( .A(KEYINPUT91), .B(KEYINPUT23), .Z(n324) );
  XNOR2_X1 U383 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n352), .B(n325), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n450), .B(n328), .ZN(n472) );
  XOR2_X1 U388 ( .A(G57GAT), .B(KEYINPUT13), .Z(n366) );
  XOR2_X1 U389 ( .A(G8GAT), .B(KEYINPUT79), .Z(n414) );
  XOR2_X1 U390 ( .A(n366), .B(n414), .Z(n331) );
  XOR2_X1 U391 ( .A(KEYINPUT70), .B(G1GAT), .Z(n351) );
  XNOR2_X1 U392 ( .A(n351), .B(n329), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n331), .B(n330), .ZN(n344) );
  XOR2_X1 U394 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n333) );
  NAND2_X1 U395 ( .A1(G231GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U396 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U397 ( .A(n334), .B(KEYINPUT80), .Z(n342) );
  XOR2_X1 U398 ( .A(G78GAT), .B(G211GAT), .Z(n336) );
  XNOR2_X1 U399 ( .A(G22GAT), .B(G155GAT), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U401 ( .A(KEYINPUT14), .B(G64GAT), .Z(n338) );
  XNOR2_X1 U402 ( .A(G183GAT), .B(G71GAT), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U406 ( .A(n344), .B(n343), .ZN(n559) );
  INV_X1 U407 ( .A(n559), .ZN(n587) );
  XOR2_X1 U408 ( .A(G8GAT), .B(G113GAT), .Z(n346) );
  XNOR2_X1 U409 ( .A(G169GAT), .B(G15GAT), .ZN(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U411 ( .A(KEYINPUT71), .B(KEYINPUT68), .Z(n348) );
  XNOR2_X1 U412 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n363) );
  XOR2_X1 U415 ( .A(G197GAT), .B(G43GAT), .Z(n354) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U418 ( .A(n355), .B(G50GAT), .Z(n361) );
  XNOR2_X1 U419 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n356), .B(KEYINPUT7), .ZN(n394) );
  XOR2_X1 U421 ( .A(n394), .B(KEYINPUT69), .Z(n358) );
  NAND2_X1 U422 ( .A1(G229GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n359), .B(G36GAT), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U426 ( .A(n363), .B(n362), .Z(n552) );
  XOR2_X1 U427 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n365) );
  XNOR2_X1 U428 ( .A(KEYINPUT76), .B(KEYINPUT32), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n383) );
  XOR2_X1 U430 ( .A(G204GAT), .B(G64GAT), .Z(n426) );
  XOR2_X1 U431 ( .A(n426), .B(n366), .Z(n368) );
  XNOR2_X1 U432 ( .A(G176GAT), .B(G92GAT), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n368), .B(n367), .ZN(n375) );
  XOR2_X1 U434 ( .A(KEYINPUT74), .B(G85GAT), .Z(n370) );
  XNOR2_X1 U435 ( .A(G99GAT), .B(G106GAT), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(n369), .ZN(n393) );
  XOR2_X1 U437 ( .A(n393), .B(n371), .Z(n373) );
  NAND2_X1 U438 ( .A1(G230GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U439 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U440 ( .A(n375), .B(n374), .Z(n381) );
  XOR2_X1 U441 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n377) );
  XNOR2_X1 U442 ( .A(KEYINPUT73), .B(KEYINPUT77), .ZN(n376) );
  XNOR2_X1 U443 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U444 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n581) );
  XOR2_X1 U447 ( .A(n581), .B(KEYINPUT41), .Z(n554) );
  NOR2_X1 U448 ( .A1(n552), .A2(n554), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n384), .B(KEYINPUT46), .ZN(n385) );
  NOR2_X1 U450 ( .A1(n587), .A2(n385), .ZN(n402) );
  XOR2_X1 U451 ( .A(G92GAT), .B(G218GAT), .Z(n387) );
  XNOR2_X1 U452 ( .A(G36GAT), .B(G190GAT), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n419) );
  XNOR2_X1 U454 ( .A(n389), .B(KEYINPUT65), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n390), .B(KEYINPUT11), .ZN(n391) );
  XOR2_X1 U456 ( .A(n392), .B(n391), .Z(n399) );
  XNOR2_X1 U457 ( .A(n394), .B(n393), .ZN(n397) );
  NAND2_X1 U458 ( .A1(G232GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n562) );
  NAND2_X1 U460 ( .A1(n402), .A2(n562), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n403), .B(KEYINPUT47), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n404), .B(KEYINPUT114), .ZN(n411) );
  XNOR2_X1 U463 ( .A(KEYINPUT36), .B(n546), .ZN(n590) );
  NAND2_X1 U464 ( .A1(n587), .A2(n590), .ZN(n407) );
  XNOR2_X1 U465 ( .A(KEYINPUT115), .B(KEYINPUT45), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n405), .B(KEYINPUT66), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n408) );
  NAND2_X1 U468 ( .A1(n408), .A2(n581), .ZN(n409) );
  INV_X1 U469 ( .A(n552), .ZN(n576) );
  NOR2_X1 U470 ( .A1(n409), .A2(n576), .ZN(n410) );
  NOR2_X1 U471 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n412), .B(KEYINPUT48), .ZN(n535) );
  XOR2_X1 U473 ( .A(n414), .B(n413), .Z(n418) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n416) );
  INV_X1 U475 ( .A(KEYINPUT98), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n419), .B(KEYINPUT96), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n423) );
  INV_X1 U478 ( .A(KEYINPUT99), .ZN(n422) );
  NAND2_X1 U479 ( .A1(n423), .A2(n422), .ZN(n425) );
  OR2_X1 U480 ( .A1(n423), .A2(n422), .ZN(n424) );
  NAND2_X1 U481 ( .A1(n425), .A2(n424), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n426), .B(KEYINPUT97), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n463) );
  XNOR2_X1 U484 ( .A(n461), .B(n463), .ZN(n507) );
  INV_X1 U485 ( .A(n507), .ZN(n527) );
  XNOR2_X1 U486 ( .A(KEYINPUT119), .B(n527), .ZN(n429) );
  NOR2_X1 U487 ( .A1(n535), .A2(n429), .ZN(n430) );
  XNOR2_X1 U488 ( .A(KEYINPUT54), .B(n430), .ZN(n453) );
  XOR2_X1 U489 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n432) );
  XNOR2_X1 U490 ( .A(KEYINPUT92), .B(KEYINPUT95), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U492 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n434) );
  XNOR2_X1 U493 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U495 ( .A(n436), .B(n435), .Z(n442) );
  XOR2_X1 U496 ( .A(G85GAT), .B(n437), .Z(n439) );
  NAND2_X1 U497 ( .A1(G225GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U499 ( .A(G29GAT), .B(n440), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U501 ( .A(G148GAT), .B(G162GAT), .Z(n444) );
  XNOR2_X1 U502 ( .A(G141GAT), .B(G134GAT), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U504 ( .A(n446), .B(n445), .Z(n452) );
  XOR2_X1 U505 ( .A(G57GAT), .B(G127GAT), .Z(n448) );
  XNOR2_X1 U506 ( .A(G1GAT), .B(G120GAT), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U509 ( .A(n452), .B(n451), .Z(n525) );
  INV_X1 U510 ( .A(n525), .ZN(n503) );
  NAND2_X1 U511 ( .A1(n453), .A2(n503), .ZN(n574) );
  NOR2_X1 U512 ( .A1(n472), .A2(n574), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n454), .B(KEYINPUT55), .ZN(n455) );
  NOR2_X2 U514 ( .A1(n511), .A2(n455), .ZN(n571) );
  NAND2_X1 U515 ( .A1(n571), .A2(n546), .ZN(n459) );
  XOR2_X1 U516 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n457) );
  NOR2_X1 U517 ( .A1(n546), .A2(n559), .ZN(n460) );
  XNOR2_X1 U518 ( .A(n460), .B(KEYINPUT16), .ZN(n481) );
  NOR2_X1 U519 ( .A1(n503), .A2(n474), .ZN(n465) );
  INV_X1 U520 ( .A(KEYINPUT100), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n465), .B(n464), .ZN(n536) );
  XOR2_X1 U522 ( .A(KEYINPUT28), .B(KEYINPUT67), .Z(n466) );
  XOR2_X1 U523 ( .A(n472), .B(n466), .Z(n513) );
  INV_X1 U524 ( .A(n513), .ZN(n540) );
  NOR2_X1 U525 ( .A1(n536), .A2(n540), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n467), .B(KEYINPUT101), .ZN(n469) );
  XOR2_X1 U527 ( .A(n537), .B(KEYINPUT87), .Z(n468) );
  NOR2_X1 U528 ( .A1(n469), .A2(n468), .ZN(n479) );
  NOR2_X1 U529 ( .A1(n511), .A2(n507), .ZN(n470) );
  NOR2_X1 U530 ( .A1(n472), .A2(n470), .ZN(n471) );
  XOR2_X1 U531 ( .A(KEYINPUT25), .B(n471), .Z(n476) );
  NAND2_X1 U532 ( .A1(n472), .A2(n511), .ZN(n473) );
  XOR2_X1 U533 ( .A(n473), .B(KEYINPUT26), .Z(n550) );
  INV_X1 U534 ( .A(n550), .ZN(n575) );
  NOR2_X1 U535 ( .A1(n575), .A2(n474), .ZN(n475) );
  NOR2_X1 U536 ( .A1(n476), .A2(n475), .ZN(n477) );
  NOR2_X1 U537 ( .A1(n525), .A2(n477), .ZN(n478) );
  NOR2_X1 U538 ( .A1(n479), .A2(n478), .ZN(n494) );
  INV_X1 U539 ( .A(n494), .ZN(n480) );
  NAND2_X1 U540 ( .A1(n481), .A2(n480), .ZN(n515) );
  NAND2_X1 U541 ( .A1(n576), .A2(n581), .ZN(n500) );
  NOR2_X1 U542 ( .A1(n515), .A2(n500), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n482), .B(KEYINPUT102), .ZN(n491) );
  NAND2_X1 U544 ( .A1(n491), .A2(n525), .ZN(n486) );
  XOR2_X1 U545 ( .A(KEYINPUT34), .B(KEYINPUT104), .Z(n484) );
  XNOR2_X1 U546 ( .A(G1GAT), .B(KEYINPUT103), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(G1324GAT) );
  NAND2_X1 U549 ( .A1(n491), .A2(n527), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n487), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT35), .B(KEYINPUT105), .Z(n489) );
  NAND2_X1 U552 ( .A1(n491), .A2(n537), .ZN(n488) );
  XNOR2_X1 U553 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U554 ( .A(G15GAT), .B(n490), .Z(G1326GAT) );
  NAND2_X1 U555 ( .A1(n491), .A2(n540), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n492), .B(KEYINPUT106), .ZN(n493) );
  XNOR2_X1 U557 ( .A(G22GAT), .B(n493), .ZN(G1327GAT) );
  XNOR2_X1 U558 ( .A(KEYINPUT39), .B(KEYINPUT110), .ZN(n505) );
  NOR2_X1 U559 ( .A1(n587), .A2(n494), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(n497) );
  NAND2_X1 U561 ( .A1(n497), .A2(n590), .ZN(n499) );
  XOR2_X1 U562 ( .A(KEYINPUT108), .B(KEYINPUT37), .Z(n498) );
  XNOR2_X1 U563 ( .A(n499), .B(n498), .ZN(n524) );
  NOR2_X1 U564 ( .A1(n524), .A2(n500), .ZN(n502) );
  XNOR2_X1 U565 ( .A(KEYINPUT38), .B(KEYINPUT109), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(n510) );
  NOR2_X1 U567 ( .A1(n503), .A2(n510), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U569 ( .A(G29GAT), .B(n506), .ZN(G1328GAT) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(KEYINPUT111), .ZN(n509) );
  NOR2_X1 U571 ( .A1(n507), .A2(n510), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1329GAT) );
  NOR2_X1 U573 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G43GAT), .B(n293), .ZN(G1330GAT) );
  NOR2_X1 U575 ( .A1(n510), .A2(n513), .ZN(n514) );
  XOR2_X1 U576 ( .A(G50GAT), .B(n514), .Z(G1331GAT) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n517) );
  INV_X1 U578 ( .A(n554), .ZN(n566) );
  NAND2_X1 U579 ( .A1(n566), .A2(n552), .ZN(n523) );
  NOR2_X1 U580 ( .A1(n523), .A2(n515), .ZN(n520) );
  NAND2_X1 U581 ( .A1(n520), .A2(n525), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1332GAT) );
  NAND2_X1 U583 ( .A1(n527), .A2(n520), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U585 ( .A1(n537), .A2(n520), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n519), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(G78GAT), .B(KEYINPUT43), .Z(n522) );
  NAND2_X1 U588 ( .A1(n520), .A2(n540), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(G1335GAT) );
  NOR2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n531) );
  NAND2_X1 U591 ( .A1(n531), .A2(n525), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(n526), .ZN(G1336GAT) );
  NAND2_X1 U593 ( .A1(n527), .A2(n531), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n531), .A2(n537), .ZN(n529) );
  XNOR2_X1 U596 ( .A(KEYINPUT112), .B(n529), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G99GAT), .B(n530), .ZN(G1338GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n533) );
  NAND2_X1 U599 ( .A1(n531), .A2(n540), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  NOR2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n551) );
  NAND2_X1 U603 ( .A1(n551), .A2(n537), .ZN(n538) );
  XNOR2_X1 U604 ( .A(KEYINPUT116), .B(n538), .ZN(n539) );
  NOR2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n576), .A2(n547), .ZN(n541) );
  XNOR2_X1 U607 ( .A(G113GAT), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U609 ( .A1(n547), .A2(n566), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  NAND2_X1 U611 ( .A1(n547), .A2(n587), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n544), .B(KEYINPUT50), .ZN(n545) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n561) );
  NOR2_X1 U618 ( .A1(n552), .A2(n561), .ZN(n553) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n553), .Z(G1344GAT) );
  NOR2_X1 U620 ( .A1(n561), .A2(n554), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n556) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n561), .ZN(n560) );
  XOR2_X1 U626 ( .A(G155GAT), .B(n560), .Z(G1346GAT) );
  NOR2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT118), .B(n563), .Z(n564) );
  XNOR2_X1 U629 ( .A(G162GAT), .B(n564), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n576), .A2(n571), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(n565), .ZN(G1348GAT) );
  XNOR2_X1 U632 ( .A(KEYINPUT57), .B(KEYINPUT120), .ZN(n570) );
  XOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT56), .Z(n568) );
  NAND2_X1 U634 ( .A1(n571), .A2(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  XOR2_X1 U637 ( .A(G183GAT), .B(KEYINPUT121), .Z(n573) );
  NAND2_X1 U638 ( .A1(n571), .A2(n587), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1350GAT) );
  XOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT60), .Z(n578) );
  NOR2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n591) );
  NAND2_X1 U642 ( .A1(n591), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n584) );
  INV_X1 U647 ( .A(n581), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n591), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n586) );
  XOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT124), .Z(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n591), .A2(n587), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(KEYINPUT126), .ZN(n589) );
  XNOR2_X1 U654 ( .A(G211GAT), .B(n589), .ZN(G1354GAT) );
  XOR2_X1 U655 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n593) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

