//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT65), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n212), .A2(new_n213), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n219), .A2(G13), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT64), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n221), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XOR2_X1   g0033(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G226), .B(G232), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT67), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XOR2_X1   g0047(.A(G50), .B(G58), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n224), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n252), .B1(new_n253), .B2(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G50), .ZN(new_n255));
  INV_X1    g0055(.A(G13), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n256), .A2(new_n225), .A3(G1), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n255), .B1(G50), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT68), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n225), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n259), .B1(new_n267), .B2(new_n252), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G222), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G223), .A2(G1698), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n279), .B(new_n280), .C1(G77), .C2(new_n275), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  OAI211_X1 g0084(.A(G1), .B(G13), .C1(new_n272), .C2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n285), .A3(G274), .ZN(new_n286));
  INV_X1    g0086(.A(G226), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n282), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n281), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(G200), .B2(new_n289), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n270), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT10), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n265), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(new_n201), .ZN(new_n298));
  INV_X1    g0098(.A(G77), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n262), .A2(new_n299), .B1(new_n225), .B2(G68), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n252), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT11), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n301), .A2(new_n302), .ZN(new_n304));
  OR3_X1    g0104(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT70), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT70), .B1(new_n303), .B2(new_n304), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n257), .A2(new_n203), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT12), .B1(new_n307), .B2(KEYINPUT71), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(KEYINPUT71), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n307), .A2(KEYINPUT71), .A3(KEYINPUT12), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n310), .A2(new_n311), .B1(G68), .B2(new_n254), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n305), .A2(new_n306), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT14), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(KEYINPUT72), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n287), .A2(new_n276), .ZN(new_n317));
  INV_X1    g0117(.A(G232), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G1698), .ZN(new_n319));
  AND2_X1   g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(KEYINPUT3), .A2(G33), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n317), .B(new_n319), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G97), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT69), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT69), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n322), .A2(new_n326), .A3(new_n323), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n280), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT13), .ZN(new_n329));
  INV_X1    g0129(.A(G238), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n286), .B1(new_n288), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n328), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n329), .B1(new_n328), .B2(new_n332), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n314), .B(new_n316), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n322), .A2(new_n326), .A3(new_n323), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n326), .B1(new_n322), .B2(new_n323), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n336), .A2(new_n337), .A3(new_n285), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT13), .B1(new_n338), .B2(new_n331), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n328), .A2(new_n329), .A3(new_n332), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(new_n340), .A3(G179), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n340), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n314), .B1(new_n343), .B2(new_n316), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n313), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n313), .B1(G200), .B2(new_n343), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n339), .A2(G190), .A3(new_n340), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G238), .A2(G1698), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n275), .B(new_n349), .C1(new_n318), .C2(G1698), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n280), .C1(G107), .C2(new_n275), .ZN(new_n351));
  INV_X1    g0151(.A(G244), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n351), .B(new_n286), .C1(new_n352), .C2(new_n288), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(G179), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n315), .B2(new_n353), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n258), .A2(G77), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(new_n254), .B2(G77), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT15), .B(G87), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n358), .A2(new_n262), .B1(new_n225), .B2(new_n299), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n260), .A2(new_n297), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n252), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n289), .A2(new_n315), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(G179), .B2(new_n289), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(new_n268), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n353), .A2(G200), .ZN(new_n368));
  INV_X1    g0168(.A(new_n362), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n368), .B(new_n369), .C1(new_n290), .C2(new_n353), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n363), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n296), .A2(new_n345), .A3(new_n348), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n261), .A2(new_n254), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n258), .B2(new_n261), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n273), .A2(new_n225), .A3(new_n274), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT73), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n273), .A2(KEYINPUT7), .A3(new_n225), .A4(new_n274), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n376), .A2(KEYINPUT73), .A3(new_n377), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(G68), .A3(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n202), .A2(new_n203), .ZN(new_n384));
  NOR2_X1   g0184(.A1(G58), .A2(G68), .ZN(new_n385));
  OAI21_X1  g0185(.A(G20), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n265), .A2(G159), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT16), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n320), .A2(new_n321), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT7), .B1(new_n391), .B2(new_n225), .ZN(new_n392));
  INV_X1    g0192(.A(new_n380), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(KEYINPUT16), .A3(new_n389), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n252), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n375), .B1(new_n390), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT74), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT74), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n375), .B(new_n399), .C1(new_n390), .C2(new_n396), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n287), .A2(G1698), .ZN(new_n401));
  OAI221_X1 g0201(.A(new_n401), .B1(G223), .B2(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT75), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT75), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(G33), .A3(G87), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n285), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT76), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT76), .ZN(new_n411));
  NOR2_X1   g0211(.A1(G223), .A2(G1698), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n287), .B2(G1698), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n407), .B1(new_n275), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n411), .B1(new_n414), .B2(new_n285), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n286), .B1(new_n288), .B2(new_n318), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(G179), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n409), .A2(new_n417), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n416), .A2(new_n418), .B1(new_n315), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n398), .A2(new_n400), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT18), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n398), .A2(new_n423), .A3(new_n400), .A4(new_n420), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n417), .A2(G190), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(new_n410), .A3(new_n415), .ZN(new_n426));
  INV_X1    g0226(.A(G200), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n409), .B2(new_n417), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n375), .C1(new_n390), .C2(new_n396), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT17), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n395), .A2(new_n252), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n383), .A2(new_n389), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT16), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n374), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n429), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n431), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n422), .A2(new_n424), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n372), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n257), .A2(new_n210), .ZN(new_n443));
  INV_X1    g0243(.A(new_n252), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n258), .B(new_n444), .C1(G1), .C2(new_n272), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n445), .B2(new_n210), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n381), .A2(G107), .A3(new_n382), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT77), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT77), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n381), .A2(new_n449), .A3(G107), .A4(new_n382), .ZN(new_n450));
  INV_X1    g0250(.A(G107), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(KEYINPUT6), .A3(G97), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n210), .A2(new_n451), .ZN(new_n453));
  NOR2_X1   g0253(.A1(G97), .A2(G107), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n452), .B1(new_n455), .B2(KEYINPUT6), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(G20), .B1(G77), .B2(new_n265), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n448), .A2(new_n450), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n446), .B1(new_n458), .B2(new_n252), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n253), .B(G45), .C1(new_n284), .C2(KEYINPUT5), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT5), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G41), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(G274), .A3(new_n285), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n285), .B(G257), .C1(new_n460), .C2(new_n462), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n209), .B1(new_n273), .B2(new_n274), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT4), .ZN(new_n468));
  OAI21_X1  g0268(.A(G1698), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n391), .B2(new_n352), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n468), .A2(G1698), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n275), .A2(G244), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G283), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n469), .A2(new_n470), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n466), .B1(new_n474), .B2(new_n280), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n290), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(G200), .B2(new_n475), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n459), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT78), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G179), .ZN(new_n481));
  AOI211_X1 g0281(.A(new_n481), .B(new_n466), .C1(new_n280), .C2(new_n474), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n474), .A2(new_n280), .ZN(new_n483));
  INV_X1    g0283(.A(new_n466), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n315), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n459), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n459), .A2(new_n477), .A3(KEYINPUT78), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n480), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(G257), .B(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n490));
  OAI211_X1 g0290(.A(G250), .B(new_n276), .C1(new_n320), .C2(new_n321), .ZN(new_n491));
  INV_X1    g0291(.A(G294), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n490), .B(new_n491), .C1(new_n272), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n280), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n285), .B(G264), .C1(new_n460), .C2(new_n462), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n464), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n315), .ZN(new_n497));
  INV_X1    g0297(.A(new_n495), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n280), .B2(new_n493), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(new_n481), .A3(new_n464), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT84), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(new_n225), .B2(G107), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT23), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT23), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n501), .B(new_n504), .C1(new_n225), .C2(G107), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n503), .A2(new_n505), .B1(G116), .B2(new_n263), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n225), .B(G87), .C1(new_n320), .C2(new_n321), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n507), .A2(KEYINPUT22), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(KEYINPUT22), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT24), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT24), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n512), .B(new_n506), .C1(new_n508), .C2(new_n509), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n444), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n257), .A2(new_n451), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n515), .A2(KEYINPUT25), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(KEYINPUT25), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n516), .B(new_n517), .C1(new_n445), .C2(new_n451), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n497), .B(new_n500), .C1(new_n514), .C2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT21), .ZN(new_n520));
  OAI211_X1 g0320(.A(G257), .B(new_n276), .C1(new_n320), .C2(new_n321), .ZN(new_n521));
  INV_X1    g0321(.A(G303), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n521), .B1(new_n522), .B2(new_n275), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(G264), .A2(G1698), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n320), .B2(new_n321), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT82), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT82), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n275), .A2(new_n528), .A3(new_n525), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n285), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n285), .B(G270), .C1(new_n460), .C2(new_n462), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n464), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(G169), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G116), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n257), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n445), .B2(new_n535), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n251), .A2(new_n224), .B1(G20), .B2(new_n535), .ZN(new_n538));
  AOI21_X1  g0338(.A(G20), .B1(G33), .B2(G283), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n272), .A2(G97), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT83), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT83), .B1(new_n539), .B2(new_n540), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n538), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT20), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(KEYINPUT20), .B(new_n538), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n537), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n520), .B1(new_n534), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n537), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n545), .A2(new_n546), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n531), .A2(new_n533), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(G179), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n523), .B1(new_n529), .B2(new_n527), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n464), .B(new_n532), .C1(new_n554), .C2(new_n285), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n551), .A2(new_n555), .A3(KEYINPUT21), .A4(G169), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n519), .A2(new_n548), .A3(new_n553), .A4(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n514), .A2(new_n518), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n496), .A2(new_n290), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n427), .B1(new_n499), .B2(new_n464), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n551), .B1(G200), .B2(new_n555), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n552), .A2(G190), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(G250), .B1(new_n253), .B2(G45), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n280), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(G274), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n253), .A2(new_n570), .A3(G45), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n330), .A2(G1698), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI22_X1  g0374(.A1(new_n391), .A2(new_n574), .B1(new_n272), .B2(new_n535), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT79), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n275), .A2(new_n576), .A3(G244), .A4(G1698), .ZN(new_n577));
  OAI211_X1 g0377(.A(G244), .B(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT79), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n575), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT80), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n280), .B1(new_n580), .B2(KEYINPUT80), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n572), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G200), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n225), .B1(new_n323), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n208), .A2(new_n210), .A3(new_n451), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT81), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n587), .A2(KEYINPUT81), .A3(new_n588), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n275), .A2(new_n225), .A3(G68), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n586), .B1(new_n262), .B2(new_n210), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n252), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n358), .A2(new_n257), .ZN(new_n598));
  INV_X1    g0398(.A(new_n445), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G87), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(G190), .B(new_n572), .C1(new_n582), .C2(new_n583), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n585), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n481), .B(new_n572), .C1(new_n582), .C2(new_n583), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n597), .B(new_n598), .C1(new_n445), .C2(new_n358), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n579), .A2(new_n577), .ZN(new_n607));
  INV_X1    g0407(.A(new_n575), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT80), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n285), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n611), .A2(new_n581), .B1(new_n571), .B2(new_n569), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n605), .B(new_n606), .C1(new_n612), .C2(G169), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n558), .A2(new_n567), .A3(new_n604), .A4(new_n613), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n442), .A2(new_n489), .A3(new_n614), .ZN(G372));
  NAND2_X1  g0415(.A1(new_n604), .A2(new_n613), .ZN(new_n616));
  OAI21_X1  g0416(.A(KEYINPUT26), .B1(new_n616), .B2(new_n487), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT86), .B1(new_n482), .B2(new_n485), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n475), .A2(G179), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT86), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n619), .B(new_n620), .C1(new_n315), .C2(new_n475), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n459), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT85), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n597), .A2(new_n623), .A3(new_n598), .A4(new_n600), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n601), .A2(KEYINPUT85), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n585), .A2(new_n603), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n622), .A2(new_n626), .A3(new_n627), .A4(new_n613), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n617), .A2(new_n613), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n557), .A2(new_n563), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n603), .B1(new_n612), .B2(new_n427), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n625), .A2(new_n624), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n613), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n489), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n441), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n295), .B(KEYINPUT87), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n397), .A2(new_n420), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT18), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n397), .A2(new_n420), .A3(new_n423), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n345), .ZN(new_n643));
  INV_X1    g0443(.A(new_n363), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n348), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n439), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n366), .B1(new_n637), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n636), .A2(new_n648), .ZN(G369));
  NAND3_X1  g0449(.A1(new_n548), .A2(new_n553), .A3(new_n556), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n253), .A2(new_n225), .A3(G13), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT88), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n655));
  INV_X1    g0455(.A(G213), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G343), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT89), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n658), .A2(KEYINPUT89), .A3(G343), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n551), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n650), .B(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n565), .B2(new_n564), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n511), .A2(new_n513), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n252), .ZN(new_n669));
  INV_X1    g0469(.A(new_n518), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n663), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n563), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n519), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n519), .A2(new_n663), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n667), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n663), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n650), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n675), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n679), .A2(new_n683), .ZN(G399));
  NAND2_X1  g0484(.A1(new_n229), .A2(new_n284), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n588), .A2(G116), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n686), .A2(new_n253), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n223), .B2(new_n686), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT28), .Z(new_n691));
  NAND2_X1  g0491(.A1(new_n635), .A2(new_n680), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT29), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n618), .A2(new_n621), .ZN(new_n695));
  INV_X1    g0495(.A(new_n459), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT26), .B1(new_n633), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT91), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n613), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n459), .A2(new_n486), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n604), .A2(new_n701), .A3(new_n613), .A4(new_n627), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n698), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(KEYINPUT29), .B(new_n680), .C1(new_n703), .C2(new_n634), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n694), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n614), .A2(new_n489), .A3(new_n663), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n552), .A2(new_n475), .A3(G179), .A4(new_n499), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(new_n584), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n555), .A2(new_n481), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n475), .A2(new_n499), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n612), .A2(new_n710), .A3(new_n711), .A4(KEYINPUT30), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n552), .A2(new_n475), .A3(G179), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n584), .A3(new_n496), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n709), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n663), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT31), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g0518(.A(KEYINPUT90), .B(KEYINPUT31), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n718), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(G330), .B1(new_n706), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n705), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n691), .B1(new_n723), .B2(G1), .ZN(G364));
  NOR2_X1   g0524(.A1(new_n256), .A2(G20), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n253), .B1(new_n725), .B2(G45), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n686), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n229), .A2(new_n275), .ZN(new_n729));
  INV_X1    g0529(.A(G355), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n729), .A2(new_n730), .B1(G116), .B2(new_n229), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n229), .A2(new_n391), .ZN(new_n732));
  INV_X1    g0532(.A(G45), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n732), .B1(new_n733), .B2(new_n223), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n249), .A2(G45), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n224), .B1(G20), .B2(new_n315), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n728), .B1(new_n736), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n225), .B1(new_n744), .B2(G190), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n492), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n225), .A2(new_n290), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n481), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n225), .A2(G190), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n748), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI22_X1  g0553(.A1(G322), .A2(new_n750), .B1(new_n753), .B2(G311), .ZN(new_n754));
  INV_X1    g0554(.A(G283), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n427), .A2(G179), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n751), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n754), .B(new_n391), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n290), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n746), .B(new_n758), .C1(G326), .C2(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT33), .B(G317), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n762), .A2(KEYINPUT96), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n759), .A2(G190), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n762), .A2(KEYINPUT96), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n751), .A2(new_n744), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT95), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(KEYINPUT95), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n747), .A2(new_n756), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT94), .Z(new_n774));
  AOI22_X1  g0574(.A1(new_n772), .A2(G329), .B1(G303), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n761), .A2(new_n766), .A3(new_n775), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n749), .A2(new_n202), .B1(new_n752), .B2(new_n299), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT92), .ZN(new_n778));
  INV_X1    g0578(.A(new_n760), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n777), .A2(new_n778), .B1(new_n201), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n778), .B2(new_n777), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT93), .Z(new_n782));
  NAND2_X1  g0582(.A1(new_n768), .A2(G159), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT32), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n275), .B1(new_n757), .B2(new_n451), .C1(new_n208), .C2(new_n773), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n745), .A2(new_n210), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n764), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n788), .B2(new_n203), .ZN(new_n789));
  OR3_X1    g0589(.A1(new_n784), .A2(new_n785), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n776), .B1(new_n782), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n743), .B1(new_n791), .B2(new_n740), .ZN(new_n792));
  INV_X1    g0592(.A(new_n739), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n666), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n728), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n667), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n666), .A2(G330), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(G396));
  NAND2_X1  g0598(.A1(new_n644), .A2(new_n680), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n370), .B1(new_n680), .B2(new_n369), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n363), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n692), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n802), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n680), .B(new_n804), .C1(new_n629), .C2(new_n634), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n806), .A2(new_n721), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n728), .B1(new_n806), .B2(new_n721), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n740), .A2(new_n737), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n795), .B1(new_n299), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n804), .A2(new_n738), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n787), .B1(new_n779), .B2(new_n522), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n391), .B1(new_n749), .B2(new_n492), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n208), .A2(new_n757), .B1(new_n752), .B2(new_n535), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(new_n774), .C2(G107), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(new_n771), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n814), .B(new_n819), .C1(G283), .C2(new_n764), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n821), .A2(KEYINPUT97), .ZN(new_n822));
  XNOR2_X1  g0622(.A(KEYINPUT98), .B(G143), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n750), .A2(new_n823), .B1(new_n753), .B2(G159), .ZN(new_n824));
  INV_X1    g0624(.A(G137), .ZN(new_n825));
  INV_X1    g0625(.A(G150), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n824), .B1(new_n779), .B2(new_n825), .C1(new_n826), .C2(new_n788), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT34), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n772), .A2(G132), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n275), .B1(new_n745), .B2(new_n202), .C1(new_n203), .C2(new_n757), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n774), .B2(G50), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n821), .A2(KEYINPUT97), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n822), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n812), .B(new_n813), .C1(new_n740), .C2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n809), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G384));
  NOR2_X1   g0639(.A1(new_n725), .A2(new_n253), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT103), .ZN(new_n841));
  INV_X1    g0641(.A(new_n719), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n715), .B2(new_n663), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n715), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n841), .B1(new_n706), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n558), .A2(new_n567), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n480), .A2(new_n488), .A3(new_n487), .ZN(new_n849));
  INV_X1    g0649(.A(new_n616), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n680), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n851), .A2(KEYINPUT103), .A3(new_n845), .A4(new_n844), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT100), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n345), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(KEYINPUT100), .B(new_n313), .C1(new_n342), .C2(new_n344), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n663), .A2(new_n313), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n347), .B2(new_n346), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT101), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT101), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n855), .A2(new_n858), .A3(new_n861), .A4(new_n856), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n857), .B1(new_n344), .B2(new_n342), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n802), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n203), .B1(new_n378), .B2(new_n380), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n434), .B1(new_n867), .B2(new_n388), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n374), .B1(new_n432), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n658), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n421), .A2(KEYINPUT18), .B1(new_n431), .B2(new_n438), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n872), .B1(new_n873), .B2(new_n424), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n398), .A2(new_n400), .A3(new_n658), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT37), .B1(new_n436), .B2(new_n429), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n421), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n416), .A2(new_n418), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n419), .A2(new_n315), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n658), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n430), .B1(new_n880), .B2(new_n869), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n866), .B1(new_n874), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT102), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n440), .A2(new_n871), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n877), .A2(new_n882), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n884), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n885), .B1(new_n884), .B2(new_n888), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n853), .B(new_n865), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT40), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT104), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT104), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n891), .A2(new_n895), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n877), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n638), .A2(new_n430), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n875), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n898), .B1(KEYINPUT37), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n875), .B1(new_n642), .B2(new_n439), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n866), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n888), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n853), .A2(new_n865), .A3(new_n905), .A4(KEYINPUT40), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n897), .A2(new_n906), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT105), .Z(new_n908));
  AND2_X1   g0708(.A1(new_n853), .A2(new_n441), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(G330), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n884), .A2(new_n888), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT39), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n904), .A2(new_n915), .A3(new_n888), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n855), .A2(new_n856), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n920), .A2(new_n663), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n799), .B(KEYINPUT99), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n805), .A2(new_n923), .B1(new_n863), .B2(new_n864), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n890), .B2(new_n889), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n641), .A2(new_n870), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n694), .A2(new_n441), .A3(new_n704), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n648), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n927), .B(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n840), .B1(new_n912), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n930), .B2(new_n912), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n456), .A2(KEYINPUT35), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n456), .A2(KEYINPUT35), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n933), .A2(G116), .A3(new_n226), .A4(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT36), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n384), .A2(new_n222), .A3(new_n299), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n203), .A2(G50), .ZN(new_n938));
  OAI211_X1 g0738(.A(G1), .B(new_n256), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n932), .A2(new_n936), .A3(new_n939), .ZN(G367));
  OAI21_X1  g0740(.A(new_n849), .B1(new_n459), .B2(new_n680), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n622), .A2(new_n663), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n943), .A2(new_n682), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT42), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n519), .B1(new_n941), .B2(new_n942), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n680), .B1(new_n947), .B2(new_n701), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n944), .A2(new_n945), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n632), .A2(new_n663), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(new_n613), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n626), .A2(new_n951), .A3(new_n613), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n950), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n950), .A2(new_n957), .A3(new_n955), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n678), .A2(new_n943), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT106), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n959), .A2(new_n960), .B1(KEYINPUT106), .B2(new_n961), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n685), .B(KEYINPUT41), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n683), .A2(new_n943), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT44), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT45), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT107), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n683), .A2(new_n970), .A3(new_n943), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n970), .B1(new_n683), .B2(new_n943), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n973), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n975), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n968), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n678), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n677), .B(new_n681), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(new_n667), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n722), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n968), .A2(new_n974), .A3(new_n976), .A4(new_n679), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n978), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n966), .B1(new_n983), .B2(new_n723), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n965), .B1(new_n984), .B2(new_n727), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(KEYINPUT108), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT108), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n965), .B(new_n987), .C1(new_n984), .C2(new_n727), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n732), .A2(new_n241), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n741), .B1(new_n229), .B2(new_n358), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n728), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n745), .A2(new_n203), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n391), .B(new_n993), .C1(G150), .C2(new_n750), .ZN(new_n994));
  INV_X1    g0794(.A(new_n757), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n995), .A2(G77), .B1(new_n768), .B2(G137), .ZN(new_n996));
  INV_X1    g0796(.A(new_n773), .ZN(new_n997));
  AOI22_X1  g0797(.A1(G58), .A2(new_n997), .B1(new_n753), .B2(G50), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n760), .A2(new_n823), .B1(new_n764), .B2(G159), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n994), .A2(new_n996), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n275), .B1(new_n768), .B2(G317), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n788), .B2(new_n492), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n779), .A2(new_n818), .B1(new_n745), .B2(new_n451), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G303), .A2(new_n750), .B1(new_n995), .B2(G97), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(new_n755), .C2(new_n752), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n773), .A2(KEYINPUT46), .A3(new_n535), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n774), .A2(G116), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1007), .B1(new_n1008), .B2(KEYINPUT46), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1000), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT47), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n992), .B1(new_n1011), .B2(new_n740), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n952), .A2(new_n739), .A3(new_n953), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n989), .A2(new_n1014), .ZN(G387));
  INV_X1    g0815(.A(new_n980), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n677), .A2(new_n739), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n729), .A2(new_n687), .B1(G107), .B2(new_n229), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n238), .A2(new_n733), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n260), .A2(new_n1020), .A3(G50), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n733), .B1(new_n203), .B2(new_n299), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1021), .A2(new_n688), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1020), .B1(new_n260), .B2(G50), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n732), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1018), .B1(new_n1019), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n728), .B1(new_n1026), .B2(new_n742), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n773), .A2(new_n299), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n749), .A2(new_n201), .B1(new_n767), .B2(new_n826), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G68), .C2(new_n753), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n760), .A2(G159), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n745), .A2(new_n358), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n391), .B(new_n1032), .C1(G97), .C2(new_n995), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n261), .A2(new_n764), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1030), .A2(new_n1031), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n275), .B1(new_n768), .B2(G326), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n773), .A2(new_n492), .B1(new_n745), .B2(new_n755), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G317), .A2(new_n750), .B1(new_n753), .B2(G303), .ZN(new_n1038));
  XOR2_X1   g0838(.A(KEYINPUT110), .B(G322), .Z(new_n1039));
  OAI221_X1 g0839(.A(new_n1038), .B1(new_n779), .B2(new_n1039), .C1(new_n818), .C2(new_n788), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT49), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1036), .B1(new_n535), .B2(new_n757), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1035), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1027), .B1(new_n1047), .B2(new_n740), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1016), .A2(new_n727), .B1(new_n1017), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n723), .A2(new_n1016), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n686), .B1(new_n722), .B2(new_n980), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(G393));
  NAND3_X1  g0852(.A1(new_n978), .A2(new_n727), .A3(new_n982), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n246), .A2(new_n732), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n741), .B1(new_n229), .B2(new_n210), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n728), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n275), .B1(new_n757), .B2(new_n208), .C1(new_n788), .C2(new_n201), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n745), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1057), .B1(G77), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n752), .A2(new_n260), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n768), .B2(new_n823), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1059), .B(new_n1061), .C1(new_n203), .C2(new_n773), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n750), .A2(G159), .B1(G150), .B2(new_n760), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT51), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n750), .A2(G311), .B1(G317), .B2(new_n760), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT52), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n745), .A2(new_n535), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n391), .B1(new_n757), .B2(new_n451), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(G303), .C2(new_n764), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n753), .A2(G294), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1039), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n768), .A2(new_n1071), .B1(new_n997), .B2(G283), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1069), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1062), .A2(new_n1064), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1056), .B1(new_n1074), .B2(new_n740), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n943), .B2(new_n793), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n983), .A2(new_n686), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n981), .B1(new_n978), .B2(new_n982), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1053), .B(new_n1076), .C1(new_n1077), .C2(new_n1078), .ZN(G390));
  OAI211_X1 g0879(.A(new_n914), .B(new_n916), .C1(new_n924), .C2(new_n921), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n721), .A2(new_n802), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n863), .A2(new_n864), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n680), .B(new_n801), .C1(new_n703), .C2(new_n634), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT111), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1084), .A2(new_n1085), .A3(new_n799), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n1084), .B2(new_n799), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n863), .A2(new_n864), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n921), .B1(new_n904), .B2(new_n888), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1080), .B(new_n1083), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n865), .A2(G330), .A3(new_n853), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1084), .A2(new_n799), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(KEYINPUT111), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1084), .A2(new_n1085), .A3(new_n799), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(new_n1082), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n1090), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1095), .B1(new_n1100), .B2(new_n1080), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1093), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n853), .A2(G330), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n928), .B(new_n648), .C1(new_n442), .C2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1088), .B1(new_n1103), .B2(new_n802), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n1107), .A3(new_n1083), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n805), .A2(new_n923), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1110), .B1(new_n1094), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1102), .A2(new_n1105), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1105), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n1093), .B2(new_n1101), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1114), .A2(new_n1116), .A3(new_n686), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT116), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1109), .A2(new_n1088), .B1(new_n920), .B2(new_n663), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1099), .A2(new_n1090), .B1(new_n1119), .B2(new_n917), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n727), .B(new_n1092), .C1(new_n1120), .C2(new_n1095), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(KEYINPUT112), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1100), .A2(new_n1080), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1094), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT112), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1124), .A2(new_n1125), .A3(new_n727), .A4(new_n1092), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n917), .A2(new_n737), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n810), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n728), .B1(new_n261), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n772), .A2(G125), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1132), .A2(new_n752), .B1(new_n757), .B2(new_n201), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n391), .B(new_n1133), .C1(G132), .C2(new_n750), .ZN(new_n1134));
  INV_X1    g0934(.A(G128), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n788), .A2(new_n825), .B1(new_n779), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G159), .B2(new_n1058), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n773), .A2(new_n826), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1131), .A2(new_n1134), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n275), .B1(new_n774), .B2(G87), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT113), .Z(new_n1142));
  AOI22_X1  g0942(.A1(G68), .A2(new_n995), .B1(new_n753), .B2(G97), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n779), .B2(new_n755), .C1(new_n451), .C2(new_n788), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G294), .B2(new_n772), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n749), .A2(new_n535), .B1(new_n745), .B2(new_n299), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT114), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1140), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1130), .B1(new_n1149), .B2(new_n740), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT115), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1128), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1118), .B1(new_n1127), .B2(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(KEYINPUT116), .B(new_n1152), .C1(new_n1122), .C2(new_n1126), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1117), .B1(new_n1154), .B2(new_n1155), .ZN(G378));
  AOI21_X1  g0956(.A(new_n1104), .B1(new_n1102), .B2(new_n1113), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n295), .A2(KEYINPUT87), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n295), .A2(KEYINPUT87), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n367), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n268), .A2(new_n870), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT55), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1162), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n637), .A2(new_n367), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1163), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n906), .A2(G330), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n897), .B2(new_n1172), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n891), .A2(new_n895), .A3(new_n892), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n895), .B1(new_n891), .B2(new_n892), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1172), .B(new_n1171), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n927), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1172), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n1170), .A3(new_n1169), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n927), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n1181), .A3(new_n1176), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1157), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n686), .B1(new_n1183), .B2(KEYINPUT57), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT57), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1185), .B(new_n1157), .C1(new_n1182), .C2(new_n1178), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1169), .A2(new_n737), .A3(new_n1170), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n772), .A2(G283), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n779), .A2(new_n535), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n993), .B(new_n1191), .C1(G97), .C2(new_n764), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n749), .A2(new_n451), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT117), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n202), .A2(new_n757), .B1(new_n752), .B2(new_n358), .ZN(new_n1195));
  NOR4_X1   g0995(.A1(new_n1195), .A2(new_n1028), .A3(G41), .A4(new_n275), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1190), .A2(new_n1192), .A3(new_n1194), .A4(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT58), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n201), .B1(new_n320), .B2(G41), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT118), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n753), .A2(G137), .B1(G132), .B2(new_n764), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT119), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n760), .A2(G125), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n745), .A2(new_n826), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n1135), .A2(new_n749), .B1(new_n773), .B2(new_n1132), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(KEYINPUT59), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n768), .A2(G124), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G33), .B(G41), .C1(new_n995), .C2(G159), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT59), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1211), .B(new_n1212), .C1(new_n1208), .C2(new_n1213), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n1210), .A2(new_n1214), .B1(new_n1198), .B2(new_n1197), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n740), .B1(new_n1202), .B2(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT120), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n795), .B(new_n1217), .C1(new_n201), .C2(new_n810), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1188), .A2(new_n727), .B1(new_n1189), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1187), .A2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n772), .A2(G128), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n749), .A2(new_n825), .B1(new_n752), .B2(new_n826), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n391), .B(new_n1222), .C1(G58), .C2(new_n995), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n788), .A2(new_n1132), .B1(new_n201), .B2(new_n745), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G132), .B2(new_n760), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n774), .A2(G159), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1221), .A2(new_n1223), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n749), .A2(new_n755), .B1(new_n752), .B2(new_n451), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n275), .B(new_n1228), .C1(G77), .C2(new_n995), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n774), .A2(G97), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(new_n522), .C2(new_n771), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1032), .B1(new_n764), .B2(G116), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n492), .B2(new_n779), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1227), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n740), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1235), .B(new_n728), .C1(G68), .C2(new_n1129), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1088), .B2(new_n737), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1113), .B2(new_n727), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n966), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1115), .A2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1113), .A2(new_n1105), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1238), .B1(new_n1240), .B2(new_n1241), .ZN(G381));
  INV_X1    g1042(.A(G390), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n989), .A2(new_n1014), .A3(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(G393), .A2(G396), .ZN(new_n1245));
  OR4_X1    g1045(.A1(G384), .A2(new_n1244), .A3(G381), .A4(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1187), .A2(new_n1219), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1117), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1127), .A2(new_n1153), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(KEYINPUT116), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1127), .A2(new_n1118), .A3(new_n1153), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1248), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1247), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT122), .ZN(new_n1254));
  OR3_X1    g1054(.A1(new_n1246), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1254), .B1(new_n1246), .B2(new_n1253), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(G407));
  INV_X1    g1057(.A(new_n1253), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n656), .A2(G343), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n1259), .B(KEYINPUT123), .Z(new_n1260));
  AOI21_X1  g1060(.A(new_n656), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G407), .A2(new_n1261), .ZN(G409));
  INV_X1    g1062(.A(KEYINPUT126), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G378), .B(new_n1219), .C1(new_n1184), .C2(new_n1186), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1157), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1188), .A2(new_n1239), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1188), .A2(new_n727), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1189), .A2(new_n1218), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1252), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1259), .B1(new_n1264), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1113), .B2(new_n1105), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1108), .A2(new_n1104), .A3(new_n1112), .A4(KEYINPUT60), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1273), .A2(new_n686), .A3(new_n1115), .A4(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(G384), .A3(new_n1238), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1275), .B2(new_n1238), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n1263), .B(KEYINPUT62), .C1(new_n1271), .C2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1264), .A2(new_n1270), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1259), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n1282), .A3(new_n1279), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT126), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT127), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1260), .B1(new_n1264), .B2(new_n1270), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1279), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1288), .A2(new_n1284), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1286), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1287), .A2(new_n1286), .A3(new_n1289), .ZN(new_n1291));
  OAI22_X1  g1091(.A1(new_n1280), .A2(new_n1285), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1260), .A2(G2897), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1278), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1259), .A2(G2897), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1295), .A2(new_n1276), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1287), .B1(new_n1294), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G387), .A2(G390), .ZN(new_n1299));
  XOR2_X1   g1099(.A(G393), .B(G396), .Z(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1299), .A2(new_n1244), .A3(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1243), .B1(new_n989), .B2(new_n1014), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1014), .ZN(new_n1304));
  AOI211_X1 g1104(.A(new_n1304), .B(G390), .C1(new_n986), .C2(new_n988), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1300), .B1(new_n1303), .B2(new_n1305), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1298), .A2(new_n1307), .A3(KEYINPUT61), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT124), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1294), .A2(new_n1297), .A3(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1310), .B1(new_n1294), .B2(new_n1297), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT61), .B1(new_n1309), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1283), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1260), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1288), .A2(new_n1315), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1281), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT125), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1287), .A2(KEYINPUT125), .A3(new_n1318), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1314), .A2(new_n1316), .A3(new_n1321), .A4(new_n1322), .ZN(new_n1323));
  AOI22_X1  g1123(.A1(new_n1292), .A2(new_n1308), .B1(new_n1323), .B2(new_n1307), .ZN(G405));
  NAND2_X1  g1124(.A1(G375), .A2(new_n1252), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1264), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1307), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1328), .A2(new_n1264), .A3(new_n1325), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1327), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1288), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1327), .A2(new_n1279), .A3(new_n1329), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(G402));
endmodule


