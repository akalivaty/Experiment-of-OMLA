//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G97), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT64), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  OR3_X1    g0034(.A1(new_n228), .A2(new_n207), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n212), .A2(new_n226), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n221), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT2), .B(G226), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT67), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G58), .B(G77), .Z(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(KEYINPUT7), .B1(new_n257), .B2(new_n207), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(G68), .B1(new_n258), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n220), .A2(new_n214), .ZN(new_n266));
  OAI21_X1  g0066(.A(G20), .B1(new_n266), .B2(new_n201), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G159), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(KEYINPUT16), .B1(new_n265), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n231), .A2(new_n232), .A3(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n261), .A2(new_n207), .A3(new_n262), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT7), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n214), .B1(new_n277), .B2(new_n263), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n267), .A2(KEYINPUT16), .A3(new_n269), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT77), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n274), .ZN(new_n282));
  INV_X1    g0082(.A(new_n279), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n282), .B1(new_n265), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT77), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT16), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(new_n278), .B2(new_n270), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  XOR2_X1   g0092(.A(KEYINPUT8), .B(G58), .Z(new_n293));
  NAND2_X1  g0093(.A1(new_n206), .A2(G20), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n231), .A2(new_n290), .A3(new_n232), .A4(new_n273), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT78), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT78), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n281), .A2(new_n288), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT79), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n281), .A2(new_n288), .A3(new_n302), .A4(KEYINPUT79), .ZN(new_n306));
  INV_X1    g0106(.A(G41), .ZN(new_n307));
  INV_X1    g0107(.A(G45), .ZN(new_n308));
  AOI21_X1  g0108(.A(G1), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G41), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n310), .A2(G1), .A3(G13), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n311), .A3(G274), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(G232), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(G226), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G87), .ZN(new_n317));
  OR2_X1    g0117(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n318));
  NAND2_X1  g0118(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n318), .B(new_n319), .C1(new_n255), .C2(new_n256), .ZN(new_n320));
  INV_X1    g0120(.A(G223), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n316), .B(new_n317), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n233), .A2(new_n310), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n315), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G179), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n326), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n305), .A2(new_n306), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT18), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT17), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n322), .A2(new_n324), .ZN(new_n333));
  INV_X1    g0133(.A(new_n315), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G190), .ZN(new_n336));
  AOI211_X1 g0136(.A(new_n336), .B(new_n315), .C1(new_n322), .C2(new_n324), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n331), .B1(new_n303), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n284), .A2(new_n287), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n340), .A2(KEYINPUT77), .B1(new_n301), .B2(new_n299), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n335), .A2(new_n337), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n341), .A2(KEYINPUT17), .A3(new_n288), .A4(new_n342), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT18), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n305), .A2(new_n345), .A3(new_n306), .A4(new_n328), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n330), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  XOR2_X1   g0148(.A(KEYINPUT68), .B(G1698), .Z(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G226), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G232), .A2(G1698), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n257), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G33), .A2(G97), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT75), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT75), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(G33), .A3(G97), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n324), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT13), .ZN(new_n359));
  INV_X1    g0159(.A(new_n312), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n311), .A2(new_n313), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(G238), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n358), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n359), .B1(new_n358), .B2(new_n362), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT14), .B1(new_n366), .B2(new_n327), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(G179), .ZN(new_n368));
  INV_X1    g0168(.A(new_n365), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n363), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT14), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(G169), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n367), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n268), .A2(G50), .B1(G20), .B2(new_n214), .ZN(new_n374));
  INV_X1    g0174(.A(G77), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n207), .A2(G33), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n377), .A2(new_n274), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n378), .A2(KEYINPUT11), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n291), .A2(new_n214), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT12), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(KEYINPUT11), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n296), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(G68), .A3(new_n294), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n385), .B(KEYINPUT76), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n373), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n370), .A2(G200), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n369), .A2(G190), .A3(new_n363), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n390), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n293), .A2(new_n268), .B1(G20), .B2(G77), .ZN(new_n395));
  XNOR2_X1  g0195(.A(KEYINPUT15), .B(G87), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n260), .A2(G20), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n282), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n384), .A2(G77), .A3(new_n294), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n290), .A2(G77), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n360), .B1(G244), .B2(new_n361), .ZN(new_n404));
  INV_X1    g0204(.A(G1698), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(new_n261), .B2(new_n262), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G238), .ZN(new_n407));
  INV_X1    g0207(.A(G107), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n261), .A2(new_n262), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT72), .B1(new_n320), .B2(new_n221), .ZN(new_n411));
  OR3_X1    g0211(.A1(new_n320), .A2(KEYINPUT72), .A3(new_n221), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n404), .B1(new_n413), .B2(new_n323), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n403), .B1(new_n414), .B2(new_n336), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(G200), .B2(new_n414), .ZN(new_n416));
  OR2_X1    g0216(.A1(new_n414), .A2(G179), .ZN(new_n417));
  INV_X1    g0217(.A(new_n403), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n414), .A2(new_n327), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n394), .A2(new_n416), .A3(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n294), .A2(G50), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n296), .A2(new_n424), .B1(G50), .B2(new_n290), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n203), .A2(G20), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n268), .A2(G150), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n289), .B2(new_n376), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT70), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n426), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n429), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n282), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n425), .B1(new_n433), .B2(KEYINPUT71), .ZN(new_n434));
  INV_X1    g0234(.A(new_n432), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n274), .B1(new_n435), .B2(new_n430), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT71), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n434), .A2(KEYINPUT9), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT73), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n434), .A2(KEYINPUT73), .A3(KEYINPUT9), .A4(new_n438), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n434), .A2(new_n438), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT9), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n257), .A2(G77), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n349), .A2(G222), .B1(G223), .B2(G1698), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n447), .B1(new_n448), .B2(new_n257), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT69), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(KEYINPUT69), .B(new_n447), .C1(new_n448), .C2(new_n257), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n324), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n360), .B1(G226), .B2(new_n361), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(G190), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n454), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G200), .ZN(new_n457));
  NAND2_X1  g0257(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n446), .A2(new_n455), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n423), .B1(new_n443), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n441), .A2(new_n442), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n457), .A2(new_n455), .A3(new_n458), .ZN(new_n462));
  INV_X1    g0262(.A(new_n423), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .A4(new_n446), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n456), .A2(new_n327), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n467), .B(new_n444), .C1(G179), .C2(new_n456), .ZN(new_n468));
  AND4_X1   g0268(.A1(new_n348), .A2(new_n422), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n308), .A2(G1), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT81), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(new_n307), .A3(KEYINPUT5), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT5), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT81), .B1(new_n473), .B2(G41), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(G41), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n470), .B(new_n472), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(G257), .A3(new_n311), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT82), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT4), .ZN(new_n480));
  INV_X1    g0280(.A(G244), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n320), .B2(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n406), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n320), .A2(new_n480), .A3(new_n481), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n324), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n311), .A2(G274), .ZN(new_n487));
  OR2_X1    g0287(.A1(new_n476), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n479), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G169), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n479), .A2(new_n486), .A3(G179), .A4(new_n488), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n222), .A2(new_n408), .ZN(new_n493));
  NOR2_X1   g0293(.A1(G97), .A2(G107), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n408), .A2(KEYINPUT6), .A3(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(G20), .B1(G77), .B2(new_n268), .ZN(new_n498));
  OAI21_X1  g0298(.A(G107), .B1(new_n258), .B2(new_n264), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n274), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT85), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n260), .A2(G1), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n296), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G97), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n290), .A2(G97), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT80), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n501), .A2(new_n502), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n282), .B1(new_n498), .B2(new_n499), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(new_n507), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT85), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n490), .A2(new_n491), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n479), .A2(new_n486), .A3(G190), .A4(new_n488), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n509), .A2(new_n510), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n489), .A2(KEYINPUT83), .A3(G200), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT83), .B1(new_n489), .B2(G200), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT84), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(KEYINPUT84), .B(new_n515), .C1(new_n516), .C2(new_n517), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n512), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(G244), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G116), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n523), .B(new_n524), .C1(new_n320), .C2(new_n215), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n324), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n206), .A2(G45), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n311), .A2(G250), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n487), .B2(new_n527), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT86), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(G179), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n526), .A2(KEYINPUT86), .A3(new_n530), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI211_X1 g0336(.A(new_n532), .B(new_n529), .C1(new_n324), .C2(new_n525), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT86), .B1(new_n526), .B2(new_n530), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n327), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT88), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n494), .A2(new_n216), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT19), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT87), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT87), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT19), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n354), .A2(new_n356), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n541), .B1(new_n546), .B2(G20), .ZN(new_n547));
  AOI21_X1  g0347(.A(G20), .B1(new_n261), .B2(new_n262), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n398), .A2(G97), .ZN(new_n549));
  XNOR2_X1  g0349(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n548), .A2(G68), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n282), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n397), .A2(new_n290), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n296), .A2(new_n396), .A3(new_n503), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n540), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NOR4_X1   g0357(.A1(new_n552), .A2(KEYINPUT88), .A3(new_n553), .A4(new_n555), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n536), .B(new_n539), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n504), .A2(G87), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n533), .A2(G190), .A3(new_n535), .ZN(new_n562));
  OAI21_X1  g0362(.A(G200), .B1(new_n537), .B2(new_n538), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT23), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(new_n408), .A3(G20), .ZN(new_n568));
  INV_X1    g0368(.A(G116), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n566), .B(new_n568), .C1(new_n569), .C2(new_n376), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT90), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n398), .A2(G116), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n573), .A2(KEYINPUT90), .A3(new_n568), .A4(new_n566), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT24), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT22), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n548), .A2(new_n577), .A3(G87), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n207), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT22), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n575), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n576), .B1(new_n575), .B2(new_n581), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n274), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT25), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n290), .B2(G107), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n408), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n504), .A2(G107), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n409), .A2(G257), .A3(G1698), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G294), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n217), .C2(new_n320), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n591), .A2(new_n324), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n476), .A2(G264), .A3(new_n311), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n488), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(G200), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n324), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n596), .A2(G190), .A3(new_n488), .A4(new_n593), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n584), .A2(new_n588), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n588), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n575), .A2(new_n581), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT24), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n575), .A2(new_n576), .A3(new_n581), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n599), .B1(new_n603), .B2(new_n274), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n596), .A2(new_n488), .A3(new_n593), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n327), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n596), .A2(new_n534), .A3(new_n488), .A4(new_n593), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n598), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT21), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n257), .A2(new_n223), .ZN(new_n611));
  XNOR2_X1  g0411(.A(KEYINPUT89), .B(G303), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n611), .A2(new_n349), .B1(new_n257), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n406), .A2(G264), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n323), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n476), .A2(G270), .A3(new_n311), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n488), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(G169), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n504), .A2(G116), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n291), .A2(new_n569), .ZN(new_n620));
  AOI21_X1  g0420(.A(G20), .B1(G33), .B2(G283), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n260), .A2(G97), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n621), .A2(new_n622), .B1(G20), .B2(new_n569), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n623), .A2(new_n274), .A3(KEYINPUT20), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT20), .B1(new_n623), .B2(new_n274), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n619), .B(new_n620), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n610), .B1(new_n618), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n617), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n611), .A2(new_n349), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n257), .A2(new_n612), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n614), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n324), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n629), .A2(new_n633), .A3(G190), .ZN(new_n634));
  OAI21_X1  g0434(.A(G200), .B1(new_n615), .B2(new_n617), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(new_n635), .A3(new_n627), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n629), .A2(new_n633), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n637), .A2(KEYINPUT21), .A3(G169), .A4(new_n626), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n615), .A2(new_n617), .A3(new_n534), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n626), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n628), .A2(new_n636), .A3(new_n638), .A4(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n565), .A2(new_n609), .A3(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n469), .A2(new_n522), .A3(new_n642), .ZN(G372));
  NAND2_X1  g0443(.A1(new_n520), .A2(new_n521), .ZN(new_n644));
  INV_X1    g0444(.A(new_n512), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n628), .A2(new_n640), .A3(new_n638), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT91), .ZN(new_n647));
  INV_X1    g0447(.A(new_n608), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n584), .A2(new_n588), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n604), .A2(new_n608), .A3(KEYINPUT91), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n531), .A2(new_n327), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n536), .B(new_n653), .C1(new_n557), .C2(new_n558), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n531), .A2(G200), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n561), .A2(new_n562), .A3(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n654), .A2(new_n598), .A3(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n644), .A2(new_n645), .A3(new_n652), .A4(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n559), .A2(new_n564), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n512), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n514), .B1(new_n490), .B2(new_n491), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n654), .A3(new_n656), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n654), .B1(new_n663), .B2(KEYINPUT26), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n469), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT92), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n303), .A2(new_n328), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(new_n345), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n389), .B1(new_n392), .B2(new_n420), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n672), .B1(new_n673), .B2(new_n344), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n468), .B1(new_n674), .B2(new_n465), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT93), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n668), .A2(KEYINPUT92), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n669), .A2(new_n677), .A3(new_n678), .ZN(G369));
  NAND3_X1  g0479(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT27), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n682), .A2(new_n206), .A3(new_n207), .A4(G13), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n681), .A2(G213), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT94), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT95), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(G343), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(G343), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OR3_X1    g0491(.A1(new_n646), .A2(new_n627), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT96), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n691), .A2(new_n627), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n692), .B(new_n693), .C1(new_n641), .C2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G330), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n609), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n604), .B2(new_n691), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n648), .A2(new_n649), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n701), .B1(new_n702), .B2(new_n691), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  OR3_X1    g0504(.A1(new_n650), .A2(new_n651), .A3(new_n690), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n646), .A2(new_n690), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n700), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n210), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n541), .A2(G116), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G1), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n227), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n690), .B1(new_n658), .B2(new_n665), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n663), .A2(KEYINPUT26), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n512), .A2(new_n659), .A3(new_n559), .A4(new_n564), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(new_n654), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT97), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n646), .A2(new_n702), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n644), .A2(new_n645), .A3(new_n657), .A4(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT97), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n719), .A2(new_n725), .A3(new_n654), .A4(new_n720), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n722), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n717), .B1(new_n727), .B2(new_n691), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n718), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n644), .A2(new_n645), .A3(new_n642), .A4(new_n691), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n479), .A2(new_n486), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n537), .A2(new_n538), .ZN(new_n732));
  INV_X1    g0532(.A(new_n605), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n731), .A2(new_n732), .A3(new_n639), .A4(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n479), .A2(new_n486), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n605), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n738), .A2(KEYINPUT30), .A3(new_n639), .A4(new_n732), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n605), .A2(new_n534), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n531), .B1(new_n615), .B2(new_n617), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n489), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n736), .A2(new_n739), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n690), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n734), .A2(new_n735), .B1(new_n489), .B2(new_n742), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n691), .B1(new_n748), .B2(new_n739), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT31), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n730), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G330), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n729), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n715), .B1(new_n754), .B2(G1), .ZN(G364));
  INV_X1    g0555(.A(G13), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n206), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n710), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n699), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n697), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(G330), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n760), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n709), .A2(new_n257), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n770), .A2(G355), .B1(new_n569), .B2(new_n709), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n709), .A2(new_n409), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n228), .B2(G45), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n253), .A2(new_n308), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n234), .B1(G20), .B2(new_n327), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n766), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n769), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n207), .A2(new_n534), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G190), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  INV_X1    g0582(.A(G322), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n779), .A2(G190), .A3(new_n332), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n257), .B1(new_n781), .B2(new_n782), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n779), .A2(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G190), .ZN(new_n787));
  XNOR2_X1  g0587(.A(KEYINPUT33), .B(G317), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT100), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n789), .B2(new_n788), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n207), .A2(G179), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n792), .A2(new_n780), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT98), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(KEYINPUT98), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n785), .B(new_n791), .C1(G329), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n786), .A2(new_n336), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n792), .A2(new_n336), .A3(G200), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n799), .A2(G326), .B1(new_n801), .B2(G283), .ZN(new_n802));
  INV_X1    g0602(.A(G294), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n336), .A2(G179), .A3(G200), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n207), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n792), .A2(G190), .A3(G200), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(KEYINPUT99), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(KEYINPUT99), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n806), .B1(G303), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G159), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n796), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT32), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n811), .A2(G87), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n409), .B1(new_n784), .B2(new_n220), .ZN(new_n817));
  INV_X1    g0617(.A(new_n781), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(G77), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n805), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G97), .A2(new_n820), .B1(new_n799), .B2(G50), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n800), .A2(new_n408), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G68), .B2(new_n787), .ZN(new_n823));
  AND4_X1   g0623(.A1(new_n816), .A2(new_n819), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n798), .A2(new_n812), .B1(new_n815), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n776), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n778), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n763), .B1(new_n768), .B2(new_n827), .ZN(G396));
  NAND2_X1  g0628(.A1(new_n418), .A2(new_n690), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT103), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n829), .B(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n420), .B1(new_n831), .B2(new_n416), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n421), .A2(new_n691), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n716), .B(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n760), .B1(new_n835), .B2(new_n752), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n752), .B2(new_n835), .ZN(new_n837));
  INV_X1    g0637(.A(new_n784), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n409), .B1(new_n838), .B2(G294), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n839), .B1(new_n569), .B2(new_n781), .C1(new_n796), .C2(new_n782), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n787), .A2(G283), .B1(new_n799), .B2(G303), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n841), .B1(new_n216), .B2(new_n800), .C1(new_n222), .C2(new_n805), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n840), .B(new_n842), .C1(G107), .C2(new_n811), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n838), .A2(G143), .B1(new_n818), .B2(G159), .ZN(new_n844));
  INV_X1    g0644(.A(new_n787), .ZN(new_n845));
  INV_X1    g0645(.A(G150), .ZN(new_n846));
  INV_X1    g0646(.A(G137), .ZN(new_n847));
  INV_X1    g0647(.A(new_n799), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n844), .B1(new_n845), .B2(new_n846), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT101), .Z(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(KEYINPUT34), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n257), .B1(new_n797), .B2(G132), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT102), .Z(new_n853));
  NOR2_X1   g0653(.A1(new_n800), .A2(new_n214), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(G58), .B2(new_n820), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n810), .B2(new_n202), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n851), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n850), .A2(KEYINPUT34), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n843), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n826), .A2(new_n765), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n859), .A2(new_n826), .B1(G77), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n834), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(new_n765), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n760), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n837), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT104), .Z(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(G384));
  NOR2_X1   g0667(.A1(new_n757), .A2(new_n206), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n305), .A2(new_n306), .A3(new_n685), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n281), .A2(new_n288), .A3(new_n302), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT37), .B1(new_n870), .B2(new_n342), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n329), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n328), .ZN(new_n873));
  INV_X1    g0673(.A(new_n685), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n873), .A2(new_n874), .B1(new_n340), .B2(new_n298), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n342), .A2(new_n288), .A3(new_n281), .A4(new_n302), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT37), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT105), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n874), .B1(new_n340), .B2(new_n298), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n347), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n872), .A2(KEYINPUT105), .A3(new_n878), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n881), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n881), .A2(new_n883), .A3(KEYINPUT38), .A4(new_n884), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(KEYINPUT106), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT108), .B1(new_n749), .B2(KEYINPUT31), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT108), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n745), .A2(new_n891), .A3(new_n746), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n730), .A2(new_n750), .A3(new_n890), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n388), .A2(new_n690), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n389), .A2(new_n393), .A3(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n388), .B(new_n690), .C1(new_n392), .C2(new_n373), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n834), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT106), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n885), .A2(new_n899), .A3(new_n886), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n889), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n329), .A2(new_n871), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT107), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n876), .A2(new_n904), .B1(new_n303), .B2(new_n328), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n870), .A2(KEYINPUT107), .A3(new_n342), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n869), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n903), .A2(new_n869), .B1(new_n907), .B2(KEYINPUT37), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n869), .B1(new_n671), .B2(new_n344), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n886), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n888), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n893), .A2(KEYINPUT40), .A3(new_n897), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n901), .A2(new_n902), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n469), .A2(new_n893), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n698), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n914), .B2(new_n915), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n917), .B(KEYINPUT109), .Z(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n889), .A2(KEYINPUT39), .A3(new_n900), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n911), .A2(KEYINPUT39), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n373), .A2(new_n388), .A3(new_n691), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n895), .A2(new_n896), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n666), .A2(new_n691), .A3(new_n862), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n926), .B1(new_n927), .B2(new_n833), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(new_n900), .A3(new_n889), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n672), .A2(new_n874), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n925), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n469), .B1(new_n718), .B2(new_n728), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n677), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n932), .B(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n868), .B1(new_n919), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n919), .B2(new_n935), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n234), .A2(new_n207), .A3(new_n569), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT36), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n266), .A2(new_n227), .A3(new_n375), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n214), .A2(G50), .ZN(new_n944));
  OAI211_X1 g0744(.A(G1), .B(new_n756), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n937), .A2(new_n942), .A3(new_n945), .ZN(G367));
  OAI21_X1  g0746(.A(new_n690), .B1(new_n509), .B2(new_n510), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n522), .A2(new_n947), .B1(new_n662), .B2(new_n690), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n948), .A2(new_n707), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT42), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n645), .B1(new_n948), .B2(new_n702), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n691), .ZN(new_n952));
  OR3_X1    g0752(.A1(new_n654), .A2(new_n561), .A3(new_n691), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n654), .B(new_n656), .C1(new_n561), .C2(new_n691), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n950), .A2(new_n952), .B1(KEYINPUT43), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n955), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n956), .B(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n704), .A2(new_n948), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n705), .A2(new_n707), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n948), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT44), .Z(new_n965));
  NOR2_X1   g0765(.A1(new_n948), .A2(new_n963), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT45), .ZN(new_n967));
  AND3_X1   g0767(.A1(new_n965), .A2(new_n704), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n704), .B1(new_n965), .B2(new_n967), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n707), .B1(new_n703), .B2(new_n706), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n699), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n753), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n710), .B(KEYINPUT41), .Z(new_n974));
  OAI21_X1  g0774(.A(new_n758), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n962), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n772), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n241), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n777), .B1(new_n210), .B2(new_n396), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n760), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n409), .B1(new_n781), .B2(new_n202), .C1(new_n846), .C2(new_n784), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n797), .B2(G137), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n811), .A2(G58), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n787), .A2(G159), .B1(new_n799), .B2(G143), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n800), .A2(new_n375), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G68), .B2(new_n820), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n982), .A2(new_n983), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT110), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT46), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n810), .A2(new_n989), .A3(new_n569), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n409), .B1(new_n838), .B2(new_n612), .ZN(new_n991));
  INV_X1    g0791(.A(G283), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n991), .B1(new_n992), .B2(new_n781), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G317), .B2(new_n797), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n989), .B1(new_n810), .B2(new_n569), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n848), .A2(new_n782), .B1(new_n408), .B2(new_n805), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n845), .A2(new_n803), .B1(new_n222), .B2(new_n800), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n994), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n988), .B1(new_n990), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT47), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n980), .B1(new_n1001), .B2(new_n776), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n957), .A2(new_n766), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n976), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(G387));
  OR2_X1    g0806(.A1(new_n703), .A2(new_n767), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n712), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n770), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(G107), .B2(new_n210), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n245), .A2(new_n308), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT111), .ZN(new_n1012));
  AOI211_X1 g0812(.A(G45), .B(new_n1008), .C1(G68), .C2(G77), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n289), .A2(G50), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT50), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n977), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1010), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n777), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n760), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n257), .B1(new_n801), .B2(G97), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n810), .B2(new_n375), .C1(new_n796), .C2(new_n846), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT112), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n805), .A2(new_n396), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n838), .A2(G50), .B1(new_n818), .B2(G68), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n289), .B2(new_n845), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1023), .B(new_n1025), .C1(G159), .C2(new_n799), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT113), .Z(new_n1028));
  OAI22_X1  g0828(.A1(new_n810), .A2(new_n803), .B1(new_n992), .B2(new_n805), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT114), .Z(new_n1030));
  AOI22_X1  g0830(.A1(new_n838), .A2(G317), .B1(new_n818), .B2(new_n612), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n845), .B2(new_n782), .C1(new_n783), .C2(new_n848), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT48), .ZN(new_n1033));
  AOI21_X1  g0833(.A(KEYINPUT49), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1030), .A2(new_n1033), .A3(KEYINPUT49), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n797), .A2(G326), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n409), .B1(new_n801), .B2(G116), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1028), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1019), .B1(new_n1039), .B2(new_n776), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n972), .A2(new_n759), .B1(new_n1007), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n754), .A2(new_n972), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n710), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n754), .A2(new_n972), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(G393));
  OR2_X1    g0845(.A1(new_n970), .A2(KEYINPUT115), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n970), .A2(KEYINPUT115), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(new_n1047), .A3(new_n759), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n970), .A2(new_n754), .A3(new_n972), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1042), .B1(new_n968), .B2(new_n969), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n710), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n948), .A2(new_n766), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n409), .B(new_n822), .C1(G294), .C2(new_n818), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G116), .A2(new_n820), .B1(new_n787), .B2(new_n612), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n992), .B2(new_n810), .C1(new_n783), .C2(new_n796), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G317), .A2(new_n799), .B1(new_n838), .B2(G311), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G150), .A2(new_n799), .B1(new_n838), .B2(G159), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT51), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n797), .A2(G143), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n811), .A2(G68), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n409), .B1(new_n781), .B2(new_n289), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G87), .B2(new_n801), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G77), .A2(new_n820), .B1(new_n787), .B2(G50), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1056), .A2(new_n1058), .B1(new_n1060), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n776), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1018), .B1(G97), .B2(new_n709), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n250), .A2(new_n772), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n769), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1052), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1048), .A2(new_n1051), .A3(new_n1072), .ZN(G390));
  OAI21_X1  g0873(.A(new_n760), .B1(new_n860), .B2(new_n293), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n845), .A2(new_n408), .B1(new_n848), .B2(new_n992), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n854), .B(new_n1075), .C1(G77), .C2(new_n820), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n797), .A2(G294), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n257), .B1(new_n784), .B2(new_n569), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G97), .B2(new_n818), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1076), .A2(new_n816), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(G128), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n845), .A2(new_n847), .B1(new_n848), .B2(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n805), .A2(new_n813), .B1(new_n800), .B2(new_n202), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n797), .A2(G125), .ZN(new_n1085));
  OAI21_X1  g0885(.A(KEYINPUT53), .B1(new_n810), .B2(new_n846), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(KEYINPUT54), .B(G143), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n781), .A2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n257), .B(new_n1088), .C1(G132), .C2(new_n838), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .A4(new_n1089), .ZN(new_n1090));
  NOR3_X1   g0890(.A1(new_n810), .A2(KEYINPUT53), .A3(new_n846), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1080), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1074), .B1(new_n1092), .B2(new_n776), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n922), .B2(new_n765), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n893), .A2(G330), .A3(new_n897), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n833), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n716), .B2(new_n862), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n923), .B1(new_n1097), .B2(new_n926), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n920), .A2(new_n1098), .A3(new_n921), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n888), .A2(new_n910), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1100), .A2(new_n924), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n727), .A2(new_n691), .A3(new_n832), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1102), .A2(new_n833), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1101), .B1(new_n1103), .B2(new_n926), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1095), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n751), .A2(G330), .A3(new_n862), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1108), .A2(new_n926), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1105), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1094), .B1(new_n1111), .B2(new_n758), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n469), .A2(G330), .A3(new_n893), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n677), .A2(new_n933), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n893), .A2(G330), .A3(new_n862), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n926), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1103), .A2(new_n1109), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1097), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1108), .A2(new_n926), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1095), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1115), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n711), .B1(new_n1111), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1114), .B1(new_n1122), .B2(new_n1118), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1099), .A2(new_n1104), .A3(new_n1109), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1126), .B(new_n1127), .C1(new_n1107), .C2(new_n1095), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1112), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(G378));
  INV_X1    g0930(.A(KEYINPUT119), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n460), .A2(new_n464), .A3(new_n468), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n444), .A2(new_n685), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n460), .A2(new_n464), .A3(new_n468), .A4(new_n1133), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1137), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(G330), .B1(new_n1100), .B2(new_n912), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1140), .B(new_n1141), .C1(new_n902), .C2(new_n901), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1140), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n901), .A2(new_n902), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1141), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n932), .A2(new_n1142), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n923), .B1(new_n920), .B2(new_n921), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n929), .A2(new_n930), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n1140), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1144), .A2(new_n1145), .A3(new_n1143), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1150), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT57), .B1(new_n1147), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1114), .B1(new_n1110), .B2(new_n1123), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1131), .B(new_n710), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n932), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1152), .A2(new_n1150), .A3(new_n1153), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT118), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1158), .A2(new_n1159), .A3(KEYINPUT118), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1156), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1157), .B1(new_n1164), .B2(KEYINPUT57), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1128), .A2(new_n1115), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(KEYINPUT57), .A3(new_n1160), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1131), .B1(new_n1167), .B2(new_n710), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n760), .B1(new_n860), .B2(G50), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1143), .A2(new_n765), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n799), .A2(G116), .B1(new_n801), .B2(G58), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n214), .B2(new_n805), .C1(new_n222), .C2(new_n845), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n257), .A2(new_n307), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n838), .B2(G107), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n396), .B2(new_n781), .C1(new_n796), .C2(new_n992), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1173), .B(new_n1176), .C1(G77), .C2(new_n811), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT58), .Z(new_n1178));
  OAI211_X1 g0978(.A(new_n1174), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n784), .A2(new_n1081), .B1(new_n781), .B2(new_n847), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G132), .B2(new_n787), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G150), .A2(new_n820), .B1(new_n799), .B2(G125), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n810), .C2(new_n1087), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n797), .A2(G124), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G33), .B(G41), .C1(new_n801), .C2(G159), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1178), .B(new_n1179), .C1(new_n1184), .C2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT116), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n826), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1170), .B(new_n1171), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT117), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1195), .B2(new_n759), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1169), .A2(new_n1196), .ZN(G375));
  NAND2_X1  g0997(.A1(new_n926), .A2(new_n764), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n760), .B1(new_n860), .B2(G68), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n799), .A2(G132), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n220), .B2(new_n800), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n796), .A2(new_n1081), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n845), .A2(new_n1087), .B1(new_n202), .B2(new_n805), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n409), .B1(new_n781), .B2(new_n846), .C1(new_n847), .C2(new_n784), .ZN(new_n1204));
  OR4_X1    g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n810), .A2(new_n813), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1023), .B1(G283), .B2(new_n838), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT120), .Z(new_n1208));
  NAND2_X1  g1008(.A1(new_n797), .A2(G303), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n811), .A2(G97), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n409), .B(new_n985), .C1(G107), .C2(new_n818), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n787), .A2(G116), .B1(new_n799), .B2(G294), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n1205), .A2(new_n1206), .B1(new_n1208), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1199), .B1(new_n1214), .B2(new_n776), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1123), .A2(new_n759), .B1(new_n1198), .B2(new_n1215), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1126), .A2(new_n974), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1115), .A2(new_n1123), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(G381));
  NAND3_X1  g1019(.A1(new_n1169), .A2(new_n1129), .A3(new_n1196), .ZN(new_n1220));
  OR4_X1    g1020(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1221));
  OR4_X1    g1021(.A1(G387), .A2(new_n1220), .A3(new_n1221), .A4(G381), .ZN(G407));
  OAI211_X1 g1022(.A(G407), .B(G213), .C1(new_n689), .C2(new_n1220), .ZN(G409));
  NAND3_X1  g1023(.A1(new_n687), .A2(new_n688), .A3(G213), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(G378), .B(new_n1196), .C1(new_n1165), .C2(new_n1168), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1193), .B1(new_n1160), .B2(new_n759), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1195), .A2(new_n1166), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n974), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n1129), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1225), .B1(new_n1226), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1216), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1124), .A2(KEYINPUT60), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1233), .A2(new_n1218), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n711), .B1(new_n1233), .B2(new_n1218), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1232), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT121), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n866), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n866), .B(KEYINPUT121), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1239), .B1(new_n1236), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1231), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT122), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT63), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1231), .A2(KEYINPUT122), .A3(new_n1242), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT61), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1225), .A2(G2897), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1241), .B(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1249), .B1(new_n1251), .B2(new_n1231), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1005), .A2(G390), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1005), .A2(G390), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(G393), .B(G396), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT123), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1258), .A2(KEYINPUT123), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1257), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1254), .A2(KEYINPUT124), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1258), .B1(new_n1254), .B2(KEYINPUT124), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1256), .B(KEYINPUT125), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1261), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1231), .A2(KEYINPUT63), .A3(new_n1242), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1248), .A2(new_n1253), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1226), .A2(new_n1230), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1269), .A2(KEYINPUT62), .A3(new_n1224), .A4(new_n1242), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(KEYINPUT126), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT126), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1231), .A2(new_n1272), .A3(KEYINPUT62), .A4(new_n1242), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT62), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1245), .A2(new_n1275), .A3(new_n1247), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1252), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1268), .B1(new_n1277), .B2(new_n1266), .ZN(G405));
  AOI21_X1  g1078(.A(G378), .B1(new_n1169), .B2(new_n1196), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1226), .ZN(new_n1280));
  OR3_X1    g1080(.A1(new_n1279), .A2(new_n1280), .A3(new_n1242), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1242), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  XOR2_X1   g1083(.A(new_n1283), .B(new_n1266), .Z(G402));
endmodule


