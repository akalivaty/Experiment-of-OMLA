//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT87), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G128), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(G125), .B1(new_n191), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n199), .B1(new_n189), .B2(G146), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n192), .A2(KEYINPUT64), .A3(G143), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n193), .B(new_n198), .C1(new_n200), .C2(new_n201), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n196), .A2(KEYINPUT84), .A3(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT84), .B1(new_n196), .B2(new_n202), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n193), .B(new_n207), .C1(new_n200), .C2(new_n201), .ZN(new_n208));
  OR2_X1    g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n195), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n205), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n203), .A2(new_n204), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G953), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G224), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT7), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT85), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g031(.A1(KEYINPUT79), .A2(G107), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT79), .A2(G107), .ZN(new_n219));
  AOI21_X1  g033(.A(G104), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G104), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT80), .B1(new_n221), .B2(G107), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n223));
  INV_X1    g037(.A(G107), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(G104), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(G101), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n224), .A2(G104), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G101), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n224), .A2(G104), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT3), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n218), .A2(new_n219), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n229), .B(new_n231), .C1(new_n232), .C2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n227), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G116), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G119), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT5), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G116), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(G119), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n240), .B(G113), .C1(new_n244), .C2(new_n239), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT2), .B(G113), .Z(new_n246));
  XNOR2_X1  g060(.A(G116), .B(G119), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n236), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n227), .A2(new_n235), .A3(new_n245), .A4(new_n248), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G110), .B(G122), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT8), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n211), .B1(new_n202), .B2(new_n196), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n252), .A2(new_n254), .B1(new_n255), .B2(new_n216), .ZN(new_n256));
  INV_X1    g070(.A(G101), .ZN(new_n257));
  INV_X1    g071(.A(new_n219), .ZN(new_n258));
  NOR2_X1   g072(.A1(KEYINPUT79), .A2(G107), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n260), .A2(new_n233), .B1(KEYINPUT3), .B2(new_n230), .ZN(new_n261));
  INV_X1    g075(.A(new_n228), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n235), .A2(KEYINPUT4), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n231), .B1(new_n232), .B2(new_n234), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n266), .B(G101), .C1(new_n267), .C2(new_n228), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT2), .B(G113), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n244), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n248), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n251), .B(new_n253), .C1(new_n265), .C2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT85), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n196), .A2(new_n202), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT84), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n208), .A2(new_n210), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G125), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n274), .B(new_n215), .C1(new_n280), .C2(new_n203), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n217), .A2(new_n256), .A3(new_n273), .A4(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT86), .ZN(new_n283));
  INV_X1    g097(.A(G902), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n251), .B1(new_n265), .B2(new_n272), .ZN(new_n286));
  INV_X1    g100(.A(new_n253), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(KEYINPUT6), .A3(new_n273), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n286), .A2(new_n290), .A3(new_n287), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n255), .B(new_n214), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n285), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n283), .B1(new_n282), .B2(new_n284), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n188), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G210), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n282), .A2(new_n284), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT86), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n300), .A2(KEYINPUT87), .A3(new_n293), .A4(new_n285), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n296), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n300), .A2(new_n297), .A3(new_n293), .A4(new_n285), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT9), .B(G234), .ZN(new_n305));
  OAI21_X1  g119(.A(G221), .B1(new_n305), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G469), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(new_n284), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n191), .A2(new_n195), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n202), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT82), .B1(new_n312), .B2(new_n236), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n227), .A2(new_n235), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT82), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT10), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(new_n202), .B2(new_n310), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G137), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT66), .B1(new_n320), .B2(G134), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT66), .ZN(new_n322));
  INV_X1    g136(.A(G134), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(G137), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT65), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n323), .B2(G137), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT11), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n320), .A2(G134), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT11), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n325), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G131), .ZN(new_n333));
  INV_X1    g147(.A(G131), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n325), .A2(new_n328), .A3(new_n334), .A4(new_n331), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT1), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(G143), .B2(new_n192), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n197), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n190), .A2(KEYINPUT81), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT64), .B1(new_n192), .B2(G143), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n199), .A2(new_n189), .A3(G146), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n341), .A2(new_n342), .B1(new_n193), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n202), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n316), .B1(new_n348), .B2(new_n236), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n208), .A2(new_n210), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n268), .B(new_n350), .C1(new_n263), .C2(new_n264), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n319), .A2(new_n337), .A3(new_n349), .A4(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT83), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(new_n314), .B2(new_n311), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n314), .B1(new_n347), .B2(new_n346), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n236), .A2(KEYINPUT83), .A3(new_n202), .A4(new_n310), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n357), .A2(KEYINPUT12), .A3(new_n336), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT12), .B1(new_n357), .B2(new_n336), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n352), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(G110), .B(G140), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n213), .A2(G227), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n361), .B(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT78), .ZN(new_n364));
  INV_X1    g178(.A(new_n363), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n352), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n312), .A2(new_n236), .A3(KEYINPUT82), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n315), .B1(new_n314), .B2(new_n317), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n349), .B(new_n351), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n336), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n360), .A2(new_n364), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n309), .B1(new_n372), .B2(G469), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n357), .A2(KEYINPUT12), .A3(new_n336), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n357), .A2(new_n336), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT12), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n366), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n365), .B1(new_n371), .B2(new_n352), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n308), .B(new_n284), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n307), .B1(new_n373), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(G237), .A2(G953), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(G143), .A3(G214), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(G143), .B1(new_n382), .B2(G214), .ZN(new_n385));
  OAI211_X1 g199(.A(KEYINPUT18), .B(G131), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(G214), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n189), .ZN(new_n388));
  NAND2_X1  g202(.A1(KEYINPUT18), .A2(G131), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n383), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G125), .B(G140), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n391), .A2(new_n192), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n192), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n386), .B(new_n390), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n384), .A2(new_n385), .A3(G131), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n334), .B1(new_n388), .B2(new_n383), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT17), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(new_n391), .B2(KEYINPUT16), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G146), .ZN(new_n400));
  OAI211_X1 g214(.A(KEYINPUT17), .B(G131), .C1(new_n384), .C2(new_n385), .ZN(new_n401));
  INV_X1    g215(.A(G140), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G125), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n205), .A2(G140), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT16), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n192), .B1(new_n405), .B2(new_n398), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n400), .A2(new_n401), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n394), .B1(new_n397), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G113), .B(G122), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(new_n221), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n410), .B(new_n394), .C1(new_n397), .C2(new_n407), .ZN(new_n413));
  AOI21_X1  g227(.A(G902), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT89), .B(G475), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT19), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT19), .B1(new_n403), .B2(new_n404), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n192), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n400), .B(new_n421), .C1(new_n395), .C2(new_n396), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n394), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n411), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n424), .A2(new_n413), .A3(KEYINPUT88), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT88), .B1(new_n424), .B2(new_n413), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(G475), .A2(G902), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n418), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n424), .A2(new_n413), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n430), .A2(new_n418), .A3(new_n428), .ZN(new_n431));
  OAI211_X1 g245(.A(KEYINPUT90), .B(new_n417), .C1(new_n429), .C2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT90), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n424), .A2(new_n413), .A3(KEYINPUT88), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n428), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n431), .B1(new_n437), .B2(KEYINPUT20), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n433), .B1(new_n438), .B2(new_n416), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n189), .A2(G128), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT13), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n441), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n197), .A2(G143), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT92), .A4(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT92), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n323), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n440), .A2(new_n445), .A3(new_n323), .ZN(new_n450));
  INV_X1    g264(.A(G122), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G116), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n237), .A2(G122), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n454), .B1(new_n452), .B2(new_n453), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n456), .A2(new_n260), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n457), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n232), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n449), .B(new_n450), .C1(new_n458), .C2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n460), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n440), .A2(new_n445), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G134), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n450), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n237), .A2(KEYINPUT14), .A3(G122), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n452), .A2(new_n453), .ZN(new_n467));
  OAI211_X1 g281(.A(G107), .B(new_n466), .C1(new_n467), .C2(KEYINPUT14), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n462), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G217), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n305), .A2(new_n470), .A3(G953), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n461), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n471), .B1(new_n461), .B2(new_n469), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n284), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G478), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(KEYINPUT15), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OAI221_X1 g291(.A(new_n284), .B1(KEYINPUT15), .B2(new_n475), .C1(new_n472), .C2(new_n473), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT21), .B(G898), .ZN(new_n480));
  NAND2_X1  g294(.A1(G234), .A2(G237), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n480), .A2(G902), .A3(G953), .A4(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(KEYINPUT93), .A2(G952), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(KEYINPUT93), .A2(G952), .ZN(new_n485));
  AOI21_X1  g299(.A(G953), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n481), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n479), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n432), .A2(new_n439), .A3(new_n488), .ZN(new_n489));
  AND4_X1   g303(.A1(new_n187), .A2(new_n304), .A3(new_n381), .A4(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(G472), .A2(G902), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT32), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n382), .A2(G210), .ZN(new_n495));
  XOR2_X1   g309(.A(new_n495), .B(KEYINPUT70), .Z(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT26), .B(G101), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n496), .B(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT67), .ZN(new_n502));
  AOI211_X1 g316(.A(new_n502), .B(new_n278), .C1(new_n335), .C2(new_n333), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT67), .B1(new_n336), .B2(new_n350), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT68), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n246), .A2(new_n247), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n244), .A2(new_n269), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n248), .A2(KEYINPUT68), .A3(new_n270), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n323), .A2(G137), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n329), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G131), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n311), .A2(new_n335), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n503), .A2(new_n504), .A3(new_n515), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n202), .A2(new_n310), .B1(G131), .B2(new_n512), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n336), .A2(new_n350), .B1(new_n335), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n271), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT28), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT73), .ZN(new_n522));
  INV_X1    g336(.A(new_n514), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n278), .B1(new_n333), .B2(new_n335), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n330), .B1(new_n329), .B2(new_n326), .ZN(new_n526));
  AOI211_X1 g340(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n320), .C2(G134), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n334), .B1(new_n528), .B2(new_n325), .ZN(new_n529));
  INV_X1    g343(.A(new_n335), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n350), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT73), .A3(new_n514), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n525), .A2(new_n532), .A3(new_n510), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT28), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n501), .B1(new_n521), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n503), .A2(new_n504), .ZN(new_n537));
  INV_X1    g351(.A(new_n515), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n500), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n531), .A2(new_n514), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n519), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n531), .A2(new_n502), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n524), .A2(KEYINPUT67), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n541), .B1(new_n517), .B2(new_n335), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g361(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n548));
  AND3_X1   g362(.A1(new_n539), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n536), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT71), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n514), .A2(KEYINPUT30), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n503), .A2(new_n504), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n271), .B1(new_n518), .B2(KEYINPUT30), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n538), .A2(new_n543), .A3(new_n544), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n501), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n551), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n539), .A2(new_n547), .A3(KEYINPUT71), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(KEYINPUT31), .A3(new_n559), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n550), .A2(KEYINPUT74), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT74), .B1(new_n550), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n494), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n510), .B1(new_n537), .B2(new_n514), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT28), .B1(new_n564), .B2(new_n516), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT29), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n500), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n535), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT75), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT75), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n565), .A2(new_n570), .A3(new_n535), .A4(new_n567), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n547), .A2(new_n556), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n500), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n521), .A2(new_n501), .A3(new_n535), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n574), .A3(new_n566), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n569), .A2(new_n284), .A3(new_n571), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G472), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT74), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n539), .A2(new_n547), .A3(KEYINPUT71), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT71), .B1(new_n539), .B2(new_n547), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT31), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n533), .A2(new_n534), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n540), .A2(new_n271), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n534), .B1(new_n556), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n500), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n539), .A2(new_n547), .A3(new_n548), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n578), .B1(new_n582), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n550), .A2(KEYINPUT74), .A3(new_n560), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n492), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n563), .B(new_n577), .C1(new_n591), .C2(KEYINPUT32), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n470), .B1(G234), .B2(new_n284), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n400), .A2(new_n406), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n241), .A2(G128), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n197), .A2(G119), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n596), .B(new_n597), .C1(new_n599), .C2(KEYINPUT23), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G110), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n596), .A2(new_n598), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT24), .B(G110), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n595), .B(new_n601), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n392), .B1(new_n399), .B2(G146), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT76), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n602), .A2(new_n603), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(new_n600), .B2(G110), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n606), .B1(new_n605), .B2(new_n608), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n604), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT22), .B(G137), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n213), .A2(G221), .A3(G234), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n604), .B(new_n614), .C1(new_n609), .C2(new_n610), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n284), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT25), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n616), .A2(KEYINPUT25), .A3(new_n284), .A4(new_n617), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n594), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n593), .A2(G902), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n616), .A2(new_n617), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT77), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n490), .A2(new_n592), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G101), .ZN(G3));
  OAI21_X1  g444(.A(new_n284), .B1(new_n561), .B2(new_n562), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n591), .B1(G472), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n360), .A2(new_n364), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n367), .A2(new_n371), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(G469), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n309), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n380), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n306), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n627), .A2(new_n638), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n472), .A2(new_n473), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT33), .ZN(new_n641));
  OR3_X1    g455(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT33), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(G478), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n640), .A2(new_n475), .A3(new_n284), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n475), .A2(new_n284), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n432), .B2(new_n439), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n487), .A2(new_n482), .ZN(new_n649));
  INV_X1    g463(.A(new_n187), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n298), .B1(new_n294), .B2(new_n295), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n650), .B1(new_n651), .B2(new_n303), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n648), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n632), .A2(new_n639), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  XOR2_X1   g470(.A(new_n649), .B(KEYINPUT94), .Z(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n416), .A2(new_n658), .ZN(new_n659));
  AND4_X1   g473(.A1(new_n418), .A2(new_n435), .A3(new_n428), .A4(new_n436), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n479), .B(new_n659), .C1(new_n429), .C2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT95), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n651), .A2(new_n303), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n427), .A2(new_n418), .A3(new_n428), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n437), .A2(KEYINPUT20), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT95), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n666), .A2(new_n667), .A3(new_n479), .A4(new_n659), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n662), .A2(new_n663), .A3(new_n187), .A4(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT96), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n652), .A2(KEYINPUT96), .A3(new_n662), .A4(new_n668), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n632), .A3(new_n639), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT35), .B(G107), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  OR2_X1    g490(.A1(new_n615), .A2(KEYINPUT36), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n611), .B(new_n677), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n678), .A2(G902), .A3(new_n593), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n622), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n490), .A2(new_n632), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT37), .B(G110), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G12));
  AND3_X1   g498(.A1(new_n381), .A2(new_n652), .A3(new_n681), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n481), .A2(G902), .A3(G953), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n487), .B1(G900), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT97), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n688), .B1(new_n414), .B2(new_n415), .ZN(new_n689));
  INV_X1    g503(.A(new_n479), .ZN(new_n690));
  AOI211_X1 g504(.A(new_n689), .B(new_n690), .C1(new_n665), .C2(new_n664), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n592), .A2(new_n685), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  NOR2_X1   g507(.A1(new_n579), .A2(new_n580), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n500), .B1(new_n564), .B2(new_n516), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT98), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n558), .A2(KEYINPUT98), .A3(new_n695), .A4(new_n559), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n284), .ZN(new_n698));
  OAI21_X1  g512(.A(G472), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n563), .B(new_n699), .C1(new_n591), .C2(KEYINPUT32), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT99), .Z(new_n701));
  XOR2_X1   g515(.A(new_n304), .B(KEYINPUT38), .Z(new_n702));
  NAND2_X1  g516(.A1(new_n432), .A2(new_n439), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(new_n187), .A3(new_n479), .A4(new_n680), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n688), .B(KEYINPUT39), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n381), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n704), .B1(new_n706), .B2(KEYINPUT40), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(KEYINPUT40), .B2(new_n706), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n701), .A2(new_n702), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n189), .ZN(G45));
  NAND2_X1  g524(.A1(new_n648), .A2(new_n688), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n592), .A2(new_n685), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  NAND2_X1  g528(.A1(new_n377), .A2(new_n374), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n371), .A2(new_n352), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n715), .A2(new_n367), .B1(new_n716), .B2(new_n363), .ZN(new_n717));
  OAI21_X1  g531(.A(G469), .B1(new_n717), .B2(G902), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n306), .A3(new_n380), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT100), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT100), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n718), .A2(new_n721), .A3(new_n306), .A4(new_n380), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n592), .A3(new_n628), .A4(new_n653), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND4_X1  g540(.A1(new_n673), .A2(new_n592), .A3(new_n723), .A4(new_n628), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  AND3_X1   g542(.A1(new_n720), .A2(new_n652), .A3(new_n722), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n489), .A2(new_n681), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n592), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G119), .ZN(G21));
  AND3_X1   g546(.A1(new_n720), .A2(new_n657), .A3(new_n722), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n543), .A2(new_n544), .A3(new_n514), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n509), .A3(new_n508), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n534), .B1(new_n735), .B2(new_n556), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n500), .B1(new_n736), .B2(new_n583), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n560), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT101), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n560), .A2(new_n737), .A3(KEYINPUT101), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n587), .A3(new_n741), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n631), .A2(G472), .B1(new_n742), .B2(new_n491), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n652), .A2(new_n703), .A3(new_n479), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n733), .A2(new_n743), .A3(new_n626), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G122), .ZN(G24));
  NAND4_X1  g560(.A1(new_n729), .A2(new_n743), .A3(new_n681), .A4(new_n712), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  AND2_X1   g562(.A1(new_n303), .A2(new_n187), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n302), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n638), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n592), .A2(new_n628), .A3(new_n712), .A4(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n753));
  INV_X1    g567(.A(new_n626), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n589), .A2(new_n590), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n755), .A2(new_n494), .B1(G472), .B2(new_n576), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n491), .B1(new_n561), .B2(new_n562), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n493), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n754), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  NOR4_X1   g574(.A1(new_n711), .A2(new_n750), .A3(new_n638), .A4(new_n760), .ZN(new_n761));
  AOI22_X1  g575(.A1(new_n752), .A2(new_n753), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n334), .ZN(G33));
  NAND4_X1  g577(.A1(new_n592), .A2(new_n628), .A3(new_n691), .A4(new_n751), .ZN(new_n764));
  XOR2_X1   g578(.A(KEYINPUT103), .B(G134), .Z(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G36));
  OAI21_X1  g580(.A(G469), .B1(new_n372), .B2(KEYINPUT45), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(KEYINPUT45), .B2(new_n372), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n768), .A2(new_n309), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT46), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(new_n380), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n769), .A2(new_n770), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n307), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n705), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT104), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n703), .B(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n647), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(KEYINPUT43), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n703), .A2(new_n647), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n780), .B1(KEYINPUT43), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n632), .A2(new_n680), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n775), .B1(new_n776), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT105), .ZN(new_n786));
  INV_X1    g600(.A(new_n750), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n787), .B1(new_n784), .B2(new_n776), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n785), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n788), .A2(new_n786), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n320), .ZN(G39));
  NAND2_X1  g606(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n774), .A2(new_n793), .ZN(new_n794));
  XOR2_X1   g608(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n795));
  OAI21_X1  g609(.A(new_n794), .B1(new_n774), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n712), .A2(new_n627), .A3(new_n787), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n796), .A2(new_n592), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n402), .ZN(G42));
  NAND2_X1  g613(.A1(new_n718), .A2(new_n380), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n800), .A2(KEYINPUT49), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(KEYINPUT49), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n779), .A2(new_n626), .A3(new_n187), .A4(new_n306), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n701), .A2(new_n702), .A3(new_n778), .A4(new_n804), .ZN(new_n805));
  XOR2_X1   g619(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n806));
  OAI211_X1 g620(.A(new_n592), .B(new_n685), .C1(new_n691), .C2(new_n712), .ZN(new_n807));
  INV_X1    g621(.A(new_n688), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n622), .A2(new_n679), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n637), .A2(new_n306), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(KEYINPUT110), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT110), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n381), .B2(new_n809), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n700), .B(new_n744), .C1(new_n811), .C2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n747), .A2(new_n807), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT52), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n747), .A2(new_n807), .A3(new_n814), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n816), .A2(KEYINPUT111), .A3(new_n818), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n745), .A2(new_n731), .A3(new_n629), .A4(new_n682), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT107), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n825), .B1(new_n703), .B2(new_n690), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n703), .A2(new_n779), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n432), .A2(new_n439), .A3(KEYINPUT107), .A4(new_n479), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n650), .B(new_n658), .C1(new_n302), .C2(new_n303), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n632), .A2(new_n639), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n727), .A2(new_n724), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n824), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n762), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n631), .A2(G472), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n742), .A2(new_n491), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(new_n681), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n751), .A2(new_n712), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT109), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n711), .A2(new_n750), .A3(new_n638), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT109), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n743), .A3(new_n841), .A4(new_n681), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT108), .ZN(new_n844));
  AOI211_X1 g658(.A(new_n689), .B(new_n479), .C1(new_n664), .C2(new_n665), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n637), .A2(new_n681), .A3(new_n845), .A4(new_n306), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n750), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n592), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n844), .B1(new_n592), .B2(new_n847), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n764), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n833), .A2(new_n834), .A3(new_n843), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n823), .A2(new_n853), .A3(KEYINPUT53), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  OAI211_X1 g669(.A(KEYINPUT112), .B(new_n855), .C1(new_n852), .C2(new_n819), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n839), .A2(new_n842), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n858), .A2(new_n850), .A3(new_n762), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n833), .A3(new_n818), .A4(new_n816), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT112), .B1(new_n860), .B2(new_n855), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n806), .B(new_n854), .C1(new_n857), .C2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT53), .B1(new_n823), .B2(new_n853), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n860), .A2(new_n855), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT54), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT114), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n862), .A2(new_n865), .A3(KEYINPUT114), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n796), .B1(new_n306), .B2(new_n800), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n743), .A2(new_n626), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n782), .A2(new_n481), .A3(new_n486), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n872), .A2(new_n873), .A3(new_n787), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n873), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n702), .A2(new_n650), .A3(new_n723), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n876), .A2(KEYINPUT50), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n723), .A2(new_n787), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT115), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(new_n837), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT50), .B1(new_n876), .B2(new_n877), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n875), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n627), .A2(new_n487), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n880), .A2(new_n701), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n703), .A2(new_n779), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n871), .B1(new_n885), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n889), .A2(new_n648), .A3(new_n890), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n874), .A2(new_n880), .A3(new_n759), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT48), .Z(new_n897));
  XNOR2_X1  g711(.A(new_n486), .B(KEYINPUT117), .ZN(new_n898));
  INV_X1    g712(.A(new_n729), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n898), .B1(new_n876), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n894), .A2(new_n895), .A3(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n885), .A2(new_n871), .A3(new_n893), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n870), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(G952), .A2(G953), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n805), .B1(new_n904), .B2(new_n905), .ZN(G75));
  NOR2_X1   g720(.A1(new_n213), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n854), .B1(new_n857), .B2(new_n861), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(G902), .ZN(new_n910));
  INV_X1    g724(.A(G210), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n289), .A2(new_n291), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n292), .ZN(new_n914));
  XNOR2_X1  g728(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n910), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n909), .A2(KEYINPUT119), .A3(G902), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n298), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n916), .A2(KEYINPUT56), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n907), .B(new_n917), .C1(new_n921), .C2(new_n922), .ZN(G51));
  INV_X1    g737(.A(new_n806), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n909), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n926), .A3(new_n862), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n909), .A2(KEYINPUT120), .A3(new_n924), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n309), .B(KEYINPUT57), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n378), .B2(new_n379), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n919), .A2(new_n768), .A3(new_n920), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n907), .B1(new_n931), .B2(new_n932), .ZN(G54));
  NAND4_X1  g747(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .A4(new_n920), .ZN(new_n934));
  INV_X1    g748(.A(new_n427), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n907), .ZN(G60));
  AND2_X1   g752(.A1(new_n641), .A2(new_n642), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  XNOR2_X1  g754(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n646), .B(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n940), .B1(new_n870), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n939), .A2(new_n942), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n927), .A2(new_n928), .A3(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n907), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT122), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n862), .A2(KEYINPUT114), .A3(new_n865), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT114), .B1(new_n862), .B2(new_n865), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n943), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n939), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT122), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n953), .A2(new_n954), .A3(new_n947), .A4(new_n946), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n949), .A2(new_n955), .ZN(G63));
  NAND2_X1  g770(.A1(G217), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT60), .Z(new_n958));
  NAND2_X1  g772(.A1(new_n909), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n616), .A2(new_n617), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT124), .Z(new_n961));
  AOI21_X1  g775(.A(new_n907), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT61), .B1(new_n962), .B2(KEYINPUT123), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n962), .B1(new_n678), .B2(new_n959), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(G66));
  INV_X1    g779(.A(G224), .ZN(new_n966));
  OAI21_X1  g780(.A(G953), .B1(new_n480), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT125), .Z(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n833), .B2(G953), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT126), .Z(new_n970));
  INV_X1    g784(.A(G898), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n913), .B1(new_n971), .B2(G953), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n970), .B(new_n972), .ZN(G69));
  OAI21_X1  g787(.A(new_n546), .B1(KEYINPUT30), .B2(new_n518), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n419), .A2(new_n420), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(G900), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n976), .B1(new_n977), .B2(new_n213), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n791), .A2(new_n798), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n774), .A2(new_n705), .A3(new_n744), .A4(new_n759), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n747), .A2(new_n807), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n980), .A2(new_n834), .A3(new_n764), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n978), .B1(new_n984), .B2(new_n213), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n213), .B1(G227), .B2(G900), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n791), .A2(new_n798), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n709), .A2(new_n981), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT62), .Z(new_n989));
  NAND3_X1  g803(.A1(new_n592), .A2(new_n628), .A3(new_n751), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n829), .A2(new_n705), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n987), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n976), .B1(new_n994), .B2(new_n213), .ZN(new_n995));
  OR3_X1    g809(.A1(new_n985), .A2(new_n986), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n986), .B1(new_n985), .B2(new_n995), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(G72));
  XOR2_X1   g812(.A(new_n572), .B(KEYINPUT127), .Z(new_n999));
  NOR2_X1   g813(.A1(new_n999), .A2(new_n501), .ZN(new_n1000));
  NOR4_X1   g814(.A1(new_n979), .A2(new_n824), .A3(new_n832), .A4(new_n983), .ZN(new_n1001));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1000), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1004), .B1(new_n694), .B2(new_n573), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1006), .B1(new_n863), .B2(new_n864), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n987), .A2(new_n993), .A3(new_n833), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n501), .B(new_n999), .C1(new_n1008), .C2(new_n1004), .ZN(new_n1009));
  AND4_X1   g823(.A1(new_n947), .A2(new_n1005), .A3(new_n1007), .A4(new_n1009), .ZN(G57));
endmodule


