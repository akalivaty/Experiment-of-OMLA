

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U321 ( .A(n377), .B(n376), .ZN(n543) );
  XNOR2_X1 U322 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n376) );
  XOR2_X1 U323 ( .A(n326), .B(n325), .Z(n289) );
  XNOR2_X1 U324 ( .A(n336), .B(n321), .ZN(n322) );
  XNOR2_X1 U325 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U326 ( .A(n327), .B(n289), .ZN(n328) );
  XNOR2_X1 U327 ( .A(n329), .B(n328), .ZN(n369) );
  XNOR2_X1 U328 ( .A(n455), .B(G183GAT), .ZN(n456) );
  XNOR2_X1 U329 ( .A(n457), .B(n456), .ZN(G1350GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n291) );
  XNOR2_X1 U331 ( .A(G57GAT), .B(G64GAT), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n291), .B(n290), .ZN(n306) );
  XOR2_X1 U333 ( .A(G1GAT), .B(G127GAT), .Z(n406) );
  XOR2_X1 U334 ( .A(G78GAT), .B(G211GAT), .Z(n293) );
  XNOR2_X1 U335 ( .A(G183GAT), .B(G155GAT), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U337 ( .A(n406), .B(n294), .Z(n296) );
  NAND2_X1 U338 ( .A1(G231GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U340 ( .A(KEYINPUT81), .B(KEYINPUT15), .Z(n298) );
  XNOR2_X1 U341 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U343 ( .A(n300), .B(n299), .Z(n304) );
  XNOR2_X1 U344 ( .A(G15GAT), .B(G22GAT), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n301), .B(G8GAT), .ZN(n362) );
  XNOR2_X1 U346 ( .A(G71GAT), .B(KEYINPUT74), .ZN(n302) );
  XNOR2_X1 U347 ( .A(n302), .B(KEYINPUT13), .ZN(n333) );
  XNOR2_X1 U348 ( .A(n362), .B(n333), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U350 ( .A(n306), .B(n305), .Z(n477) );
  INV_X1 U351 ( .A(n477), .ZN(n577) );
  INV_X1 U352 ( .A(G50GAT), .ZN(n307) );
  NAND2_X1 U353 ( .A1(n307), .A2(G43GAT), .ZN(n310) );
  INV_X1 U354 ( .A(G43GAT), .ZN(n308) );
  NAND2_X1 U355 ( .A1(n308), .A2(G50GAT), .ZN(n309) );
  NAND2_X1 U356 ( .A1(n310), .A2(n309), .ZN(n312) );
  XNOR2_X1 U357 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n363) );
  INV_X1 U359 ( .A(n363), .ZN(n313) );
  XOR2_X1 U360 ( .A(G36GAT), .B(G190GAT), .Z(n388) );
  NAND2_X1 U361 ( .A1(n313), .A2(n388), .ZN(n316) );
  INV_X1 U362 ( .A(n388), .ZN(n314) );
  NAND2_X1 U363 ( .A1(n314), .A2(n363), .ZN(n315) );
  NAND2_X1 U364 ( .A1(n316), .A2(n315), .ZN(n318) );
  NAND2_X1 U365 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n323) );
  XOR2_X1 U367 ( .A(G92GAT), .B(KEYINPUT76), .Z(n320) );
  XNOR2_X1 U368 ( .A(G99GAT), .B(G85GAT), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n320), .B(n319), .ZN(n336) );
  XOR2_X1 U370 ( .A(KEYINPUT10), .B(KEYINPUT80), .Z(n321) );
  XOR2_X1 U371 ( .A(KEYINPUT9), .B(n324), .Z(n329) );
  XOR2_X1 U372 ( .A(G29GAT), .B(G134GAT), .Z(n408) );
  XNOR2_X1 U373 ( .A(G218GAT), .B(n408), .ZN(n327) );
  XOR2_X1 U374 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n326) );
  XNOR2_X1 U375 ( .A(G162GAT), .B(G106GAT), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n369), .B(KEYINPUT36), .ZN(n580) );
  NOR2_X1 U377 ( .A1(n577), .A2(n580), .ZN(n330) );
  XNOR2_X1 U378 ( .A(KEYINPUT45), .B(n330), .ZN(n367) );
  XOR2_X1 U379 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n332) );
  XNOR2_X1 U380 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n331) );
  XOR2_X1 U381 ( .A(n332), .B(n331), .Z(n346) );
  XOR2_X1 U382 ( .A(G176GAT), .B(G64GAT), .Z(n389) );
  XOR2_X1 U383 ( .A(n389), .B(KEYINPUT77), .Z(n335) );
  XNOR2_X1 U384 ( .A(n333), .B(KEYINPUT75), .ZN(n334) );
  XNOR2_X1 U385 ( .A(n335), .B(n334), .ZN(n340) );
  XOR2_X1 U386 ( .A(n336), .B(KEYINPUT31), .Z(n338) );
  NAND2_X1 U387 ( .A1(G230GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U388 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U389 ( .A(n340), .B(n339), .Z(n344) );
  XNOR2_X1 U390 ( .A(G106GAT), .B(G78GAT), .ZN(n341) );
  XNOR2_X1 U391 ( .A(n341), .B(G204GAT), .ZN(n426) );
  XNOR2_X1 U392 ( .A(G120GAT), .B(G148GAT), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n342), .B(G57GAT), .ZN(n409) );
  XNOR2_X1 U394 ( .A(n426), .B(n409), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U396 ( .A(n346), .B(n345), .ZN(n572) );
  XOR2_X1 U397 ( .A(G113GAT), .B(G29GAT), .Z(n348) );
  XNOR2_X1 U398 ( .A(G169GAT), .B(G36GAT), .ZN(n347) );
  XNOR2_X1 U399 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U400 ( .A(KEYINPUT70), .B(G1GAT), .Z(n350) );
  XNOR2_X1 U401 ( .A(G141GAT), .B(G197GAT), .ZN(n349) );
  XNOR2_X1 U402 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U403 ( .A(n352), .B(n351), .Z(n357) );
  XOR2_X1 U404 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n354) );
  NAND2_X1 U405 ( .A1(G229GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U406 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U407 ( .A(KEYINPUT68), .B(n355), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U409 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n359) );
  XNOR2_X1 U410 ( .A(KEYINPUT30), .B(KEYINPUT71), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U412 ( .A(n361), .B(n360), .Z(n365) );
  XNOR2_X1 U413 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U414 ( .A(n365), .B(n364), .Z(n507) );
  NOR2_X1 U415 ( .A1(n572), .A2(n507), .ZN(n366) );
  AND2_X1 U416 ( .A1(n367), .A2(n366), .ZN(n368) );
  XNOR2_X1 U417 ( .A(n368), .B(KEYINPUT114), .ZN(n375) );
  NAND2_X1 U418 ( .A1(n369), .A2(n577), .ZN(n372) );
  INV_X1 U419 ( .A(n507), .ZN(n567) );
  XNOR2_X1 U420 ( .A(KEYINPUT41), .B(n572), .ZN(n546) );
  NOR2_X1 U421 ( .A1(n567), .A2(n546), .ZN(n370) );
  XNOR2_X1 U422 ( .A(n370), .B(KEYINPUT46), .ZN(n371) );
  NOR2_X1 U423 ( .A1(n372), .A2(n371), .ZN(n373) );
  XOR2_X1 U424 ( .A(KEYINPUT47), .B(n373), .Z(n374) );
  NOR2_X1 U425 ( .A1(n375), .A2(n374), .ZN(n377) );
  XOR2_X1 U426 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n379) );
  XNOR2_X1 U427 ( .A(KEYINPUT88), .B(KEYINPUT18), .ZN(n378) );
  XNOR2_X1 U428 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U429 ( .A(n380), .B(KEYINPUT89), .Z(n382) );
  XNOR2_X1 U430 ( .A(G169GAT), .B(G183GAT), .ZN(n381) );
  XNOR2_X1 U431 ( .A(n382), .B(n381), .ZN(n439) );
  XOR2_X1 U432 ( .A(KEYINPUT93), .B(G218GAT), .Z(n384) );
  XNOR2_X1 U433 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n383) );
  XNOR2_X1 U434 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U435 ( .A(G197GAT), .B(n385), .Z(n430) );
  XNOR2_X1 U436 ( .A(n439), .B(n430), .ZN(n397) );
  XOR2_X1 U437 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n387) );
  XNOR2_X1 U438 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n386) );
  XNOR2_X1 U439 ( .A(n387), .B(n386), .ZN(n393) );
  XOR2_X1 U440 ( .A(n389), .B(n388), .Z(n391) );
  XNOR2_X1 U441 ( .A(G204GAT), .B(G92GAT), .ZN(n390) );
  XNOR2_X1 U442 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U443 ( .A(n393), .B(n392), .Z(n395) );
  NAND2_X1 U444 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U445 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U446 ( .A(n397), .B(n396), .ZN(n521) );
  NOR2_X1 U447 ( .A1(n543), .A2(n521), .ZN(n398) );
  XNOR2_X1 U448 ( .A(n398), .B(KEYINPUT54), .ZN(n418) );
  XOR2_X1 U449 ( .A(KEYINPUT2), .B(G162GAT), .Z(n400) );
  XNOR2_X1 U450 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n399) );
  XNOR2_X1 U451 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U452 ( .A(G141GAT), .B(n401), .ZN(n433) );
  XOR2_X1 U453 ( .A(KEYINPUT96), .B(KEYINPUT4), .Z(n403) );
  XNOR2_X1 U454 ( .A(KEYINPUT97), .B(KEYINPUT1), .ZN(n402) );
  XNOR2_X1 U455 ( .A(n403), .B(n402), .ZN(n416) );
  XOR2_X1 U456 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n405) );
  XNOR2_X1 U457 ( .A(G85GAT), .B(KEYINPUT95), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n405), .B(n404), .ZN(n407) );
  XOR2_X1 U459 ( .A(n407), .B(n406), .Z(n414) );
  XOR2_X1 U460 ( .A(G113GAT), .B(KEYINPUT0), .Z(n449) );
  XOR2_X1 U461 ( .A(n409), .B(n408), .Z(n411) );
  NAND2_X1 U462 ( .A1(G225GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U463 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U464 ( .A(n449), .B(n412), .ZN(n413) );
  XNOR2_X1 U465 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U466 ( .A(n416), .B(n415), .Z(n417) );
  XNOR2_X1 U467 ( .A(n433), .B(n417), .ZN(n467) );
  XOR2_X1 U468 ( .A(KEYINPUT98), .B(n467), .Z(n471) );
  INV_X1 U469 ( .A(n471), .ZN(n519) );
  NAND2_X1 U470 ( .A1(n418), .A2(n519), .ZN(n419) );
  XNOR2_X1 U471 ( .A(n419), .B(KEYINPUT65), .ZN(n566) );
  XOR2_X1 U472 ( .A(KEYINPUT24), .B(KEYINPUT91), .Z(n421) );
  XNOR2_X1 U473 ( .A(G50GAT), .B(KEYINPUT92), .ZN(n420) );
  XNOR2_X1 U474 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U475 ( .A(G148GAT), .B(KEYINPUT23), .Z(n423) );
  XNOR2_X1 U476 ( .A(KEYINPUT22), .B(KEYINPUT94), .ZN(n422) );
  XNOR2_X1 U477 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U478 ( .A(n425), .B(n424), .Z(n432) );
  XOR2_X1 U479 ( .A(G22GAT), .B(n426), .Z(n428) );
  NAND2_X1 U480 ( .A1(G228GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U483 ( .A(n432), .B(n431), .ZN(n434) );
  XNOR2_X1 U484 ( .A(n434), .B(n433), .ZN(n472) );
  NAND2_X1 U485 ( .A1(n566), .A2(n472), .ZN(n435) );
  XNOR2_X1 U486 ( .A(KEYINPUT55), .B(n435), .ZN(n454) );
  XOR2_X1 U487 ( .A(KEYINPUT90), .B(KEYINPUT87), .Z(n437) );
  XNOR2_X1 U488 ( .A(G120GAT), .B(KEYINPUT85), .ZN(n436) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n453) );
  XOR2_X1 U491 ( .A(G99GAT), .B(G134GAT), .Z(n441) );
  XNOR2_X1 U492 ( .A(G43GAT), .B(G190GAT), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U494 ( .A(G71GAT), .B(KEYINPUT86), .Z(n443) );
  XNOR2_X1 U495 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U497 ( .A(n445), .B(n444), .Z(n451) );
  XOR2_X1 U498 ( .A(G176GAT), .B(G127GAT), .Z(n447) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U503 ( .A(n453), .B(n452), .Z(n523) );
  INV_X1 U504 ( .A(n523), .ZN(n532) );
  NAND2_X1 U505 ( .A1(n454), .A2(n532), .ZN(n560) );
  NOR2_X1 U506 ( .A1(n577), .A2(n560), .ZN(n457) );
  XNOR2_X1 U507 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n455) );
  NOR2_X1 U508 ( .A1(n560), .A2(n369), .ZN(n458) );
  XNOR2_X1 U509 ( .A(KEYINPUT58), .B(n458), .ZN(n460) );
  INV_X1 U510 ( .A(G190GAT), .ZN(n459) );
  XNOR2_X1 U511 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  NOR2_X1 U512 ( .A1(n567), .A2(n572), .ZN(n495) );
  XOR2_X1 U513 ( .A(n521), .B(KEYINPUT27), .Z(n470) );
  XNOR2_X1 U514 ( .A(KEYINPUT26), .B(KEYINPUT102), .ZN(n462) );
  NOR2_X1 U515 ( .A1(n532), .A2(n472), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n462), .B(n461), .ZN(n565) );
  NAND2_X1 U517 ( .A1(n470), .A2(n565), .ZN(n466) );
  OR2_X1 U518 ( .A1(n523), .A2(n521), .ZN(n463) );
  NAND2_X1 U519 ( .A1(n472), .A2(n463), .ZN(n464) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(n464), .Z(n465) );
  NAND2_X1 U521 ( .A1(n466), .A2(n465), .ZN(n468) );
  NAND2_X1 U522 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U523 ( .A(n469), .B(KEYINPUT103), .ZN(n476) );
  NAND2_X1 U524 ( .A1(n471), .A2(n470), .ZN(n542) );
  INV_X1 U525 ( .A(n542), .ZN(n474) );
  XOR2_X1 U526 ( .A(n472), .B(KEYINPUT28), .Z(n473) );
  XNOR2_X1 U527 ( .A(KEYINPUT67), .B(n473), .ZN(n526) );
  NAND2_X1 U528 ( .A1(n474), .A2(n526), .ZN(n530) );
  NOR2_X1 U529 ( .A1(n530), .A2(n532), .ZN(n475) );
  NOR2_X1 U530 ( .A1(n476), .A2(n475), .ZN(n491) );
  NAND2_X1 U531 ( .A1(n477), .A2(n369), .ZN(n478) );
  XNOR2_X1 U532 ( .A(n478), .B(KEYINPUT84), .ZN(n479) );
  XNOR2_X1 U533 ( .A(n479), .B(KEYINPUT16), .ZN(n480) );
  NOR2_X1 U534 ( .A1(n491), .A2(n480), .ZN(n481) );
  XNOR2_X1 U535 ( .A(KEYINPUT104), .B(n481), .ZN(n508) );
  NAND2_X1 U536 ( .A1(n495), .A2(n508), .ZN(n489) );
  NOR2_X1 U537 ( .A1(n519), .A2(n489), .ZN(n482) );
  XOR2_X1 U538 ( .A(G1GAT), .B(n482), .Z(n483) );
  XNOR2_X1 U539 ( .A(KEYINPUT34), .B(n483), .ZN(G1324GAT) );
  NOR2_X1 U540 ( .A1(n521), .A2(n489), .ZN(n485) );
  XNOR2_X1 U541 ( .A(G8GAT), .B(KEYINPUT105), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n485), .B(n484), .ZN(G1325GAT) );
  NOR2_X1 U543 ( .A1(n523), .A2(n489), .ZN(n487) );
  XNOR2_X1 U544 ( .A(KEYINPUT106), .B(KEYINPUT35), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(n488), .ZN(G1326GAT) );
  NOR2_X1 U547 ( .A1(n526), .A2(n489), .ZN(n490) );
  XOR2_X1 U548 ( .A(G22GAT), .B(n490), .Z(G1327GAT) );
  NOR2_X1 U549 ( .A1(n491), .A2(n580), .ZN(n492) );
  NAND2_X1 U550 ( .A1(n492), .A2(n577), .ZN(n494) );
  XOR2_X1 U551 ( .A(KEYINPUT107), .B(KEYINPUT37), .Z(n493) );
  XNOR2_X1 U552 ( .A(n494), .B(n493), .ZN(n518) );
  NAND2_X1 U553 ( .A1(n495), .A2(n518), .ZN(n496) );
  XNOR2_X1 U554 ( .A(n496), .B(KEYINPUT108), .ZN(n497) );
  XNOR2_X1 U555 ( .A(KEYINPUT38), .B(n497), .ZN(n505) );
  NOR2_X1 U556 ( .A1(n519), .A2(n505), .ZN(n499) );
  XNOR2_X1 U557 ( .A(KEYINPUT109), .B(KEYINPUT39), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U559 ( .A(G29GAT), .B(n500), .Z(G1328GAT) );
  NOR2_X1 U560 ( .A1(n521), .A2(n505), .ZN(n501) );
  XOR2_X1 U561 ( .A(KEYINPUT110), .B(n501), .Z(n502) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n502), .ZN(G1329GAT) );
  NOR2_X1 U563 ( .A1(n523), .A2(n505), .ZN(n503) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(n503), .Z(n504) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n504), .ZN(G1330GAT) );
  NOR2_X1 U566 ( .A1(n526), .A2(n505), .ZN(n506) );
  XOR2_X1 U567 ( .A(G50GAT), .B(n506), .Z(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT111), .B(n546), .Z(n559) );
  NOR2_X1 U569 ( .A1(n507), .A2(n559), .ZN(n517) );
  NAND2_X1 U570 ( .A1(n517), .A2(n508), .ZN(n513) );
  NOR2_X1 U571 ( .A1(n519), .A2(n513), .ZN(n509) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n509), .Z(n510) );
  XNOR2_X1 U573 ( .A(KEYINPUT42), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U574 ( .A1(n521), .A2(n513), .ZN(n511) );
  XOR2_X1 U575 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U576 ( .A1(n523), .A2(n513), .ZN(n512) );
  XOR2_X1 U577 ( .A(G71GAT), .B(n512), .Z(G1334GAT) );
  NOR2_X1 U578 ( .A1(n526), .A2(n513), .ZN(n515) );
  XNOR2_X1 U579 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n525) );
  NOR2_X1 U583 ( .A1(n519), .A2(n525), .ZN(n520) );
  XOR2_X1 U584 ( .A(G85GAT), .B(n520), .Z(G1336GAT) );
  NOR2_X1 U585 ( .A1(n521), .A2(n525), .ZN(n522) );
  XOR2_X1 U586 ( .A(G92GAT), .B(n522), .Z(G1337GAT) );
  NOR2_X1 U587 ( .A1(n523), .A2(n525), .ZN(n524) );
  XOR2_X1 U588 ( .A(G99GAT), .B(n524), .Z(G1338GAT) );
  NOR2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NOR2_X1 U593 ( .A1(n543), .A2(n530), .ZN(n531) );
  NAND2_X1 U594 ( .A1(n532), .A2(n531), .ZN(n539) );
  NOR2_X1 U595 ( .A1(n567), .A2(n539), .ZN(n533) );
  XOR2_X1 U596 ( .A(G113GAT), .B(n533), .Z(G1340GAT) );
  NOR2_X1 U597 ( .A1(n559), .A2(n539), .ZN(n535) );
  XNOR2_X1 U598 ( .A(KEYINPUT49), .B(KEYINPUT115), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U600 ( .A(G120GAT), .B(n536), .Z(G1341GAT) );
  NOR2_X1 U601 ( .A1(n577), .A2(n539), .ZN(n537) );
  XOR2_X1 U602 ( .A(KEYINPUT50), .B(n537), .Z(n538) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  NOR2_X1 U604 ( .A1(n369), .A2(n539), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NOR2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U608 ( .A1(n565), .A2(n544), .ZN(n555) );
  NOR2_X1 U609 ( .A1(n567), .A2(n555), .ZN(n545) );
  XOR2_X1 U610 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  NOR2_X1 U611 ( .A1(n546), .A2(n555), .ZN(n551) );
  XOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n548) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(KEYINPUT52), .B(n549), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NOR2_X1 U617 ( .A1(n577), .A2(n555), .ZN(n553) );
  XNOR2_X1 U618 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G155GAT), .B(n554), .ZN(G1346GAT) );
  NOR2_X1 U621 ( .A1(n369), .A2(n555), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT120), .B(n556), .Z(n557) );
  XNOR2_X1 U623 ( .A(G162GAT), .B(n557), .ZN(G1347GAT) );
  NOR2_X1 U624 ( .A1(n567), .A2(n560), .ZN(n558) );
  XOR2_X1 U625 ( .A(G169GAT), .B(n558), .Z(G1348GAT) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n579) );
  NOR2_X1 U633 ( .A1(n567), .A2(n579), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n575) );
  INV_X1 U638 ( .A(n579), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n576), .Z(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n579), .ZN(n578) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n578), .Z(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(G218GAT), .B(n583), .Z(G1355GAT) );
endmodule

