

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U323 ( .A(n473), .B(KEYINPUT48), .ZN(n539) );
  XNOR2_X1 U324 ( .A(n417), .B(n416), .ZN(n456) );
  XNOR2_X1 U325 ( .A(n350), .B(n349), .ZN(n352) );
  XNOR2_X1 U326 ( .A(KEYINPUT45), .B(KEYINPUT65), .ZN(n461) );
  XNOR2_X1 U327 ( .A(n462), .B(n461), .ZN(n463) );
  INV_X1 U328 ( .A(G218GAT), .ZN(n397) );
  XNOR2_X1 U329 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U330 ( .A(n437), .B(n399), .ZN(n403) );
  XNOR2_X1 U331 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U332 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n349) );
  XNOR2_X1 U333 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U334 ( .A(n377), .B(n376), .ZN(n379) );
  XNOR2_X1 U335 ( .A(KEYINPUT105), .B(KEYINPUT37), .ZN(n416) );
  NOR2_X1 U336 ( .A1(n526), .A2(n477), .ZN(n386) );
  XNOR2_X1 U337 ( .A(n410), .B(n409), .ZN(n414) );
  XNOR2_X1 U338 ( .A(n423), .B(n381), .ZN(n382) );
  XNOR2_X1 U339 ( .A(n383), .B(n382), .ZN(n480) );
  XNOR2_X1 U340 ( .A(n457), .B(KEYINPUT114), .ZN(n524) );
  XNOR2_X1 U341 ( .A(n452), .B(n451), .ZN(n503) );
  XNOR2_X1 U342 ( .A(n481), .B(G176GAT), .ZN(n482) );
  XNOR2_X1 U343 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n459) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n453) );
  XNOR2_X1 U345 ( .A(n483), .B(n482), .ZN(G1349GAT) );
  XNOR2_X1 U346 ( .A(n454), .B(n453), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(G155GAT), .B(KEYINPUT79), .Z(n292) );
  XNOR2_X1 U348 ( .A(G22GAT), .B(G127GAT), .ZN(n291) );
  XNOR2_X1 U349 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U350 ( .A(G71GAT), .B(G183GAT), .Z(n294) );
  XNOR2_X1 U351 ( .A(G8GAT), .B(G15GAT), .ZN(n293) );
  XNOR2_X1 U352 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U353 ( .A(n296), .B(n295), .Z(n301) );
  XOR2_X1 U354 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n298) );
  NAND2_X1 U355 ( .A1(G231GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U356 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U357 ( .A(KEYINPUT14), .B(n299), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n301), .B(n300), .ZN(n310) );
  XOR2_X1 U359 ( .A(KEYINPUT12), .B(G78GAT), .Z(n303) );
  XNOR2_X1 U360 ( .A(G64GAT), .B(G211GAT), .ZN(n302) );
  XNOR2_X1 U361 ( .A(n303), .B(n302), .ZN(n308) );
  XOR2_X1 U362 ( .A(KEYINPUT13), .B(G57GAT), .Z(n446) );
  XOR2_X1 U363 ( .A(n446), .B(KEYINPUT80), .Z(n306) );
  XNOR2_X1 U364 ( .A(G1GAT), .B(KEYINPUT67), .ZN(n304) );
  XNOR2_X1 U365 ( .A(n304), .B(KEYINPUT68), .ZN(n418) );
  XNOR2_X1 U366 ( .A(n418), .B(KEYINPUT78), .ZN(n305) );
  XNOR2_X1 U367 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U368 ( .A(n308), .B(n307), .Z(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n557) );
  XOR2_X1 U370 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n312) );
  XNOR2_X1 U371 ( .A(KEYINPUT4), .B(KEYINPUT93), .ZN(n311) );
  XNOR2_X1 U372 ( .A(n312), .B(n311), .ZN(n318) );
  XOR2_X1 U373 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n314) );
  XNOR2_X1 U374 ( .A(G162GAT), .B(G155GAT), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n314), .B(n313), .ZN(n358) );
  XOR2_X1 U376 ( .A(n358), .B(KEYINPUT6), .Z(n316) );
  NAND2_X1 U377 ( .A1(G225GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U378 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n333) );
  XOR2_X1 U380 ( .A(G148GAT), .B(G120GAT), .Z(n320) );
  XNOR2_X1 U381 ( .A(G113GAT), .B(G141GAT), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U383 ( .A(KEYINPUT1), .B(KEYINPUT95), .Z(n322) );
  XNOR2_X1 U384 ( .A(KEYINPUT96), .B(KEYINPUT94), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U386 ( .A(n324), .B(n323), .Z(n331) );
  XOR2_X1 U387 ( .A(G57GAT), .B(G85GAT), .Z(n328) );
  XOR2_X1 U388 ( .A(KEYINPUT0), .B(KEYINPUT81), .Z(n326) );
  XNOR2_X1 U389 ( .A(G134GAT), .B(G127GAT), .ZN(n325) );
  XNOR2_X1 U390 ( .A(n326), .B(n325), .ZN(n381) );
  XNOR2_X1 U391 ( .A(G29GAT), .B(n381), .ZN(n327) );
  XNOR2_X1 U392 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U393 ( .A(G1GAT), .B(n329), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n519) );
  XOR2_X1 U396 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n341) );
  XNOR2_X1 U397 ( .A(G169GAT), .B(G36GAT), .ZN(n334) );
  XNOR2_X1 U398 ( .A(n334), .B(G8GAT), .ZN(n424) );
  XOR2_X1 U399 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n336) );
  XNOR2_X1 U400 ( .A(G218GAT), .B(G211GAT), .ZN(n335) );
  XNOR2_X1 U401 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n337), .B(KEYINPUT89), .ZN(n339) );
  XOR2_X1 U403 ( .A(G197GAT), .B(KEYINPUT90), .Z(n338) );
  XNOR2_X1 U404 ( .A(n339), .B(n338), .ZN(n365) );
  XNOR2_X1 U405 ( .A(n424), .B(n365), .ZN(n340) );
  XNOR2_X1 U406 ( .A(n341), .B(n340), .ZN(n348) );
  XOR2_X1 U407 ( .A(G204GAT), .B(KEYINPUT74), .Z(n343) );
  XNOR2_X1 U408 ( .A(G92GAT), .B(G64GAT), .ZN(n342) );
  XNOR2_X1 U409 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U410 ( .A(G176GAT), .B(n344), .Z(n450) );
  XOR2_X1 U411 ( .A(n450), .B(KEYINPUT98), .Z(n346) );
  NAND2_X1 U412 ( .A1(G226GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U413 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U414 ( .A(n348), .B(n347), .Z(n354) );
  XNOR2_X1 U415 ( .A(KEYINPUT85), .B(KEYINPUT17), .ZN(n350) );
  XOR2_X1 U416 ( .A(KEYINPUT19), .B(G190GAT), .Z(n351) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n369) );
  XNOR2_X1 U418 ( .A(n369), .B(KEYINPUT77), .ZN(n353) );
  XOR2_X1 U419 ( .A(n354), .B(n353), .Z(n521) );
  XNOR2_X1 U420 ( .A(n521), .B(KEYINPUT27), .ZN(n387) );
  AND2_X1 U421 ( .A1(n519), .A2(n387), .ZN(n540) );
  XOR2_X1 U422 ( .A(KEYINPUT22), .B(G204GAT), .Z(n356) );
  XNOR2_X1 U423 ( .A(G50GAT), .B(G106GAT), .ZN(n355) );
  XNOR2_X1 U424 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U425 ( .A(n358), .B(n357), .Z(n360) );
  XOR2_X1 U426 ( .A(G22GAT), .B(G141GAT), .Z(n427) );
  XOR2_X1 U427 ( .A(G78GAT), .B(G148GAT), .Z(n445) );
  XNOR2_X1 U428 ( .A(n427), .B(n445), .ZN(n359) );
  XNOR2_X1 U429 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U430 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n362) );
  NAND2_X1 U431 ( .A1(G228GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U432 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U433 ( .A(n364), .B(n363), .Z(n367) );
  XNOR2_X1 U434 ( .A(n365), .B(KEYINPUT23), .ZN(n366) );
  XNOR2_X1 U435 ( .A(n367), .B(n366), .ZN(n477) );
  XNOR2_X1 U436 ( .A(n477), .B(KEYINPUT28), .ZN(n458) );
  NAND2_X1 U437 ( .A1(n540), .A2(n458), .ZN(n528) );
  XNOR2_X1 U438 ( .A(G99GAT), .B(G71GAT), .ZN(n368) );
  XNOR2_X1 U439 ( .A(n368), .B(G120GAT), .ZN(n438) );
  XNOR2_X1 U440 ( .A(n369), .B(n438), .ZN(n377) );
  XOR2_X1 U441 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n371) );
  XNOR2_X1 U442 ( .A(KEYINPUT84), .B(KEYINPUT87), .ZN(n370) );
  XNOR2_X1 U443 ( .A(n371), .B(n370), .ZN(n373) );
  XOR2_X1 U444 ( .A(G169GAT), .B(G176GAT), .Z(n372) );
  XNOR2_X1 U445 ( .A(n373), .B(n372), .ZN(n375) );
  XOR2_X1 U446 ( .A(KEYINPUT86), .B(KEYINPUT83), .Z(n374) );
  NAND2_X1 U447 ( .A1(G227GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n379), .B(n378), .ZN(n383) );
  XNOR2_X1 U449 ( .A(G43GAT), .B(G15GAT), .ZN(n380) );
  XOR2_X1 U450 ( .A(n380), .B(G113GAT), .Z(n423) );
  INV_X1 U451 ( .A(n480), .ZN(n526) );
  XNOR2_X1 U452 ( .A(KEYINPUT88), .B(n526), .ZN(n384) );
  NOR2_X1 U453 ( .A1(n528), .A2(n384), .ZN(n395) );
  XOR2_X1 U454 ( .A(KEYINPUT26), .B(KEYINPUT101), .Z(n385) );
  XNOR2_X1 U455 ( .A(n386), .B(n385), .ZN(n564) );
  NAND2_X1 U456 ( .A1(n387), .A2(n564), .ZN(n391) );
  NAND2_X1 U457 ( .A1(n526), .A2(n521), .ZN(n388) );
  NAND2_X1 U458 ( .A1(n477), .A2(n388), .ZN(n389) );
  XOR2_X1 U459 ( .A(KEYINPUT25), .B(n389), .Z(n390) );
  NAND2_X1 U460 ( .A1(n391), .A2(n390), .ZN(n392) );
  XOR2_X1 U461 ( .A(KEYINPUT102), .B(n392), .Z(n393) );
  NOR2_X1 U462 ( .A1(n519), .A2(n393), .ZN(n394) );
  NOR2_X1 U463 ( .A1(n395), .A2(n394), .ZN(n486) );
  NOR2_X1 U464 ( .A1(n557), .A2(n486), .ZN(n415) );
  XNOR2_X1 U465 ( .A(G85GAT), .B(KEYINPUT71), .ZN(n396) );
  XNOR2_X1 U466 ( .A(n396), .B(G106GAT), .ZN(n437) );
  NAND2_X1 U467 ( .A1(G232GAT), .A2(G233GAT), .ZN(n398) );
  XOR2_X1 U468 ( .A(KEYINPUT9), .B(KEYINPUT64), .Z(n401) );
  XNOR2_X1 U469 ( .A(KEYINPUT10), .B(KEYINPUT11), .ZN(n400) );
  XOR2_X1 U470 ( .A(n401), .B(n400), .Z(n402) );
  XNOR2_X1 U471 ( .A(n403), .B(n402), .ZN(n410) );
  XOR2_X1 U472 ( .A(G162GAT), .B(G134GAT), .Z(n405) );
  XNOR2_X1 U473 ( .A(G43GAT), .B(G190GAT), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U475 ( .A(G99GAT), .B(n406), .ZN(n408) );
  INV_X1 U476 ( .A(G92GAT), .ZN(n407) );
  XOR2_X1 U477 ( .A(G29GAT), .B(G50GAT), .Z(n412) );
  XNOR2_X1 U478 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n411) );
  XNOR2_X1 U479 ( .A(n412), .B(n411), .ZN(n419) );
  XNOR2_X1 U480 ( .A(n419), .B(G36GAT), .ZN(n413) );
  XNOR2_X1 U481 ( .A(n414), .B(n413), .ZN(n484) );
  XOR2_X1 U482 ( .A(n484), .B(KEYINPUT36), .Z(n579) );
  NAND2_X1 U483 ( .A1(n415), .A2(n579), .ZN(n417) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n432) );
  XOR2_X1 U485 ( .A(G197GAT), .B(KEYINPUT66), .Z(n421) );
  NAND2_X1 U486 ( .A1(G229GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U488 ( .A(n422), .B(KEYINPUT30), .Z(n426) );
  XOR2_X1 U489 ( .A(n424), .B(n423), .Z(n425) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U491 ( .A(n428), .B(n427), .Z(n430) );
  XNOR2_X1 U492 ( .A(KEYINPUT29), .B(KEYINPUT69), .ZN(n429) );
  XNOR2_X1 U493 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U494 ( .A(n432), .B(n431), .Z(n566) );
  XOR2_X1 U495 ( .A(n566), .B(KEYINPUT70), .Z(n555) );
  XOR2_X1 U496 ( .A(KEYINPUT32), .B(KEYINPUT75), .Z(n434) );
  NAND2_X1 U497 ( .A1(G230GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n436) );
  INV_X1 U499 ( .A(KEYINPUT33), .ZN(n435) );
  XNOR2_X1 U500 ( .A(n436), .B(n435), .ZN(n440) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U502 ( .A(n440), .B(n439), .Z(n444) );
  XOR2_X1 U503 ( .A(KEYINPUT31), .B(KEYINPUT76), .Z(n442) );
  XNOR2_X1 U504 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n441) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U506 ( .A(n444), .B(n443), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U508 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U509 ( .A(n450), .B(n449), .ZN(n572) );
  NAND2_X1 U510 ( .A1(n555), .A2(n572), .ZN(n489) );
  NOR2_X1 U511 ( .A1(n456), .A2(n489), .ZN(n452) );
  XNOR2_X1 U512 ( .A(KEYINPUT38), .B(KEYINPUT106), .ZN(n451) );
  NAND2_X1 U513 ( .A1(n503), .A2(n526), .ZN(n454) );
  XOR2_X1 U514 ( .A(KEYINPUT41), .B(n572), .Z(n546) );
  XNOR2_X1 U515 ( .A(KEYINPUT109), .B(n546), .ZN(n530) );
  NAND2_X1 U516 ( .A1(n566), .A2(n530), .ZN(n455) );
  XNOR2_X1 U517 ( .A(n455), .B(KEYINPUT110), .ZN(n508) );
  NOR2_X1 U518 ( .A1(n456), .A2(n508), .ZN(n457) );
  INV_X1 U519 ( .A(n458), .ZN(n514) );
  NAND2_X1 U520 ( .A1(n524), .A2(n514), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n460), .B(n459), .ZN(G1339GAT) );
  XNOR2_X1 U522 ( .A(KEYINPUT122), .B(n521), .ZN(n474) );
  NAND2_X1 U523 ( .A1(n557), .A2(n579), .ZN(n462) );
  NAND2_X1 U524 ( .A1(n463), .A2(n572), .ZN(n464) );
  NOR2_X1 U525 ( .A1(n464), .A2(n555), .ZN(n465) );
  XNOR2_X1 U526 ( .A(n465), .B(KEYINPUT117), .ZN(n472) );
  NOR2_X1 U527 ( .A1(n566), .A2(n546), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(KEYINPUT46), .ZN(n467) );
  NOR2_X1 U529 ( .A1(n557), .A2(n467), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n468), .B(KEYINPUT116), .ZN(n469) );
  AND2_X1 U531 ( .A1(n469), .A2(n484), .ZN(n470) );
  XNOR2_X1 U532 ( .A(KEYINPUT47), .B(n470), .ZN(n471) );
  NAND2_X1 U533 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U534 ( .A1(n474), .A2(n539), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n475), .B(KEYINPUT54), .ZN(n476) );
  NOR2_X2 U536 ( .A1(n476), .A2(n519), .ZN(n565) );
  NAND2_X1 U537 ( .A1(n477), .A2(n565), .ZN(n478) );
  XOR2_X1 U538 ( .A(n478), .B(KEYINPUT55), .Z(n479) );
  NOR2_X1 U539 ( .A1(n480), .A2(n479), .ZN(n561) );
  NAND2_X1 U540 ( .A1(n530), .A2(n561), .ZN(n483) );
  XOR2_X1 U541 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n481) );
  INV_X1 U542 ( .A(n557), .ZN(n575) );
  INV_X1 U543 ( .A(n484), .ZN(n560) );
  NOR2_X1 U544 ( .A1(n575), .A2(n560), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n485), .B(KEYINPUT16), .ZN(n488) );
  INV_X1 U546 ( .A(n486), .ZN(n487) );
  NAND2_X1 U547 ( .A1(n488), .A2(n487), .ZN(n507) );
  NOR2_X1 U548 ( .A1(n489), .A2(n507), .ZN(n496) );
  NAND2_X1 U549 ( .A1(n496), .A2(n519), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n490), .B(KEYINPUT34), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G1GAT), .B(n491), .ZN(G1324GAT) );
  NAND2_X1 U552 ( .A1(n521), .A2(n496), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n494) );
  NAND2_X1 U555 ( .A1(n496), .A2(n526), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U557 ( .A(G15GAT), .B(n495), .Z(G1326GAT) );
  NAND2_X1 U558 ( .A1(n496), .A2(n514), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(KEYINPUT104), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G22GAT), .B(n498), .ZN(G1327GAT) );
  XOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT39), .Z(n500) );
  NAND2_X1 U562 ( .A1(n503), .A2(n519), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  XOR2_X1 U564 ( .A(G36GAT), .B(KEYINPUT107), .Z(n502) );
  NAND2_X1 U565 ( .A1(n503), .A2(n521), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(G1329GAT) );
  NAND2_X1 U567 ( .A1(n503), .A2(n514), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n504), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n505), .B(KEYINPUT111), .ZN(n506) );
  XOR2_X1 U571 ( .A(KEYINPUT108), .B(n506), .Z(n510) );
  NOR2_X1 U572 ( .A1(n508), .A2(n507), .ZN(n515) );
  NAND2_X1 U573 ( .A1(n515), .A2(n519), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n521), .A2(n515), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n515), .A2(n526), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n512), .B(KEYINPUT112), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(n513), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT113), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U581 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U583 ( .A(G78GAT), .B(n518), .Z(G1335GAT) );
  NAND2_X1 U584 ( .A1(n524), .A2(n519), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n520), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U586 ( .A(G92GAT), .B(KEYINPUT115), .Z(n523) );
  NAND2_X1 U587 ( .A1(n524), .A2(n521), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n524), .A2(n526), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U591 ( .A1(n526), .A2(n539), .ZN(n527) );
  NOR2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n555), .A2(n535), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n529), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U596 ( .A1(n535), .A2(n530), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NAND2_X1 U598 ( .A1(n557), .A2(n535), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(KEYINPUT50), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n537) );
  NAND2_X1 U602 ( .A1(n535), .A2(n560), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(n538), .ZN(G1343GAT) );
  INV_X1 U605 ( .A(n539), .ZN(n542) );
  NAND2_X1 U606 ( .A1(n540), .A2(n564), .ZN(n541) );
  NOR2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U608 ( .A(KEYINPUT119), .B(n543), .Z(n553) );
  INV_X1 U609 ( .A(n553), .ZN(n547) );
  OR2_X1 U610 ( .A1(n547), .A2(n566), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n544), .B(KEYINPUT120), .ZN(n545) );
  XNOR2_X1 U612 ( .A(G141GAT), .B(n545), .ZN(G1344GAT) );
  NOR2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n551) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT121), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n557), .A2(n553), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n560), .A2(n553), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n561), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(G183GAT), .B(KEYINPUT123), .Z(n559) );
  NAND2_X1 U625 ( .A1(n561), .A2(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1350GAT) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1351GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n578) );
  NOR2_X1 U631 ( .A1(n566), .A2(n578), .ZN(n571) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT124), .B(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n578), .ZN(n574) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n578), .ZN(n576) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(n576), .Z(n577) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n582) );
  INV_X1 U644 ( .A(n578), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

