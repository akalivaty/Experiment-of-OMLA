//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n187));
  INV_X1    g001(.A(G131), .ZN(new_n188));
  INV_X1    g002(.A(G137), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n189), .A2(KEYINPUT11), .A3(G134), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT67), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT67), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n192), .A2(new_n189), .A3(KEYINPUT11), .A4(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n189), .A2(G134), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n197));
  OAI22_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .B1(new_n189), .B2(G134), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(KEYINPUT66), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n196), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n188), .B1(new_n195), .B2(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n201), .A2(new_n188), .A3(new_n191), .A4(new_n193), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT68), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT68), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n195), .A2(new_n205), .A3(new_n188), .A4(new_n201), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n202), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT65), .B1(new_n210), .B2(G143), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n208), .A3(G146), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n209), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT0), .B(G128), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n210), .A2(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n208), .A2(G146), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G128), .ZN(new_n219));
  OAI22_X1  g033(.A1(new_n214), .A2(new_n215), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n207), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n189), .A2(G134), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT69), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n196), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n223), .B(G131), .C1(new_n225), .C2(new_n222), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g042(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n219), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n211), .A2(new_n213), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n217), .ZN(new_n233));
  OR2_X1    g047(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n234));
  NAND2_X1  g048(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n217), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G128), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n231), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  AOI211_X1 g052(.A(new_n227), .B(new_n238), .C1(new_n204), .C2(new_n206), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n187), .B1(new_n221), .B2(new_n239), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n217), .A2(new_n232), .B1(new_n236), .B2(G128), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT74), .B1(new_n241), .B2(new_n231), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT74), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n234), .A2(new_n235), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n244), .A2(G128), .A3(new_n217), .A4(new_n218), .ZN(new_n245));
  INV_X1    g059(.A(G128), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n246), .B1(new_n230), .B2(new_n217), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n243), .B(new_n245), .C1(new_n247), .C2(new_n214), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n204), .A2(new_n206), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n250), .A3(new_n226), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n251), .B(KEYINPUT30), .C1(new_n207), .C2(new_n220), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT73), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n255));
  INV_X1    g069(.A(G119), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(G116), .ZN(new_n257));
  INV_X1    g071(.A(G116), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT71), .B1(new_n258), .B2(G119), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(G119), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n257), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT2), .B(G113), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n254), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n262), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n255), .B1(new_n256), .B2(G116), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n256), .A2(G116), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n264), .A2(KEYINPUT72), .A3(new_n267), .A4(new_n257), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n261), .A2(new_n262), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n253), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(new_n253), .A3(new_n270), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n240), .A2(new_n252), .A3(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(G237), .A2(G953), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G210), .ZN(new_n277));
  XOR2_X1   g091(.A(new_n277), .B(KEYINPUT27), .Z(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(KEYINPUT26), .ZN(new_n279));
  INV_X1    g093(.A(G101), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n202), .ZN(new_n282));
  INV_X1    g096(.A(new_n196), .ZN(new_n283));
  INV_X1    g097(.A(G134), .ZN(new_n284));
  AOI22_X1  g098(.A1(KEYINPUT66), .A2(new_n199), .B1(new_n284), .B2(G137), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n197), .A2(KEYINPUT11), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n283), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(new_n194), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n205), .B1(new_n288), .B2(new_n188), .ZN(new_n289));
  NOR4_X1   g103(.A1(new_n287), .A2(new_n194), .A3(KEYINPUT68), .A4(G131), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n282), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n220), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n227), .B1(new_n204), .B2(new_n206), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n291), .A2(new_n292), .B1(new_n293), .B2(new_n249), .ZN(new_n294));
  INV_X1    g108(.A(new_n273), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(new_n271), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT75), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n226), .B1(new_n289), .B2(new_n290), .ZN(new_n298));
  INV_X1    g112(.A(new_n248), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n233), .A2(new_n237), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n243), .B1(new_n300), .B2(new_n245), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  OAI22_X1  g116(.A1(new_n298), .A2(new_n302), .B1(new_n207), .B2(new_n220), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n303), .A2(new_n304), .A3(new_n274), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n275), .B(new_n281), .C1(new_n297), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT31), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT76), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT28), .B1(new_n294), .B2(new_n296), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n291), .A2(new_n292), .ZN(new_n312));
  INV_X1    g126(.A(new_n238), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n293), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n296), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n304), .B1(new_n303), .B2(new_n274), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n294), .A2(KEYINPUT75), .A3(new_n296), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT28), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n311), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n281), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n316), .A2(new_n317), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n323), .A2(new_n275), .A3(new_n281), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT31), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n306), .A2(KEYINPUT76), .A3(KEYINPUT31), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n309), .A2(new_n322), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(G472), .A2(G902), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT32), .ZN(new_n331));
  INV_X1    g145(.A(G472), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n303), .A2(new_n274), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n333), .B1(new_n305), .B2(new_n297), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n310), .B1(new_n334), .B2(KEYINPUT28), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT29), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n321), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(G902), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n281), .B(new_n311), .C1(new_n318), .C2(new_n319), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n323), .A2(new_n275), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n321), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n336), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n332), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n330), .A2(new_n331), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n343), .A2(new_n344), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n329), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n306), .A2(KEYINPUT76), .A3(KEYINPUT31), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT76), .B1(new_n306), .B2(KEYINPUT31), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n321), .A2(new_n320), .B1(new_n324), .B2(new_n325), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n348), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT78), .B1(new_n353), .B2(KEYINPUT32), .ZN(new_n354));
  AND4_X1   g168(.A1(KEYINPUT78), .A2(new_n328), .A3(KEYINPUT32), .A4(new_n329), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n345), .B(new_n347), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  INV_X1    g171(.A(G902), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(G234), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G953), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(G221), .A3(G234), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT22), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(G137), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT16), .ZN(new_n365));
  XNOR2_X1  g179(.A(G125), .B(G140), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT80), .ZN(new_n367));
  INV_X1    g181(.A(G140), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G125), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n369), .A2(KEYINPUT80), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n365), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n369), .A2(KEYINPUT16), .ZN(new_n372));
  OR3_X1    g186(.A1(new_n371), .A2(new_n210), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n210), .B1(new_n371), .B2(new_n372), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  OR2_X1    g190(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n377), .A2(G119), .A3(new_n246), .A4(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G119), .B(G128), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n379), .B1(new_n381), .B2(new_n378), .ZN(new_n382));
  INV_X1    g196(.A(G110), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT24), .B(G110), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n376), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n373), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n382), .A2(new_n383), .B1(new_n381), .B2(new_n385), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n366), .A2(new_n210), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n364), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  OAI221_X1 g207(.A(new_n375), .B1(new_n383), .B2(new_n382), .C1(new_n381), .C2(new_n385), .ZN(new_n394));
  INV_X1    g208(.A(new_n392), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(new_n363), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n358), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT25), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n397), .A2(new_n398), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n359), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n359), .A2(G902), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n393), .A2(new_n396), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n356), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g220(.A(KEYINPUT9), .B(G234), .Z(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G221), .B1(new_n408), .B2(G902), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G140), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n360), .A2(G227), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n207), .B(KEYINPUT82), .ZN(new_n415));
  INV_X1    g229(.A(G104), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G107), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n416), .A2(G107), .ZN(new_n419));
  OAI21_X1  g233(.A(G101), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT3), .B1(new_n416), .B2(G107), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT3), .ZN(new_n422));
  INV_X1    g236(.A(G107), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(G104), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n421), .A2(new_n424), .A3(new_n280), .A4(new_n417), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n249), .A2(KEYINPUT10), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT10), .ZN(new_n428));
  INV_X1    g242(.A(new_n219), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT1), .ZN(new_n430));
  OAI21_X1  g244(.A(G128), .B1(new_n209), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n217), .A2(new_n218), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n429), .A2(new_n244), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n420), .A2(new_n425), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n433), .A2(KEYINPUT81), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT81), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n431), .A2(new_n432), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n245), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n426), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n428), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n425), .A2(KEYINPUT4), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n421), .A2(new_n424), .A3(new_n417), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G101), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n441), .B(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n292), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n427), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n415), .A2(new_n446), .ZN(new_n447));
  OAI22_X1  g261(.A1(new_n435), .A2(new_n439), .B1(new_n313), .B2(new_n426), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT12), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n448), .A2(KEYINPUT83), .A3(new_n449), .A4(new_n291), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(KEYINPUT83), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n449), .A2(KEYINPUT83), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT81), .B1(new_n433), .B2(new_n434), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n426), .A2(new_n438), .A3(new_n436), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n453), .A2(new_n454), .B1(new_n238), .B2(new_n434), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n451), .B(new_n452), .C1(new_n455), .C2(new_n207), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n414), .B1(new_n447), .B2(new_n457), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n427), .A2(new_n440), .A3(new_n445), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT82), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n207), .B(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n414), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n446), .A2(new_n291), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n458), .A2(new_n464), .A3(G469), .ZN(new_n465));
  NAND2_X1  g279(.A1(G469), .A2(G902), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n457), .A2(KEYINPUT84), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT84), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n450), .A2(new_n456), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n462), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n459), .A2(new_n461), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n463), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n414), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G469), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(new_n358), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n410), .B1(new_n468), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(G234), .A2(G237), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(G902), .A3(G953), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n481), .B(KEYINPUT103), .Z(new_n482));
  XOR2_X1   g296(.A(KEYINPUT21), .B(G898), .Z(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT102), .B(G952), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(G953), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n480), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(G143), .B1(new_n276), .B2(G214), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n276), .A2(G143), .A3(G214), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n188), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT18), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n367), .A2(G146), .A3(new_n370), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n390), .ZN(new_n496));
  NAND2_X1  g310(.A1(KEYINPUT18), .A2(G131), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n491), .A2(new_n492), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n494), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT90), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT90), .A4(new_n498), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n491), .A2(new_n188), .A3(new_n492), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(new_n493), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n493), .A2(KEYINPUT17), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n507), .A2(new_n373), .A3(new_n374), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(G113), .B(G122), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(new_n416), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT94), .ZN(new_n514));
  INV_X1    g328(.A(new_n512), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n505), .A2(KEYINPUT91), .ZN(new_n516));
  NOR2_X1   g330(.A1(KEYINPUT92), .A2(KEYINPUT19), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n366), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n367), .A2(new_n370), .B1(KEYINPUT92), .B2(new_n366), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT19), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n210), .B(new_n518), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT91), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n504), .B2(new_n493), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n516), .A2(new_n373), .A3(new_n521), .A4(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n503), .A2(new_n515), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n513), .A2(new_n514), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT20), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(G475), .A2(G902), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT93), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n513), .A2(new_n525), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n513), .A2(new_n525), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n533), .A2(KEYINPUT94), .A3(new_n527), .A4(new_n530), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G122), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(G116), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(G116), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(new_n423), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n246), .A2(G143), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(KEYINPUT13), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n208), .A2(G128), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n543), .A2(KEYINPUT13), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT13), .ZN(new_n548));
  OAI211_X1 g362(.A(KEYINPUT97), .B(new_n548), .C1(new_n246), .C2(G143), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n544), .A2(new_n546), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G134), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n545), .A2(new_n543), .A3(G134), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT98), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n541), .A2(new_n551), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n540), .A2(new_n423), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n545), .A2(new_n543), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(new_n284), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT99), .B1(new_n538), .B2(KEYINPUT14), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n538), .A2(KEYINPUT14), .ZN(new_n561));
  OR4_X1    g375(.A1(KEYINPUT99), .A2(new_n536), .A3(KEYINPUT14), .A4(G116), .ZN(new_n562));
  AND4_X1   g376(.A1(new_n539), .A2(new_n560), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n557), .B(new_n559), .C1(new_n563), .C2(new_n423), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n556), .A2(new_n564), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n408), .A2(new_n357), .A3(G953), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT100), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n556), .A2(new_n564), .A3(new_n566), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n565), .A2(KEYINPUT100), .A3(new_n567), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n571), .A2(KEYINPUT101), .A3(new_n358), .A4(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G478), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n574), .A2(KEYINPUT15), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n573), .B(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n510), .B1(new_n577), .B2(new_n512), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n503), .A2(new_n509), .A3(KEYINPUT95), .A4(new_n515), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n358), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT96), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT96), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n578), .A2(new_n579), .A3(new_n582), .A4(new_n358), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(G475), .A3(new_n583), .ZN(new_n584));
  AND4_X1   g398(.A1(new_n489), .A2(new_n535), .A3(new_n576), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n479), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g400(.A(G110), .B(G122), .Z(new_n587));
  INV_X1    g401(.A(new_n444), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n272), .B2(new_n273), .ZN(new_n589));
  MUX2_X1   g403(.A(new_n266), .B(new_n261), .S(KEYINPUT5), .Z(new_n590));
  AOI22_X1  g404(.A1(new_n590), .A2(G113), .B1(new_n263), .B2(new_n268), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n426), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n587), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n587), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n592), .B(new_n595), .C1(new_n296), .C2(new_n588), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(KEYINPUT6), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT86), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n220), .A2(G125), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT85), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G125), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n238), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n598), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(G224), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(G953), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n599), .A2(new_n600), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT85), .B1(new_n220), .B2(G125), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n598), .B(new_n603), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n605), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n610), .ZN(new_n612));
  OAI22_X1  g426(.A1(new_n604), .A2(new_n612), .B1(new_n606), .B2(G953), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT6), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n614), .B(new_n587), .C1(new_n589), .C2(new_n593), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n597), .A2(new_n611), .A3(new_n613), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n601), .A2(new_n603), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT7), .ZN(new_n618));
  OR3_X1    g432(.A1(new_n617), .A2(new_n618), .A3(new_n607), .ZN(new_n619));
  OR2_X1    g433(.A1(new_n592), .A2(KEYINPUT88), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT87), .B(KEYINPUT8), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n587), .B(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT88), .B1(new_n591), .B2(new_n426), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n620), .B(new_n622), .C1(new_n593), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n603), .A2(new_n599), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n625), .B1(new_n618), .B2(new_n607), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n619), .A2(new_n624), .A3(new_n596), .A4(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n616), .A2(new_n627), .A3(new_n358), .ZN(new_n628));
  OAI21_X1  g442(.A(G210), .B1(G237), .B2(G902), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT89), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n616), .A2(new_n627), .A3(new_n358), .A4(new_n629), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n633), .A2(new_n632), .ZN(new_n635));
  OAI21_X1  g449(.A(G214), .B1(G237), .B2(G902), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n586), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(KEYINPUT104), .B1(new_n586), .B2(new_n637), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n406), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n280), .ZN(G3));
  AOI21_X1  g458(.A(new_n332), .B1(new_n328), .B2(new_n358), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n353), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n479), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n647), .A2(new_n404), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n631), .A2(new_n633), .ZN(new_n650));
  INV_X1    g464(.A(new_n636), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n485), .B2(new_n488), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n535), .A2(new_n584), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n571), .A2(new_n572), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n358), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n574), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT33), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n568), .A2(KEYINPUT33), .A3(new_n570), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n358), .A2(G478), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n654), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n653), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n649), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n416), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT105), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT34), .Z(G6));
  INV_X1    g483(.A(new_n576), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n531), .B(KEYINPUT20), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n584), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n653), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n649), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT35), .B(G107), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  NAND2_X1  g490(.A1(new_n394), .A2(new_n395), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n402), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n401), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n640), .A2(new_n641), .A3(new_n646), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT106), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  INV_X1    g499(.A(new_n488), .ZN(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n686), .B1(new_n687), .B2(new_n482), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n672), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n651), .B1(new_n631), .B2(new_n633), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n681), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  AND4_X1   g506(.A1(new_n356), .A2(new_n479), .A3(new_n689), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n246), .ZN(G30));
  NAND2_X1  g508(.A1(new_n634), .A2(new_n635), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT107), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT38), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n697), .A2(new_n651), .A3(new_n681), .ZN(new_n698));
  AOI21_X1  g512(.A(KEYINPUT32), .B1(new_n328), .B2(new_n329), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n324), .B1(new_n321), .B2(new_n334), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n701), .B2(G902), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n700), .B(new_n702), .C1(new_n354), .C2(new_n355), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT108), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n353), .A2(KEYINPUT78), .A3(KEYINPUT32), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n328), .A2(KEYINPUT32), .A3(new_n329), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT78), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(new_n710), .A3(new_n700), .A4(new_n702), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n688), .B(KEYINPUT39), .Z(new_n713));
  NAND2_X1  g527(.A1(new_n479), .A2(new_n713), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n714), .A2(KEYINPUT40), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(KEYINPUT40), .ZN(new_n716));
  INV_X1    g530(.A(new_n654), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n576), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n698), .A2(new_n712), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT109), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n208), .ZN(G45));
  INV_X1    g536(.A(new_n688), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n654), .A2(new_n663), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n356), .A2(new_n479), .A3(new_n692), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT110), .ZN(new_n727));
  AOI211_X1 g541(.A(KEYINPUT77), .B(new_n332), .C1(new_n338), .C2(new_n342), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n346), .A2(new_n699), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n648), .B1(new_n729), .B2(new_n709), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n731), .A3(new_n692), .A4(new_n725), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G146), .ZN(G48));
  INV_X1    g548(.A(new_n476), .ZN(new_n735));
  OAI21_X1  g549(.A(G469), .B1(new_n735), .B2(G902), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n409), .A3(new_n478), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n356), .A2(new_n405), .A3(new_n665), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT41), .B(G113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  NAND4_X1  g555(.A1(new_n356), .A2(new_n405), .A3(new_n673), .A4(new_n738), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT111), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n404), .B1(new_n729), .B2(new_n709), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(new_n745), .A3(new_n673), .A4(new_n738), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  NOR2_X1   g562(.A1(new_n691), .A2(new_n737), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n356), .A2(new_n585), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  AOI22_X1  g565(.A1(new_n316), .A2(new_n317), .B1(new_n274), .B2(new_n303), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n311), .B1(new_n752), .B2(new_n319), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g569(.A(KEYINPUT112), .B(new_n311), .C1(new_n752), .C2(new_n319), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n321), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n306), .B(new_n325), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n348), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n645), .A2(new_n759), .A3(new_n404), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n718), .A2(new_n690), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n489), .A4(new_n738), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  NOR3_X1   g577(.A1(new_n645), .A2(new_n759), .A3(new_n724), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n764), .A2(new_n765), .A3(new_n749), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n765), .B1(new_n764), .B2(new_n749), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n602), .ZN(G27));
  AOI211_X1 g583(.A(G469), .B(G902), .C1(new_n472), .C2(new_n475), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT114), .B1(new_n770), .B2(new_n467), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n468), .A2(new_n478), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n410), .A2(new_n651), .ZN(new_n775));
  AND4_X1   g589(.A1(new_n695), .A2(new_n774), .A3(new_n725), .A4(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n356), .A2(new_n405), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT115), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n744), .A2(new_n779), .A3(new_n776), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT42), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n729), .A2(new_n706), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n405), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(KEYINPUT42), .A3(new_n776), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G131), .ZN(G33));
  NAND2_X1  g602(.A1(new_n695), .A2(new_n775), .ZN(new_n789));
  INV_X1    g603(.A(new_n774), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n356), .A2(new_n405), .A3(new_n689), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G134), .ZN(G36));
  NAND2_X1  g607(.A1(new_n458), .A2(new_n464), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT45), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(G469), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT46), .B1(new_n796), .B2(new_n466), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n770), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n466), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n800), .A2(new_n409), .A3(new_n713), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n717), .A2(new_n663), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT43), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n647), .A3(new_n681), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT44), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n695), .A2(new_n636), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n804), .A2(new_n647), .A3(KEYINPUT44), .A4(new_n681), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n801), .A2(new_n807), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G137), .ZN(G39));
  NAND2_X1  g626(.A1(new_n800), .A2(new_n409), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT47), .Z(new_n814));
  NOR2_X1   g628(.A1(new_n808), .A2(new_n688), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n356), .A2(new_n405), .A3(new_n664), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  NOR2_X1   g632(.A1(new_n712), .A2(new_n404), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n736), .A2(new_n478), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n802), .B1(new_n820), .B2(KEYINPUT49), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n820), .A2(KEYINPUT49), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n821), .A2(new_n822), .A3(new_n775), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n819), .A2(new_n697), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n681), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n645), .A2(new_n825), .A3(new_n759), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n776), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n825), .A2(new_n670), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n356), .A2(new_n479), .A3(new_n815), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n584), .A2(new_n671), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n792), .B(new_n827), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n664), .B1(new_n576), .B2(new_n654), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n635), .A2(new_n832), .A3(new_n634), .A4(new_n652), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n405), .A3(new_n479), .A4(new_n646), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n682), .B(new_n834), .C1(new_n406), .C2(new_n642), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n739), .A2(new_n762), .ZN(new_n837));
  INV_X1    g651(.A(new_n750), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n743), .B2(new_n746), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n787), .A2(new_n836), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n768), .B(new_n693), .C1(new_n727), .C2(new_n732), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n761), .A2(new_n723), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n790), .A2(new_n681), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n712), .A2(new_n409), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT52), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n693), .B1(new_n727), .B2(new_n732), .ZN(new_n846));
  INV_X1    g660(.A(new_n768), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(KEYINPUT52), .A3(new_n847), .A4(new_n844), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n840), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT54), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n836), .A2(KEYINPUT116), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n831), .B2(new_n835), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n851), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n782), .A2(new_n786), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n747), .A2(new_n750), .A3(new_n837), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n787), .A2(KEYINPUT117), .A3(new_n839), .A4(new_n837), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n846), .A2(new_n847), .A3(new_n844), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT52), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n861), .A2(new_n862), .B1(new_n865), .B2(new_n848), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n857), .A2(new_n866), .B1(new_n850), .B2(new_n851), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n853), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n804), .A2(new_n686), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n872), .A2(new_n738), .A3(new_n760), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n651), .A3(new_n697), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT50), .Z(new_n875));
  NOR3_X1   g689(.A1(new_n789), .A2(new_n820), .A3(new_n488), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n804), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT119), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n826), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n819), .A2(new_n876), .ZN(new_n880));
  OR3_X1    g694(.A1(new_n880), .A2(new_n654), .A3(new_n663), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n875), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT51), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n872), .A2(new_n760), .A3(new_n809), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n820), .A2(new_n409), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n885), .B1(new_n814), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n886), .B(KEYINPUT118), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n814), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n890), .A2(new_n885), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n883), .B1(new_n882), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n878), .A2(new_n785), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT120), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT48), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n487), .B1(new_n880), .B2(new_n664), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n888), .A2(new_n892), .A3(new_n896), .A4(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n873), .A2(new_n690), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n870), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(G952), .A2(G953), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n824), .B1(new_n902), .B2(new_n903), .ZN(G75));
  INV_X1    g718(.A(new_n867), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(G210), .A3(G902), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n597), .A2(new_n615), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n611), .A2(new_n613), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n616), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT55), .Z(new_n912));
  AND3_X1   g726(.A1(new_n906), .A2(new_n907), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n906), .B2(new_n907), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n360), .A2(G952), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(G51));
  XNOR2_X1  g730(.A(new_n867), .B(new_n868), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n466), .B(KEYINPUT57), .Z(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n476), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n867), .A2(new_n358), .A3(new_n796), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n915), .B1(new_n920), .B2(new_n921), .ZN(G54));
  NAND4_X1  g736(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n923));
  INV_X1    g737(.A(new_n533), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n926), .A3(new_n915), .ZN(G60));
  INV_X1    g741(.A(new_n661), .ZN(new_n928));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT59), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n917), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n928), .B1(new_n870), .B2(new_n930), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n931), .A2(new_n932), .A3(new_n915), .ZN(G63));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n934));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT60), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n934), .B1(new_n867), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n936), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n861), .A2(new_n862), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n865), .A2(new_n848), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n857), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT53), .B1(new_n940), .B2(new_n840), .ZN(new_n942));
  OAI211_X1 g756(.A(KEYINPUT121), .B(new_n938), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n915), .B1(new_n944), .B2(new_n679), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n393), .A2(new_n396), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n937), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT123), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n937), .A2(new_n949), .A3(new_n946), .A4(new_n943), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n945), .A2(new_n948), .A3(KEYINPUT61), .A4(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT122), .B1(new_n944), .B2(new_n679), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT122), .ZN(new_n953));
  INV_X1    g767(.A(new_n679), .ZN(new_n954));
  AOI211_X1 g768(.A(new_n953), .B(new_n954), .C1(new_n937), .C2(new_n943), .ZN(new_n955));
  INV_X1    g769(.A(new_n915), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n947), .A2(new_n956), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n952), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n951), .B1(new_n958), .B2(KEYINPUT61), .ZN(G66));
  AOI21_X1  g773(.A(new_n360), .B1(new_n483), .B2(G224), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n860), .A2(new_n835), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(new_n360), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n908), .B1(G898), .B2(new_n360), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n962), .B(new_n963), .Z(G69));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n240), .A2(new_n252), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n519), .A2(new_n520), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n967), .B1(new_n366), .B2(new_n517), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n966), .B(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n360), .A2(G900), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n846), .A2(new_n847), .A3(new_n811), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n972), .A2(KEYINPUT126), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(KEYINPUT126), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n785), .A2(new_n801), .A3(new_n761), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n817), .A2(new_n976), .A3(new_n787), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n792), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n971), .B1(new_n978), .B2(new_n360), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n981));
  INV_X1    g795(.A(new_n792), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n973), .B2(new_n974), .ZN(new_n983));
  AOI21_X1  g797(.A(G953), .B1(new_n983), .B2(new_n977), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n981), .B1(new_n984), .B2(new_n971), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n970), .B1(new_n980), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n841), .ZN(new_n987));
  AND2_X1   g801(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n988));
  OR3_X1    g802(.A1(new_n721), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  XNOR2_X1  g803(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(new_n721), .B2(new_n987), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n817), .A2(new_n811), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n808), .A2(new_n714), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n744), .A2(new_n832), .A3(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n989), .A2(new_n991), .A3(new_n992), .A4(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n969), .A2(G953), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n965), .B1(new_n986), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n360), .B1(G227), .B2(G900), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n998), .B(new_n999), .ZN(G72));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT63), .Z(new_n1002));
  OAI211_X1 g816(.A(new_n281), .B(new_n1002), .C1(new_n995), .C2(new_n961), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n321), .B(new_n1002), .C1(new_n978), .C2(new_n961), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n1003), .A2(new_n306), .A3(new_n341), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n341), .A2(new_n306), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n852), .A2(new_n1002), .A3(new_n1006), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n1005), .A2(new_n956), .A3(new_n1007), .ZN(G57));
endmodule


