

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580;

  XNOR2_X1 U321 ( .A(n354), .B(n353), .ZN(n573) );
  AND2_X1 U322 ( .A1(G230GAT), .A2(G233GAT), .ZN(n289) );
  XOR2_X1 U323 ( .A(n351), .B(n350), .Z(n290) );
  NOR2_X1 U324 ( .A1(n358), .A2(n357), .ZN(n359) );
  XNOR2_X1 U325 ( .A(n426), .B(n289), .ZN(n343) );
  XNOR2_X1 U326 ( .A(n343), .B(n380), .ZN(n345) );
  XNOR2_X1 U327 ( .A(n352), .B(n290), .ZN(n353) );
  INV_X1 U328 ( .A(G218GAT), .ZN(n444) );
  XOR2_X1 U329 ( .A(n549), .B(KEYINPUT28), .Z(n520) );
  XNOR2_X1 U330 ( .A(n444), .B(KEYINPUT62), .ZN(n445) );
  XNOR2_X1 U331 ( .A(n446), .B(n445), .ZN(G1355GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT9), .B(KEYINPUT73), .Z(n292) );
  XNOR2_X1 U333 ( .A(G106GAT), .B(G92GAT), .ZN(n291) );
  XNOR2_X1 U334 ( .A(n292), .B(n291), .ZN(n309) );
  XOR2_X1 U335 ( .A(KEYINPUT10), .B(KEYINPUT64), .Z(n294) );
  XNOR2_X1 U336 ( .A(KEYINPUT74), .B(KEYINPUT11), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U338 ( .A(n295), .B(KEYINPUT76), .Z(n297) );
  XOR2_X1 U339 ( .A(G134GAT), .B(KEYINPUT75), .Z(n397) );
  XNOR2_X1 U340 ( .A(G218GAT), .B(n397), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n302) );
  XOR2_X1 U342 ( .A(G36GAT), .B(G190GAT), .Z(n373) );
  XNOR2_X1 U343 ( .A(G50GAT), .B(KEYINPUT72), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n298), .B(G162GAT), .ZN(n416) );
  XOR2_X1 U345 ( .A(n373), .B(n416), .Z(n300) );
  NAND2_X1 U346 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U348 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U349 ( .A(G29GAT), .B(G43GAT), .Z(n304) );
  XNOR2_X1 U350 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n327) );
  XNOR2_X1 U352 ( .A(G99GAT), .B(G85GAT), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n305), .B(KEYINPUT69), .ZN(n349) );
  XNOR2_X1 U354 ( .A(n327), .B(n349), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n564) );
  XNOR2_X1 U357 ( .A(KEYINPUT36), .B(n564), .ZN(n474) );
  XNOR2_X1 U358 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n367) );
  XOR2_X1 U359 ( .A(G155GAT), .B(G78GAT), .Z(n311) );
  XNOR2_X1 U360 ( .A(G22GAT), .B(G211GAT), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U362 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n313) );
  XNOR2_X1 U363 ( .A(G8GAT), .B(KEYINPUT77), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U365 ( .A(n315), .B(n314), .Z(n317) );
  XOR2_X1 U366 ( .A(G15GAT), .B(G1GAT), .Z(n338) );
  XOR2_X1 U367 ( .A(G57GAT), .B(KEYINPUT13), .Z(n344) );
  XNOR2_X1 U368 ( .A(n338), .B(n344), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U370 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n319) );
  NAND2_X1 U371 ( .A1(G231GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U373 ( .A(n321), .B(n320), .Z(n326) );
  XOR2_X1 U374 ( .A(G64GAT), .B(G127GAT), .Z(n323) );
  XNOR2_X1 U375 ( .A(G183GAT), .B(G71GAT), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n324), .B(KEYINPUT14), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n579) );
  NAND2_X1 U379 ( .A1(n579), .A2(n564), .ZN(n358) );
  XOR2_X1 U380 ( .A(G141GAT), .B(G22GAT), .Z(n412) );
  XNOR2_X1 U381 ( .A(n327), .B(n412), .ZN(n328) );
  XOR2_X1 U382 ( .A(G169GAT), .B(G8GAT), .Z(n374) );
  XNOR2_X1 U383 ( .A(n328), .B(n374), .ZN(n332) );
  XOR2_X1 U384 ( .A(KEYINPUT65), .B(KEYINPUT67), .Z(n330) );
  NAND2_X1 U385 ( .A1(G229GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U387 ( .A(n332), .B(n331), .Z(n337) );
  XOR2_X1 U388 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n334) );
  XNOR2_X1 U389 ( .A(G197GAT), .B(G113GAT), .ZN(n333) );
  XNOR2_X1 U390 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n335), .B(KEYINPUT30), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n339) );
  XOR2_X1 U393 ( .A(n339), .B(n338), .Z(n341) );
  XNOR2_X1 U394 ( .A(G36GAT), .B(G50GAT), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n568) );
  XOR2_X1 U396 ( .A(G120GAT), .B(G71GAT), .Z(n426) );
  XNOR2_X1 U397 ( .A(G176GAT), .B(G92GAT), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n342), .B(G64GAT), .ZN(n380) );
  XOR2_X1 U399 ( .A(n345), .B(n344), .Z(n347) );
  XNOR2_X1 U400 ( .A(G204GAT), .B(KEYINPUT70), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n354) );
  XNOR2_X1 U402 ( .A(G106GAT), .B(G78GAT), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n348), .B(G148GAT), .ZN(n421) );
  XNOR2_X1 U404 ( .A(n421), .B(n349), .ZN(n352) );
  XOR2_X1 U405 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n351) );
  XNOR2_X1 U406 ( .A(KEYINPUT32), .B(KEYINPUT68), .ZN(n350) );
  INV_X1 U407 ( .A(KEYINPUT41), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n573), .B(n355), .ZN(n556) );
  NOR2_X1 U409 ( .A1(n568), .A2(n556), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n356), .B(KEYINPUT46), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n359), .B(KEYINPUT47), .ZN(n365) );
  NOR2_X1 U412 ( .A1(n474), .A2(n579), .ZN(n360) );
  XNOR2_X1 U413 ( .A(KEYINPUT45), .B(n360), .ZN(n361) );
  NAND2_X1 U414 ( .A1(n361), .A2(n573), .ZN(n362) );
  XOR2_X1 U415 ( .A(KEYINPUT110), .B(n362), .Z(n363) );
  NAND2_X1 U416 ( .A1(n363), .A2(n568), .ZN(n364) );
  NAND2_X1 U417 ( .A1(n365), .A2(n364), .ZN(n366) );
  XNOR2_X1 U418 ( .A(n367), .B(n366), .ZN(n518) );
  XOR2_X1 U419 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n369) );
  XNOR2_X1 U420 ( .A(G218GAT), .B(KEYINPUT86), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U422 ( .A(n370), .B(G211GAT), .Z(n372) );
  XNOR2_X1 U423 ( .A(G197GAT), .B(G204GAT), .ZN(n371) );
  XNOR2_X1 U424 ( .A(n372), .B(n371), .ZN(n422) );
  XNOR2_X1 U425 ( .A(n374), .B(n373), .ZN(n384) );
  XOR2_X1 U426 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n376) );
  NAND2_X1 U427 ( .A1(G226GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U428 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U429 ( .A(n377), .B(KEYINPUT92), .Z(n382) );
  XOR2_X1 U430 ( .A(G183GAT), .B(KEYINPUT18), .Z(n379) );
  XNOR2_X1 U431 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n378) );
  XNOR2_X1 U432 ( .A(n379), .B(n378), .ZN(n430) );
  XNOR2_X1 U433 ( .A(n430), .B(n380), .ZN(n381) );
  XNOR2_X1 U434 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U435 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U436 ( .A(n422), .B(n385), .ZN(n510) );
  NOR2_X1 U437 ( .A1(n518), .A2(n510), .ZN(n386) );
  XNOR2_X1 U438 ( .A(n386), .B(KEYINPUT54), .ZN(n408) );
  XOR2_X1 U439 ( .A(KEYINPUT88), .B(KEYINPUT6), .Z(n388) );
  XNOR2_X1 U440 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n388), .B(n387), .ZN(n407) );
  XOR2_X1 U442 ( .A(KEYINPUT5), .B(G57GAT), .Z(n390) );
  XNOR2_X1 U443 ( .A(G141GAT), .B(G120GAT), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U445 ( .A(G85GAT), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U446 ( .A(G29GAT), .B(G148GAT), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n405) );
  XOR2_X1 U449 ( .A(G127GAT), .B(KEYINPUT0), .Z(n396) );
  XNOR2_X1 U450 ( .A(G113GAT), .B(KEYINPUT80), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n425) );
  XOR2_X1 U452 ( .A(n397), .B(n425), .Z(n399) );
  NAND2_X1 U453 ( .A1(G225GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U455 ( .A(n400), .B(KEYINPUT89), .Z(n403) );
  XNOR2_X1 U456 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n401), .B(KEYINPUT3), .ZN(n419) );
  XNOR2_X1 U458 ( .A(G1GAT), .B(n419), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n407), .B(n406), .ZN(n507) );
  NAND2_X1 U462 ( .A1(n408), .A2(n507), .ZN(n548) );
  XOR2_X1 U463 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n442) );
  XOR2_X1 U464 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n410) );
  XNOR2_X1 U465 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U467 ( .A(n412), .B(n411), .Z(n414) );
  NAND2_X1 U468 ( .A1(G228GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U470 ( .A(n415), .B(KEYINPUT24), .Z(n418) );
  XNOR2_X1 U471 ( .A(n416), .B(KEYINPUT87), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U473 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U474 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U475 ( .A(n424), .B(n423), .ZN(n549) );
  XOR2_X1 U476 ( .A(n426), .B(n425), .Z(n428) );
  NAND2_X1 U477 ( .A1(G227GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U478 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U479 ( .A(n429), .B(G176GAT), .Z(n432) );
  XNOR2_X1 U480 ( .A(G169GAT), .B(n430), .ZN(n431) );
  XNOR2_X1 U481 ( .A(n432), .B(n431), .ZN(n440) );
  XOR2_X1 U482 ( .A(G134GAT), .B(G99GAT), .Z(n434) );
  XNOR2_X1 U483 ( .A(G43GAT), .B(G190GAT), .ZN(n433) );
  XNOR2_X1 U484 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U485 ( .A(KEYINPUT81), .B(KEYINPUT20), .Z(n436) );
  XNOR2_X1 U486 ( .A(G15GAT), .B(KEYINPUT82), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U488 ( .A(n438), .B(n437), .Z(n439) );
  XNOR2_X1 U489 ( .A(n440), .B(n439), .ZN(n552) );
  INV_X1 U490 ( .A(n552), .ZN(n522) );
  NAND2_X1 U491 ( .A1(n549), .A2(n522), .ZN(n441) );
  XNOR2_X1 U492 ( .A(n442), .B(n441), .ZN(n536) );
  NOR2_X1 U493 ( .A1(n548), .A2(n536), .ZN(n443) );
  XOR2_X1 U494 ( .A(KEYINPUT124), .B(n443), .Z(n578) );
  NOR2_X1 U495 ( .A1(n474), .A2(n578), .ZN(n446) );
  INV_X1 U496 ( .A(n568), .ZN(n490) );
  NAND2_X1 U497 ( .A1(n490), .A2(n573), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n447), .B(KEYINPUT71), .ZN(n477) );
  INV_X1 U499 ( .A(n507), .ZN(n493) );
  NOR2_X1 U500 ( .A1(n522), .A2(n510), .ZN(n448) );
  NOR2_X1 U501 ( .A1(n549), .A2(n448), .ZN(n449) );
  XOR2_X1 U502 ( .A(KEYINPUT25), .B(n449), .Z(n452) );
  XOR2_X1 U503 ( .A(KEYINPUT27), .B(KEYINPUT93), .Z(n450) );
  XNOR2_X1 U504 ( .A(n510), .B(n450), .ZN(n454) );
  NOR2_X1 U505 ( .A1(n536), .A2(n454), .ZN(n451) );
  NOR2_X1 U506 ( .A1(n452), .A2(n451), .ZN(n453) );
  NOR2_X1 U507 ( .A1(n493), .A2(n453), .ZN(n458) );
  NOR2_X1 U508 ( .A1(n454), .A2(n507), .ZN(n455) );
  XOR2_X1 U509 ( .A(KEYINPUT94), .B(n455), .Z(n519) );
  NAND2_X1 U510 ( .A1(n522), .A2(n520), .ZN(n456) );
  NOR2_X1 U511 ( .A1(n519), .A2(n456), .ZN(n457) );
  NOR2_X1 U512 ( .A1(n458), .A2(n457), .ZN(n473) );
  INV_X1 U513 ( .A(n579), .ZN(n459) );
  NAND2_X1 U514 ( .A1(n564), .A2(n459), .ZN(n460) );
  XNOR2_X1 U515 ( .A(KEYINPUT16), .B(n460), .ZN(n461) );
  NOR2_X1 U516 ( .A1(n473), .A2(n461), .ZN(n491) );
  NAND2_X1 U517 ( .A1(n477), .A2(n491), .ZN(n470) );
  NOR2_X1 U518 ( .A1(n507), .A2(n470), .ZN(n463) );
  XNOR2_X1 U519 ( .A(KEYINPUT34), .B(KEYINPUT96), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U521 ( .A(G1GAT), .B(n464), .Z(G1324GAT) );
  NOR2_X1 U522 ( .A1(n510), .A2(n470), .ZN(n466) );
  XNOR2_X1 U523 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U525 ( .A(G8GAT), .B(n467), .ZN(G1325GAT) );
  NOR2_X1 U526 ( .A1(n522), .A2(n470), .ZN(n469) );
  XNOR2_X1 U527 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n469), .B(n468), .ZN(G1326GAT) );
  NOR2_X1 U529 ( .A1(n520), .A2(n470), .ZN(n472) );
  XNOR2_X1 U530 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(G1327GAT) );
  NOR2_X1 U532 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U533 ( .A1(n579), .A2(n475), .ZN(n476) );
  XNOR2_X1 U534 ( .A(KEYINPUT37), .B(n476), .ZN(n506) );
  NAND2_X1 U535 ( .A1(n477), .A2(n506), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n478), .B(KEYINPUT38), .ZN(n487) );
  NOR2_X1 U537 ( .A1(n507), .A2(n487), .ZN(n482) );
  XOR2_X1 U538 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n480) );
  XNOR2_X1 U539 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(G1328GAT) );
  NOR2_X1 U542 ( .A1(n487), .A2(n510), .ZN(n483) );
  XOR2_X1 U543 ( .A(KEYINPUT102), .B(n483), .Z(n484) );
  XNOR2_X1 U544 ( .A(G36GAT), .B(n484), .ZN(G1329GAT) );
  NOR2_X1 U545 ( .A1(n522), .A2(n487), .ZN(n485) );
  XOR2_X1 U546 ( .A(KEYINPUT40), .B(n485), .Z(n486) );
  XNOR2_X1 U547 ( .A(G43GAT), .B(n486), .ZN(G1330GAT) );
  XNOR2_X1 U548 ( .A(G50GAT), .B(KEYINPUT103), .ZN(n489) );
  NOR2_X1 U549 ( .A1(n520), .A2(n487), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(G1331GAT) );
  NOR2_X1 U551 ( .A1(n556), .A2(n490), .ZN(n505) );
  NAND2_X1 U552 ( .A1(n491), .A2(n505), .ZN(n492) );
  XOR2_X1 U553 ( .A(KEYINPUT104), .B(n492), .Z(n502) );
  NAND2_X1 U554 ( .A1(n502), .A2(n493), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n494), .B(KEYINPUT42), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G57GAT), .B(n495), .ZN(G1332GAT) );
  INV_X1 U557 ( .A(n510), .ZN(n496) );
  NAND2_X1 U558 ( .A1(n496), .A2(n502), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G64GAT), .B(n497), .ZN(G1333GAT) );
  NAND2_X1 U560 ( .A1(n502), .A2(n552), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n498), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n500) );
  XNOR2_X1 U563 ( .A(G78GAT), .B(KEYINPUT106), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(n504) );
  INV_X1 U565 ( .A(n520), .ZN(n501) );
  NAND2_X1 U566 ( .A1(n502), .A2(n501), .ZN(n503) );
  XOR2_X1 U567 ( .A(n504), .B(n503), .Z(G1335GAT) );
  NAND2_X1 U568 ( .A1(n506), .A2(n505), .ZN(n514) );
  NOR2_X1 U569 ( .A1(n507), .A2(n514), .ZN(n509) );
  XNOR2_X1 U570 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n509), .B(n508), .ZN(G1336GAT) );
  NOR2_X1 U572 ( .A1(n510), .A2(n514), .ZN(n511) );
  XOR2_X1 U573 ( .A(KEYINPUT108), .B(n511), .Z(n512) );
  XNOR2_X1 U574 ( .A(G92GAT), .B(n512), .ZN(G1337GAT) );
  NOR2_X1 U575 ( .A1(n522), .A2(n514), .ZN(n513) );
  XOR2_X1 U576 ( .A(G99GAT), .B(n513), .Z(G1338GAT) );
  NOR2_X1 U577 ( .A1(n520), .A2(n514), .ZN(n516) );
  XNOR2_X1 U578 ( .A(KEYINPUT44), .B(KEYINPUT109), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U580 ( .A(G106GAT), .B(n517), .ZN(G1339GAT) );
  XNOR2_X1 U581 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n525) );
  NOR2_X1 U582 ( .A1(n519), .A2(n518), .ZN(n537) );
  NAND2_X1 U583 ( .A1(n537), .A2(n520), .ZN(n521) );
  NOR2_X1 U584 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U585 ( .A(KEYINPUT112), .B(n523), .Z(n532) );
  NOR2_X1 U586 ( .A1(n568), .A2(n532), .ZN(n524) );
  XNOR2_X1 U587 ( .A(n525), .B(n524), .ZN(G1340GAT) );
  NOR2_X1 U588 ( .A1(n532), .A2(n556), .ZN(n529) );
  XOR2_X1 U589 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n527) );
  XNOR2_X1 U590 ( .A(G120GAT), .B(KEYINPUT115), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n529), .B(n528), .ZN(G1341GAT) );
  NOR2_X1 U593 ( .A1(n579), .A2(n532), .ZN(n530) );
  XOR2_X1 U594 ( .A(KEYINPUT50), .B(n530), .Z(n531) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(n531), .ZN(G1342GAT) );
  NOR2_X1 U596 ( .A1(n532), .A2(n564), .ZN(n534) );
  XNOR2_X1 U597 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G134GAT), .B(n535), .ZN(G1343GAT) );
  INV_X1 U600 ( .A(n536), .ZN(n538) );
  NAND2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U602 ( .A(KEYINPUT117), .B(n539), .Z(n545) );
  NOR2_X1 U603 ( .A1(n568), .A2(n545), .ZN(n540) );
  XOR2_X1 U604 ( .A(G141GAT), .B(n540), .Z(G1344GAT) );
  NOR2_X1 U605 ( .A1(n556), .A2(n545), .ZN(n542) );
  XNOR2_X1 U606 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(n543), .ZN(G1345GAT) );
  NOR2_X1 U609 ( .A1(n579), .A2(n545), .ZN(n544) );
  XOR2_X1 U610 ( .A(G155GAT), .B(n544), .Z(G1346GAT) );
  NOR2_X1 U611 ( .A1(n564), .A2(n545), .ZN(n546) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(n546), .Z(n547) );
  XNOR2_X1 U613 ( .A(G162GAT), .B(n547), .ZN(G1347GAT) );
  NOR2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U615 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n563) );
  NOR2_X1 U618 ( .A1(n568), .A2(n563), .ZN(n554) );
  XOR2_X1 U619 ( .A(G169GAT), .B(n554), .Z(n555) );
  XNOR2_X1 U620 ( .A(KEYINPUT120), .B(n555), .ZN(G1348GAT) );
  NOR2_X1 U621 ( .A1(n556), .A2(n563), .ZN(n561) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n558) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(KEYINPUT121), .B(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NOR2_X1 U627 ( .A1(n579), .A2(n563), .ZN(n562) );
  XOR2_X1 U628 ( .A(G183GAT), .B(n562), .Z(G1350GAT) );
  NOR2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n566) );
  XNOR2_X1 U630 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(n567), .ZN(G1351GAT) );
  NOR2_X1 U633 ( .A1(n578), .A2(n568), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n578), .A2(n573), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n575) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT127), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
endmodule

