

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745;

  NOR2_X1 U369 ( .A1(G953), .A2(G237), .ZN(n463) );
  NOR2_X1 U370 ( .A1(n523), .A2(n615), .ZN(n620) );
  NAND2_X1 U371 ( .A1(n620), .A2(n546), .ZN(n593) );
  OR2_X2 U372 ( .A1(n662), .A2(n414), .ZN(n413) );
  OR2_X1 U373 ( .A1(n574), .A2(n573), .ZN(n406) );
  XNOR2_X1 U374 ( .A(n352), .B(KEYINPUT103), .ZN(n634) );
  XNOR2_X1 U375 ( .A(n592), .B(KEYINPUT6), .ZN(n519) );
  XNOR2_X1 U376 ( .A(n540), .B(n487), .ZN(n619) );
  INV_X1 U377 ( .A(G953), .ZN(n735) );
  AND2_X2 U378 ( .A1(n718), .A2(n734), .ZN(n658) );
  XNOR2_X2 U379 ( .A(n726), .B(n503), .ZN(n662) );
  XNOR2_X2 U380 ( .A(n494), .B(n493), .ZN(n726) );
  NAND2_X1 U381 ( .A1(n366), .A2(n362), .ZN(n361) );
  NOR2_X1 U382 ( .A1(n579), .A2(KEYINPUT48), .ZN(n362) );
  XNOR2_X1 U383 ( .A(n460), .B(n347), .ZN(n479) );
  XNOR2_X1 U384 ( .A(n421), .B(G125), .ZN(n498) );
  NAND2_X1 U385 ( .A1(n504), .A2(n415), .ZN(n414) );
  INV_X1 U386 ( .A(n506), .ZN(n415) );
  NAND2_X1 U387 ( .A1(n453), .A2(G221), .ZN(n403) );
  XNOR2_X1 U388 ( .A(n482), .B(n481), .ZN(n493) );
  XNOR2_X1 U389 ( .A(G101), .B(KEYINPUT89), .ZN(n481) );
  XNOR2_X1 U390 ( .A(G107), .B(G104), .ZN(n480) );
  INV_X1 U391 ( .A(KEYINPUT83), .ZN(n411) );
  NAND2_X1 U392 ( .A1(n386), .A2(n351), .ZN(n385) );
  NAND2_X1 U393 ( .A1(n659), .A2(n506), .ZN(n416) );
  NOR2_X1 U394 ( .A1(n363), .A2(n365), .ZN(n611) );
  NAND2_X1 U395 ( .A1(n361), .A2(n360), .ZN(n363) );
  XNOR2_X1 U396 ( .A(n388), .B(n410), .ZN(n609) );
  XNOR2_X1 U397 ( .A(n486), .B(G469), .ZN(n540) );
  NOR2_X1 U398 ( .A1(G902), .A2(n683), .ZN(n486) );
  NOR2_X1 U399 ( .A1(G902), .A2(n671), .ZN(n474) );
  XNOR2_X1 U400 ( .A(n372), .B(n369), .ZN(n404) );
  XNOR2_X1 U401 ( .A(n424), .B(n373), .ZN(n372) );
  XNOR2_X1 U402 ( .A(n371), .B(n370), .ZN(n369) );
  XNOR2_X1 U403 ( .A(KEYINPUT93), .B(KEYINPUT23), .ZN(n424) );
  XNOR2_X1 U404 ( .A(n392), .B(n423), .ZN(n453) );
  XOR2_X1 U405 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n423) );
  NAND2_X1 U406 ( .A1(n394), .A2(n393), .ZN(n392) );
  XOR2_X1 U407 ( .A(KEYINPUT10), .B(n498), .Z(n733) );
  XOR2_X1 U408 ( .A(G113), .B(G104), .Z(n467) );
  XNOR2_X1 U409 ( .A(n468), .B(n353), .ZN(n469) );
  XNOR2_X1 U410 ( .A(G143), .B(G140), .ZN(n468) );
  XNOR2_X1 U411 ( .A(n354), .B(KEYINPUT11), .ZN(n353) );
  INV_X1 U412 ( .A(KEYINPUT12), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n479), .B(n478), .ZN(n732) );
  XNOR2_X1 U414 ( .A(n358), .B(n553), .ZN(n581) );
  XNOR2_X1 U415 ( .A(n517), .B(KEYINPUT22), .ZN(n533) );
  OR2_X1 U416 ( .A1(n714), .A2(G902), .ZN(n368) );
  INV_X1 U417 ( .A(KEYINPUT25), .ZN(n429) );
  INV_X1 U418 ( .A(n519), .ZN(n530) );
  AND2_X1 U419 ( .A1(n364), .A2(n348), .ZN(n360) );
  NAND2_X1 U420 ( .A1(n579), .A2(KEYINPUT48), .ZN(n364) );
  INV_X1 U421 ( .A(KEYINPUT46), .ZN(n367) );
  NAND2_X1 U422 ( .A1(n374), .A2(n389), .ZN(n388) );
  AND2_X1 U423 ( .A1(n601), .A2(n602), .ZN(n389) );
  XNOR2_X1 U424 ( .A(n375), .B(n411), .ZN(n374) );
  INV_X1 U425 ( .A(KEYINPUT82), .ZN(n410) );
  NAND2_X1 U426 ( .A1(G237), .A2(G234), .ZN(n433) );
  XOR2_X1 U427 ( .A(G137), .B(KEYINPUT5), .Z(n440) );
  XOR2_X1 U428 ( .A(G146), .B(G101), .Z(n419) );
  XNOR2_X1 U429 ( .A(G128), .B(KEYINPUT94), .ZN(n370) );
  XNOR2_X1 U430 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n371) );
  XNOR2_X1 U431 ( .A(KEYINPUT77), .B(KEYINPUT72), .ZN(n373) );
  NOR2_X1 U432 ( .A1(KEYINPUT78), .A2(G953), .ZN(n390) );
  AND2_X1 U433 ( .A1(n396), .A2(n395), .ZN(n394) );
  NAND2_X1 U434 ( .A1(KEYINPUT78), .A2(G953), .ZN(n395) );
  NAND2_X1 U435 ( .A1(n391), .A2(KEYINPUT78), .ZN(n396) );
  INV_X1 U436 ( .A(G234), .ZN(n391) );
  XNOR2_X1 U437 ( .A(n447), .B(G128), .ZN(n500) );
  INV_X1 U438 ( .A(G143), .ZN(n447) );
  XNOR2_X1 U439 ( .A(KEYINPUT73), .B(KEYINPUT4), .ZN(n499) );
  NAND2_X1 U440 ( .A1(n382), .A2(n588), .ZN(n381) );
  INV_X1 U441 ( .A(G237), .ZN(n488) );
  XNOR2_X1 U442 ( .A(n401), .B(KEYINPUT67), .ZN(n539) );
  NAND2_X1 U443 ( .A1(n539), .A2(n592), .ZN(n400) );
  AND2_X1 U444 ( .A1(n526), .A2(n569), .ZN(n352) );
  XNOR2_X1 U445 ( .A(n452), .B(n451), .ZN(n547) );
  XNOR2_X1 U446 ( .A(n450), .B(n449), .ZN(n451) );
  INV_X1 U447 ( .A(G472), .ZN(n449) );
  XNOR2_X1 U448 ( .A(n611), .B(n583), .ZN(n734) );
  INV_X1 U449 ( .A(KEYINPUT79), .ZN(n583) );
  XNOR2_X1 U450 ( .A(n444), .B(n443), .ZN(n376) );
  XNOR2_X1 U451 ( .A(G116), .B(G113), .ZN(n444) );
  XNOR2_X1 U452 ( .A(KEYINPUT3), .B(G119), .ZN(n443) );
  XNOR2_X1 U453 ( .A(G107), .B(G122), .ZN(n454) );
  XOR2_X1 U454 ( .A(KEYINPUT9), .B(G116), .Z(n455) );
  XNOR2_X1 U455 ( .A(n500), .B(n387), .ZN(n460) );
  INV_X1 U456 ( .A(G134), .ZN(n387) );
  XNOR2_X1 U457 ( .A(n613), .B(n612), .ZN(n379) );
  INV_X1 U458 ( .A(KEYINPUT80), .ZN(n612) );
  NAND2_X1 U459 ( .A1(n412), .A2(n417), .ZN(n377) );
  AND2_X1 U460 ( .A1(n413), .A2(n350), .ZN(n412) );
  XNOR2_X1 U461 ( .A(n359), .B(KEYINPUT71), .ZN(n567) );
  NAND2_X1 U462 ( .A1(n552), .A2(n418), .ZN(n359) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n569) );
  XNOR2_X1 U464 ( .A(n462), .B(G478), .ZN(n397) );
  OR2_X1 U465 ( .A1(n710), .A2(G902), .ZN(n398) );
  INV_X1 U466 ( .A(KEYINPUT102), .ZN(n462) );
  XNOR2_X1 U467 ( .A(n376), .B(n492), .ZN(n494) );
  XNOR2_X1 U468 ( .A(KEYINPUT16), .B(G122), .ZN(n492) );
  XNOR2_X1 U469 ( .A(n422), .B(n733), .ZN(n425) );
  XNOR2_X1 U470 ( .A(n404), .B(n403), .ZN(n402) );
  XNOR2_X1 U471 ( .A(n461), .B(n460), .ZN(n710) );
  XNOR2_X1 U472 ( .A(n459), .B(n458), .ZN(n461) );
  NAND2_X1 U473 ( .A1(n453), .A2(G217), .ZN(n459) );
  XNOR2_X1 U474 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U475 ( .A(n471), .B(n472), .ZN(n473) );
  BUF_X1 U476 ( .A(n681), .Z(n713) );
  XNOR2_X1 U477 ( .A(n732), .B(n485), .ZN(n683) );
  AND2_X1 U478 ( .A1(n665), .A2(G953), .ZN(n717) );
  XNOR2_X1 U479 ( .A(n535), .B(n534), .ZN(n587) );
  NOR2_X1 U480 ( .A1(n533), .A2(n532), .ZN(n535) );
  INV_X1 U481 ( .A(n406), .ZN(n405) );
  XOR2_X1 U482 ( .A(n430), .B(n429), .Z(n346) );
  XOR2_X1 U483 ( .A(G131), .B(KEYINPUT4), .Z(n347) );
  NAND2_X1 U484 ( .A1(n619), .A2(n620), .ZN(n386) );
  INV_X1 U485 ( .A(n386), .ZN(n588) );
  AND2_X1 U486 ( .A1(n709), .A2(n582), .ZN(n348) );
  AND2_X1 U487 ( .A1(n413), .A2(n416), .ZN(n349) );
  AND2_X1 U488 ( .A1(n416), .A2(n630), .ZN(n350) );
  XOR2_X1 U489 ( .A(n524), .B(KEYINPUT33), .Z(n351) );
  XNOR2_X1 U490 ( .A(n425), .B(n402), .ZN(n714) );
  NAND2_X1 U491 ( .A1(n390), .A2(G234), .ZN(n393) );
  NOR2_X2 U492 ( .A1(n573), .A2(n513), .ZN(n356) );
  XNOR2_X1 U493 ( .A(n355), .B(n680), .ZN(G57) );
  NOR2_X2 U494 ( .A1(n679), .A2(n717), .ZN(n355) );
  XNOR2_X2 U495 ( .A(n356), .B(n514), .ZN(n589) );
  XNOR2_X2 U496 ( .A(n357), .B(KEYINPUT45), .ZN(n718) );
  NAND2_X1 U497 ( .A1(n609), .A2(n608), .ZN(n357) );
  NAND2_X1 U498 ( .A1(n567), .A2(n631), .ZN(n358) );
  XNOR2_X1 U499 ( .A(n556), .B(n367), .ZN(n366) );
  NOR2_X1 U500 ( .A1(n366), .A2(n580), .ZN(n365) );
  XNOR2_X2 U501 ( .A(n368), .B(n346), .ZN(n523) );
  NAND2_X1 U502 ( .A1(n603), .A2(KEYINPUT44), .ZN(n375) );
  XNOR2_X1 U503 ( .A(n528), .B(KEYINPUT35), .ZN(n603) );
  XNOR2_X1 U504 ( .A(n376), .B(n419), .ZN(n445) );
  XNOR2_X2 U505 ( .A(n559), .B(KEYINPUT19), .ZN(n573) );
  XNOR2_X2 U506 ( .A(n377), .B(n509), .ZN(n559) );
  NOR2_X4 U507 ( .A1(n380), .A2(n378), .ZN(n681) );
  NAND2_X1 U508 ( .A1(n660), .A2(n659), .ZN(n378) );
  NAND2_X1 U509 ( .A1(n718), .A2(n379), .ZN(n660) );
  NOR2_X2 U510 ( .A1(n658), .A2(KEYINPUT2), .ZN(n380) );
  NAND2_X1 U511 ( .A1(n383), .A2(n381), .ZN(n409) );
  NOR2_X1 U512 ( .A1(n519), .A2(n351), .ZN(n382) );
  AND2_X1 U513 ( .A1(n385), .A2(n384), .ZN(n383) );
  NAND2_X1 U514 ( .A1(n519), .A2(n351), .ZN(n384) );
  INV_X1 U515 ( .A(n409), .ZN(n648) );
  NOR2_X2 U516 ( .A1(n666), .A2(n717), .ZN(n668) );
  NOR2_X2 U517 ( .A1(n674), .A2(n717), .ZN(n675) );
  XNOR2_X1 U518 ( .A(n400), .B(n399), .ZN(n542) );
  INV_X1 U519 ( .A(KEYINPUT28), .ZN(n399) );
  NAND2_X1 U520 ( .A1(n523), .A2(n439), .ZN(n401) );
  NAND2_X1 U521 ( .A1(n405), .A2(n636), .ZN(n575) );
  NAND2_X1 U522 ( .A1(n405), .A2(n693), .ZN(n694) );
  NAND2_X1 U523 ( .A1(n405), .A2(n697), .ZN(n698) );
  XNOR2_X1 U524 ( .A(n406), .B(KEYINPUT47), .ZN(n576) );
  NAND2_X1 U525 ( .A1(n407), .A2(n527), .ZN(n528) );
  XNOR2_X1 U526 ( .A(n408), .B(n525), .ZN(n407) );
  NAND2_X1 U527 ( .A1(n595), .A2(n409), .ZN(n408) );
  XNOR2_X1 U528 ( .A(n589), .B(KEYINPUT91), .ZN(n595) );
  NAND2_X1 U529 ( .A1(n417), .A2(n349), .ZN(n536) );
  NAND2_X1 U530 ( .A1(n662), .A2(n506), .ZN(n417) );
  BUF_X1 U531 ( .A(n603), .Z(n605) );
  AND2_X1 U532 ( .A1(n551), .A2(n550), .ZN(n418) );
  INV_X1 U533 ( .A(KEYINPUT48), .ZN(n580) );
  XNOR2_X1 U534 ( .A(n420), .B(G119), .ZN(n422) );
  XNOR2_X1 U535 ( .A(n446), .B(n445), .ZN(n448) );
  INV_X1 U536 ( .A(n477), .ZN(n478) );
  INV_X1 U537 ( .A(n533), .ZN(n586) );
  XNOR2_X1 U538 ( .A(G140), .B(G137), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n477), .B(G110), .ZN(n420) );
  INV_X1 U540 ( .A(G146), .ZN(n421) );
  XOR2_X1 U541 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n428) );
  XNOR2_X1 U542 ( .A(KEYINPUT88), .B(KEYINPUT15), .ZN(n426) );
  XNOR2_X1 U543 ( .A(n426), .B(G902), .ZN(n504) );
  NAND2_X1 U544 ( .A1(n504), .A2(G234), .ZN(n427) );
  XNOR2_X1 U545 ( .A(n428), .B(n427), .ZN(n431) );
  NAND2_X1 U546 ( .A1(G217), .A2(n431), .ZN(n430) );
  NAND2_X1 U547 ( .A1(G221), .A2(n431), .ZN(n432) );
  XNOR2_X1 U548 ( .A(KEYINPUT21), .B(n432), .ZN(n615) );
  XNOR2_X1 U549 ( .A(n433), .B(KEYINPUT14), .ZN(n434) );
  XNOR2_X1 U550 ( .A(KEYINPUT70), .B(n434), .ZN(n435) );
  NAND2_X1 U551 ( .A1(G952), .A2(n435), .ZN(n646) );
  NOR2_X1 U552 ( .A1(n646), .A2(G953), .ZN(n512) );
  NAND2_X1 U553 ( .A1(G902), .A2(n435), .ZN(n510) );
  OR2_X1 U554 ( .A1(n735), .A2(n510), .ZN(n436) );
  XNOR2_X1 U555 ( .A(KEYINPUT106), .B(n436), .ZN(n437) );
  NOR2_X1 U556 ( .A1(G900), .A2(n437), .ZN(n438) );
  NOR2_X1 U557 ( .A1(n512), .A2(n438), .ZN(n549) );
  NOR2_X1 U558 ( .A1(n615), .A2(n549), .ZN(n439) );
  NAND2_X1 U559 ( .A1(G210), .A2(n463), .ZN(n441) );
  XNOR2_X1 U560 ( .A(n440), .B(n441), .ZN(n442) );
  XOR2_X1 U561 ( .A(n442), .B(KEYINPUT96), .Z(n446) );
  XNOR2_X1 U562 ( .A(n448), .B(n479), .ZN(n676) );
  NOR2_X1 U563 ( .A1(G902), .A2(n676), .ZN(n452) );
  INV_X1 U564 ( .A(KEYINPUT97), .ZN(n450) );
  INV_X1 U565 ( .A(n547), .ZN(n618) );
  INV_X1 U566 ( .A(n618), .ZN(n592) );
  XNOR2_X1 U567 ( .A(n455), .B(n454), .ZN(n457) );
  XNOR2_X1 U568 ( .A(KEYINPUT101), .B(KEYINPUT7), .ZN(n456) );
  XNOR2_X1 U569 ( .A(KEYINPUT13), .B(G475), .ZN(n475) );
  XOR2_X1 U570 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n465) );
  NAND2_X1 U571 ( .A1(n463), .A2(G214), .ZN(n464) );
  XNOR2_X1 U572 ( .A(n465), .B(n464), .ZN(n472) );
  XNOR2_X1 U573 ( .A(G122), .B(G131), .ZN(n466) );
  XNOR2_X1 U574 ( .A(n467), .B(n466), .ZN(n470) );
  XOR2_X1 U575 ( .A(n470), .B(n469), .Z(n471) );
  XNOR2_X1 U576 ( .A(n733), .B(n473), .ZN(n671) );
  XOR2_X1 U577 ( .A(n475), .B(n474), .Z(n526) );
  INV_X1 U578 ( .A(n526), .ZN(n568) );
  NAND2_X1 U579 ( .A1(n569), .A2(n568), .ZN(n699) );
  NOR2_X1 U580 ( .A1(n519), .A2(n699), .ZN(n476) );
  NAND2_X1 U581 ( .A1(n539), .A2(n476), .ZN(n558) );
  XNOR2_X1 U582 ( .A(n480), .B(G110), .ZN(n482) );
  NAND2_X1 U583 ( .A1(G227), .A2(n735), .ZN(n483) );
  XNOR2_X1 U584 ( .A(n483), .B(G146), .ZN(n484) );
  XNOR2_X1 U585 ( .A(n493), .B(n484), .ZN(n485) );
  INV_X1 U586 ( .A(KEYINPUT1), .ZN(n487) );
  INV_X1 U587 ( .A(n619), .ZN(n518) );
  INV_X1 U588 ( .A(G902), .ZN(n489) );
  NAND2_X1 U589 ( .A1(n489), .A2(n488), .ZN(n505) );
  NAND2_X1 U590 ( .A1(n505), .A2(G214), .ZN(n630) );
  NAND2_X1 U591 ( .A1(n518), .A2(n630), .ZN(n490) );
  NOR2_X1 U592 ( .A1(n558), .A2(n490), .ZN(n491) );
  XNOR2_X1 U593 ( .A(n491), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U594 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n496) );
  NAND2_X1 U595 ( .A1(n735), .A2(G224), .ZN(n495) );
  XNOR2_X1 U596 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U597 ( .A(n498), .B(n497), .ZN(n502) );
  XNOR2_X1 U598 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U599 ( .A(n502), .B(n501), .ZN(n503) );
  INV_X1 U600 ( .A(n504), .ZN(n659) );
  NAND2_X1 U601 ( .A1(n505), .A2(G210), .ZN(n506) );
  INV_X1 U602 ( .A(n536), .ZN(n564) );
  OR2_X1 U603 ( .A1(n507), .A2(n564), .ZN(n582) );
  XNOR2_X1 U604 ( .A(n582), .B(G140), .ZN(G42) );
  NOR2_X1 U605 ( .A1(n634), .A2(n615), .ZN(n508) );
  XNOR2_X1 U606 ( .A(n508), .B(KEYINPUT104), .ZN(n516) );
  INV_X1 U607 ( .A(KEYINPUT84), .ZN(n509) );
  XOR2_X1 U608 ( .A(G898), .B(KEYINPUT90), .Z(n722) );
  NAND2_X1 U609 ( .A1(G953), .A2(n722), .ZN(n728) );
  NOR2_X1 U610 ( .A1(n510), .A2(n728), .ZN(n511) );
  NOR2_X1 U611 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U612 ( .A(KEYINPUT85), .B(KEYINPUT0), .ZN(n514) );
  INV_X1 U613 ( .A(n589), .ZN(n515) );
  NAND2_X1 U614 ( .A1(n516), .A2(n515), .ZN(n517) );
  INV_X1 U615 ( .A(n523), .ZN(n529) );
  NAND2_X1 U616 ( .A1(n518), .A2(n529), .ZN(n520) );
  NOR2_X1 U617 ( .A1(n520), .A2(n530), .ZN(n521) );
  NAND2_X1 U618 ( .A1(n586), .A2(n521), .ZN(n599) );
  XOR2_X1 U619 ( .A(G101), .B(KEYINPUT111), .Z(n522) );
  XNOR2_X1 U620 ( .A(n599), .B(n522), .ZN(G3) );
  INV_X1 U621 ( .A(KEYINPUT68), .ZN(n524) );
  INV_X1 U622 ( .A(KEYINPUT34), .ZN(n525) );
  NOR2_X1 U623 ( .A1(n569), .A2(n526), .ZN(n565) );
  XNOR2_X1 U624 ( .A(n565), .B(KEYINPUT74), .ZN(n527) );
  XOR2_X1 U625 ( .A(n605), .B(G122), .Z(G24) );
  XNOR2_X1 U626 ( .A(n619), .B(KEYINPUT86), .ZN(n557) );
  NOR2_X1 U627 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U628 ( .A1(n557), .A2(n531), .ZN(n532) );
  XOR2_X1 U629 ( .A(KEYINPUT64), .B(KEYINPUT32), .Z(n534) );
  XNOR2_X1 U630 ( .A(n587), .B(G119), .ZN(G21) );
  INV_X1 U631 ( .A(KEYINPUT42), .ZN(n545) );
  XNOR2_X1 U632 ( .A(n536), .B(KEYINPUT38), .ZN(n631) );
  NAND2_X1 U633 ( .A1(n631), .A2(n630), .ZN(n635) );
  NOR2_X1 U634 ( .A1(n634), .A2(n635), .ZN(n538) );
  XNOR2_X1 U635 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n537) );
  XNOR2_X1 U636 ( .A(n538), .B(n537), .ZN(n649) );
  INV_X1 U637 ( .A(n540), .ZN(n546) );
  XOR2_X1 U638 ( .A(n546), .B(KEYINPUT107), .Z(n541) );
  NAND2_X1 U639 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U640 ( .A(n543), .B(KEYINPUT108), .ZN(n574) );
  NOR2_X1 U641 ( .A1(n649), .A2(n574), .ZN(n544) );
  XNOR2_X1 U642 ( .A(n545), .B(n544), .ZN(n744) );
  INV_X1 U643 ( .A(n593), .ZN(n552) );
  NAND2_X1 U644 ( .A1(n547), .A2(n630), .ZN(n548) );
  XOR2_X1 U645 ( .A(KEYINPUT30), .B(n548), .Z(n551) );
  INV_X1 U646 ( .A(n549), .ZN(n550) );
  XOR2_X1 U647 ( .A(KEYINPUT69), .B(KEYINPUT39), .Z(n553) );
  INV_X1 U648 ( .A(n699), .ZN(n697) );
  NAND2_X1 U649 ( .A1(n581), .A2(n697), .ZN(n555) );
  XOR2_X1 U650 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n554) );
  XNOR2_X1 U651 ( .A(n555), .B(n554), .ZN(n745) );
  NAND2_X1 U652 ( .A1(n744), .A2(n745), .ZN(n556) );
  INV_X1 U653 ( .A(n557), .ZN(n563) );
  INV_X1 U654 ( .A(n558), .ZN(n560) );
  NAND2_X1 U655 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U656 ( .A(n561), .B(KEYINPUT36), .ZN(n562) );
  NOR2_X1 U657 ( .A1(n563), .A2(n562), .ZN(n708) );
  AND2_X1 U658 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U659 ( .A1(n567), .A2(n566), .ZN(n696) );
  NOR2_X1 U660 ( .A1(n569), .A2(n568), .ZN(n693) );
  INV_X1 U661 ( .A(n693), .ZN(n702) );
  NAND2_X1 U662 ( .A1(n699), .A2(n702), .ZN(n596) );
  INV_X1 U663 ( .A(n596), .ZN(n636) );
  NAND2_X1 U664 ( .A1(n636), .A2(KEYINPUT47), .ZN(n570) );
  NAND2_X1 U665 ( .A1(n696), .A2(n570), .ZN(n571) );
  XOR2_X1 U666 ( .A(KEYINPUT75), .B(n571), .Z(n572) );
  NOR2_X1 U667 ( .A1(n708), .A2(n572), .ZN(n578) );
  NAND2_X1 U668 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U669 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U670 ( .A1(n693), .A2(n581), .ZN(n709) );
  NAND2_X1 U671 ( .A1(n618), .A2(n523), .ZN(n584) );
  NOR2_X1 U672 ( .A1(n619), .A2(n584), .ZN(n585) );
  NAND2_X1 U673 ( .A1(n586), .A2(n585), .ZN(n692) );
  NAND2_X1 U674 ( .A1(n587), .A2(n692), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n604), .A2(KEYINPUT44), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n588), .A2(n592), .ZN(n625) );
  NOR2_X1 U677 ( .A1(n625), .A2(n589), .ZN(n591) );
  XNOR2_X1 U678 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n590) );
  XNOR2_X1 U679 ( .A(n591), .B(n590), .ZN(n703) );
  NOR2_X1 U680 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U681 ( .A1(n595), .A2(n594), .ZN(n688) );
  NAND2_X1 U682 ( .A1(n703), .A2(n688), .ZN(n597) );
  NAND2_X1 U683 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U684 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U685 ( .A(n600), .B(KEYINPUT105), .ZN(n601) );
  NOR2_X1 U686 ( .A1(n604), .A2(KEYINPUT44), .ZN(n607) );
  INV_X1 U687 ( .A(n605), .ZN(n606) );
  NAND2_X1 U688 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U689 ( .A(KEYINPUT2), .B(KEYINPUT76), .ZN(n610) );
  OR2_X1 U690 ( .A1(n658), .A2(n610), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n611), .A2(KEYINPUT2), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n614), .A2(n660), .ZN(n653) );
  AND2_X1 U693 ( .A1(n615), .A2(n523), .ZN(n616) );
  XNOR2_X1 U694 ( .A(n616), .B(KEYINPUT49), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n623) );
  NOR2_X1 U696 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n621), .B(KEYINPUT50), .ZN(n622) );
  NOR2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U699 ( .A(n624), .B(KEYINPUT115), .ZN(n626) );
  NAND2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(KEYINPUT51), .ZN(n628) );
  XNOR2_X1 U702 ( .A(KEYINPUT116), .B(n628), .ZN(n629) );
  NOR2_X1 U703 ( .A1(n649), .A2(n629), .ZN(n643) );
  NOR2_X1 U704 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U705 ( .A(KEYINPUT117), .B(n632), .Z(n633) );
  NOR2_X1 U706 ( .A1(n634), .A2(n633), .ZN(n638) );
  NOR2_X1 U707 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U708 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n639), .B(KEYINPUT118), .ZN(n640) );
  NOR2_X1 U710 ( .A1(n648), .A2(n640), .ZN(n641) );
  XOR2_X1 U711 ( .A(KEYINPUT119), .B(n641), .Z(n642) );
  NOR2_X1 U712 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U713 ( .A(KEYINPUT120), .B(n644), .Z(n645) );
  XOR2_X1 U714 ( .A(KEYINPUT52), .B(n645), .Z(n647) );
  NOR2_X1 U715 ( .A1(n647), .A2(n646), .ZN(n651) );
  NOR2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U717 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U718 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U719 ( .A(n654), .B(KEYINPUT121), .ZN(n655) );
  NAND2_X1 U720 ( .A1(n655), .A2(n735), .ZN(n657) );
  XOR2_X1 U721 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n656) );
  XNOR2_X1 U722 ( .A(n657), .B(n656), .ZN(G75) );
  NAND2_X1 U723 ( .A1(n681), .A2(G210), .ZN(n664) );
  XOR2_X1 U724 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n661) );
  XNOR2_X1 U725 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U726 ( .A(n664), .B(n663), .ZN(n666) );
  INV_X1 U727 ( .A(G952), .ZN(n665) );
  XOR2_X1 U728 ( .A(KEYINPUT81), .B(KEYINPUT56), .Z(n667) );
  XNOR2_X1 U729 ( .A(n668), .B(n667), .ZN(G51) );
  NAND2_X1 U730 ( .A1(n681), .A2(G475), .ZN(n673) );
  XNOR2_X1 U731 ( .A(KEYINPUT65), .B(KEYINPUT87), .ZN(n669) );
  XOR2_X1 U732 ( .A(n669), .B(KEYINPUT59), .Z(n670) );
  XNOR2_X1 U733 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U734 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U735 ( .A(n675), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 U736 ( .A(KEYINPUT63), .ZN(n680) );
  NAND2_X1 U737 ( .A1(n681), .A2(G472), .ZN(n678) );
  XNOR2_X1 U738 ( .A(n676), .B(KEYINPUT62), .ZN(n677) );
  XNOR2_X1 U739 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U740 ( .A1(n713), .A2(G469), .ZN(n685) );
  XOR2_X1 U741 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n682) );
  XNOR2_X1 U742 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U743 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X1 U744 ( .A1(n686), .A2(n717), .ZN(G54) );
  NOR2_X1 U745 ( .A1(n688), .A2(n699), .ZN(n687) );
  XOR2_X1 U746 ( .A(G104), .B(n687), .Z(G6) );
  NOR2_X1 U747 ( .A1(n688), .A2(n702), .ZN(n690) );
  XNOR2_X1 U748 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n689) );
  XNOR2_X1 U749 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U750 ( .A(G107), .B(n691), .ZN(G9) );
  XNOR2_X1 U751 ( .A(G110), .B(n692), .ZN(G12) );
  XOR2_X1 U752 ( .A(G128), .B(KEYINPUT29), .Z(n695) );
  XNOR2_X1 U753 ( .A(n695), .B(n694), .ZN(G30) );
  XNOR2_X1 U754 ( .A(G143), .B(n696), .ZN(G45) );
  XNOR2_X1 U755 ( .A(n698), .B(G146), .ZN(G48) );
  NOR2_X1 U756 ( .A1(n703), .A2(n699), .ZN(n700) );
  XOR2_X1 U757 ( .A(KEYINPUT112), .B(n700), .Z(n701) );
  XNOR2_X1 U758 ( .A(G113), .B(n701), .ZN(G15) );
  NOR2_X1 U759 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U760 ( .A(G116), .B(n704), .Z(G18) );
  XOR2_X1 U761 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n706) );
  XNOR2_X1 U762 ( .A(G125), .B(KEYINPUT37), .ZN(n705) );
  XNOR2_X1 U763 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U764 ( .A(n708), .B(n707), .ZN(G27) );
  XNOR2_X1 U765 ( .A(G134), .B(n709), .ZN(G36) );
  NAND2_X1 U766 ( .A1(n713), .A2(G478), .ZN(n711) );
  XNOR2_X1 U767 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U768 ( .A1(n717), .A2(n712), .ZN(G63) );
  NAND2_X1 U769 ( .A1(n713), .A2(G217), .ZN(n715) );
  XNOR2_X1 U770 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U771 ( .A1(n717), .A2(n716), .ZN(G66) );
  INV_X1 U772 ( .A(n718), .ZN(n719) );
  NOR2_X1 U773 ( .A1(n719), .A2(G953), .ZN(n724) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n720) );
  XOR2_X1 U775 ( .A(KEYINPUT61), .B(n720), .Z(n721) );
  NOR2_X1 U776 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U777 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U778 ( .A(n725), .B(KEYINPUT125), .Z(n731) );
  XNOR2_X1 U779 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n727) );
  XOR2_X1 U780 ( .A(n727), .B(n726), .Z(n729) );
  NAND2_X1 U781 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U782 ( .A(n731), .B(n730), .ZN(G69) );
  XOR2_X1 U783 ( .A(n733), .B(n732), .Z(n738) );
  XOR2_X1 U784 ( .A(n738), .B(n734), .Z(n736) );
  NAND2_X1 U785 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U786 ( .A(n737), .B(KEYINPUT126), .ZN(n742) );
  XNOR2_X1 U787 ( .A(G227), .B(n738), .ZN(n739) );
  NAND2_X1 U788 ( .A1(n739), .A2(G900), .ZN(n740) );
  NAND2_X1 U789 ( .A1(n740), .A2(G953), .ZN(n741) );
  NAND2_X1 U790 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U791 ( .A(KEYINPUT127), .B(n743), .Z(G72) );
  XNOR2_X1 U792 ( .A(G137), .B(n744), .ZN(G39) );
  XNOR2_X1 U793 ( .A(n745), .B(G131), .ZN(G33) );
endmodule

