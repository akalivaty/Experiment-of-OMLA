//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n202), .A2(G77), .A3(new_n204), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n214), .B(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n210), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n204), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n216), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G68), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g0026(.A1(new_n226), .A2(G238), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G107), .A2(G264), .ZN(new_n231));
  NAND4_X1  g0031(.A1(new_n228), .A2(new_n229), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n212), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  OR2_X1    g0033(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n221), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT67), .Z(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G226), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XOR2_X1   g0047(.A(G50), .B(G58), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n217), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n210), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n210), .B1(new_n201), .B2(new_n203), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n255), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n255), .ZN(new_n266));
  INV_X1    g0066(.A(G50), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n267), .B1(new_n209), .B2(G20), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n266), .A2(new_n268), .B1(new_n267), .B2(new_n265), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT9), .ZN(new_n271));
  AND2_X1   g0071(.A1(G1), .A2(G13), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G226), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n279), .A2(new_n280), .A3(new_n275), .ZN(new_n281));
  OR3_X1    g0081(.A1(new_n278), .A2(new_n281), .A3(KEYINPUT69), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G222), .A2(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G223), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n287), .B(new_n279), .C1(G77), .C2(new_n283), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT69), .B1(new_n278), .B2(new_n281), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n282), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G200), .ZN(new_n291));
  INV_X1    g0091(.A(G190), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n271), .B(new_n291), .C1(new_n292), .C2(new_n290), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT10), .ZN(new_n294));
  INV_X1    g0094(.A(G169), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n296), .B(new_n270), .C1(G179), .C2(new_n290), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT70), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n280), .B1(new_n272), .B2(new_n273), .ZN(new_n299));
  INV_X1    g0099(.A(new_n275), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G244), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n276), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n283), .A2(G238), .A3(G1698), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n283), .A2(G232), .A3(new_n285), .ZN(new_n305));
  INV_X1    g0105(.A(G107), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n304), .B(new_n305), .C1(new_n306), .C2(new_n283), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n303), .B1(new_n307), .B2(new_n279), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G20), .A2(G77), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n311), .B1(new_n312), .B2(new_n257), .C1(new_n260), .C2(new_n256), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n313), .A2(new_n255), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n209), .A2(G20), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n266), .A2(G77), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(G77), .B2(new_n264), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n310), .B1(G169), .B2(new_n308), .C1(new_n314), .C2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n314), .A2(new_n317), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n308), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT71), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n319), .B(KEYINPUT71), .C1(new_n308), .C2(new_n320), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n308), .A2(G190), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n294), .A2(new_n298), .A3(new_n318), .A4(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G223), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(G1698), .ZN(new_n329));
  INV_X1    g0129(.A(G33), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT3), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G33), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n329), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT76), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT76), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n283), .A2(new_n336), .A3(new_n329), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n331), .A2(new_n333), .A3(G226), .A4(G1698), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G33), .A2(G87), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n274), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G232), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n301), .B1(new_n276), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(G169), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n344), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n339), .A2(new_n340), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n337), .B2(new_n335), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n346), .B(G179), .C1(new_n348), .C2(new_n274), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(G20), .B1(new_n331), .B2(new_n333), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(KEYINPUT7), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT7), .ZN(new_n353));
  AOI211_X1 g0153(.A(new_n353), .B(G20), .C1(new_n331), .C2(new_n333), .ZN(new_n354));
  OAI21_X1  g0154(.A(G68), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT66), .B(G68), .ZN(new_n356));
  INV_X1    g0156(.A(G58), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n204), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(G20), .B1(G159), .B2(new_n259), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n355), .A2(new_n359), .A3(KEYINPUT16), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n255), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT16), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n331), .A2(new_n333), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n210), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n210), .A2(KEYINPUT7), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n332), .A2(G33), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(KEYINPUT74), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT74), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n331), .A2(new_n333), .A3(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n364), .A2(new_n353), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT75), .B1(new_n370), .B2(new_n356), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n366), .A2(KEYINPUT74), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n353), .A2(G20), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n369), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n353), .B1(new_n283), .B2(G20), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n356), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT75), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n371), .A2(new_n378), .A3(new_n359), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n361), .B1(new_n362), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n266), .ZN(new_n381));
  INV_X1    g0181(.A(new_n256), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n315), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n381), .A2(new_n383), .B1(new_n264), .B2(new_n382), .ZN(new_n384));
  OAI211_X1 g0184(.A(KEYINPUT18), .B(new_n350), .C1(new_n380), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT77), .ZN(new_n386));
  INV_X1    g0186(.A(new_n384), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n203), .B1(new_n226), .B2(G58), .ZN(new_n388));
  INV_X1    g0188(.A(G159), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n388), .A2(new_n210), .B1(new_n389), .B2(new_n260), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n331), .A2(new_n333), .A3(new_n368), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n373), .B1(new_n331), .B2(new_n368), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n391), .A2(new_n392), .B1(new_n351), .B2(KEYINPUT7), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n226), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n390), .B1(new_n394), .B2(KEYINPUT75), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT16), .B1(new_n395), .B2(new_n378), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n387), .B1(new_n396), .B2(new_n361), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT77), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT18), .A4(new_n350), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT18), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n359), .B1(new_n376), .B2(new_n377), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n370), .A2(KEYINPUT75), .A3(new_n356), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n362), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n363), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n222), .B1(new_n375), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n390), .A2(new_n405), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(KEYINPUT16), .B1(new_n217), .B2(new_n254), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n384), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n350), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n400), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n386), .A2(new_n399), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n403), .A2(new_n407), .ZN(new_n412));
  OAI21_X1  g0212(.A(G200), .B1(new_n342), .B2(new_n344), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n346), .B(G190), .C1(new_n348), .C2(new_n274), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT78), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n412), .A2(new_n415), .A3(new_n416), .A4(new_n387), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n408), .A2(new_n416), .A3(KEYINPUT17), .A4(new_n415), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n411), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n327), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n226), .A2(new_n210), .ZN(new_n424));
  INV_X1    g0224(.A(G77), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n260), .A2(new_n267), .B1(new_n257), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n255), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n428), .A2(KEYINPUT11), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(KEYINPUT11), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n266), .A2(G68), .A3(new_n315), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n356), .A2(new_n265), .A3(KEYINPUT12), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n264), .A2(G68), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n431), .B(new_n432), .C1(KEYINPUT12), .C2(new_n433), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n429), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT14), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n331), .A2(new_n333), .A3(G226), .A4(new_n285), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n331), .A2(new_n333), .A3(G232), .A4(G1698), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G97), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT72), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT72), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n437), .A2(new_n438), .A3(new_n442), .A4(new_n439), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n279), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT13), .ZN(new_n445));
  INV_X1    g0245(.A(new_n276), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n281), .B1(G238), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n444), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n445), .B1(new_n444), .B2(new_n447), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n436), .B(G169), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n444), .A2(new_n447), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT13), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n453), .A2(G179), .A3(new_n448), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n448), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n436), .B1(new_n456), .B2(G169), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT73), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(G169), .B1(new_n449), .B2(new_n450), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT14), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT73), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(new_n454), .A4(new_n451), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n435), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n456), .A2(G200), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n453), .A2(G190), .A3(new_n448), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n435), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n423), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n210), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n471), .B1(new_n330), .B2(G97), .ZN(new_n472));
  INV_X1    g0272(.A(G116), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n255), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT86), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n255), .A2(KEYINPUT86), .A3(new_n474), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n472), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT87), .B1(new_n479), .B2(KEYINPUT20), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT87), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT20), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n255), .A2(KEYINPUT86), .A3(new_n474), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT86), .B1(new_n255), .B2(new_n474), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n481), .B(new_n482), .C1(new_n485), .C2(new_n472), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n479), .A2(KEYINPUT20), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n480), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n264), .A2(new_n473), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n266), .B1(G1), .B2(new_n330), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n491), .B2(new_n473), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT5), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT81), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(G41), .ZN(new_n496));
  INV_X1    g0296(.A(G41), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n498));
  INV_X1    g0298(.A(G45), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(G1), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n496), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(G270), .A3(new_n274), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n299), .A2(new_n498), .A3(new_n496), .A4(new_n500), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT84), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT84), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n283), .A2(G257), .A3(new_n285), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n283), .A2(G264), .A3(G1698), .ZN(new_n509));
  INV_X1    g0309(.A(G303), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(new_n283), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n505), .A2(new_n507), .B1(new_n279), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n493), .A2(G179), .A3(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n488), .A2(new_n492), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n279), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n506), .B1(new_n502), .B2(new_n503), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT85), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT85), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n515), .B(new_n520), .C1(new_n516), .C2(new_n517), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(G200), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n505), .A2(new_n507), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n520), .B1(new_n523), .B2(new_n515), .ZN(new_n524));
  INV_X1    g0324(.A(new_n521), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n514), .B(new_n522), .C1(new_n526), .C2(new_n292), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n493), .A2(G169), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n519), .A2(new_n521), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n528), .A2(KEYINPUT21), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT21), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n295), .B1(new_n488), .B2(new_n492), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n513), .B(new_n527), .C1(new_n530), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n501), .A2(G257), .A3(new_n274), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n503), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n331), .A2(new_n333), .A3(G250), .A4(G1698), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n331), .A2(new_n333), .A3(G244), .A4(new_n285), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT4), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n470), .B(new_n538), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT79), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n539), .A2(KEYINPUT79), .A3(new_n540), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(G190), .B(new_n537), .C1(new_n546), .C2(new_n274), .ZN(new_n547));
  INV_X1    g0347(.A(G97), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n265), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n490), .B2(new_n548), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT6), .ZN(new_n551));
  AND2_X1   g0351(.A1(G97), .A2(G107), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(new_n552), .B2(new_n206), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n306), .A2(KEYINPUT6), .A3(G97), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n370), .B2(new_n306), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n550), .B1(new_n557), .B2(new_n255), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT80), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n546), .B2(new_n274), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n539), .A2(new_n540), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n538), .A2(new_n470), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n539), .A2(KEYINPUT79), .A3(new_n540), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT79), .B1(new_n539), .B2(new_n540), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(KEYINPUT80), .A3(new_n279), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n536), .B1(new_n560), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n547), .B(new_n558), .C1(new_n567), .C2(new_n320), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n546), .A2(new_n559), .A3(new_n274), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT80), .B1(new_n565), .B2(new_n279), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n309), .B(new_n537), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n537), .B1(new_n546), .B2(new_n274), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n558), .B1(new_n295), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n491), .A2(G87), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n283), .A2(new_n210), .A3(G68), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n210), .B1(new_n439), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(G87), .B2(new_n207), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n578), .B1(new_n257), .B2(new_n548), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n577), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n582), .A2(new_n255), .B1(new_n265), .B2(new_n312), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n285), .A2(G238), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT83), .B1(new_n363), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT83), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n283), .A2(new_n587), .A3(G238), .A4(new_n285), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n331), .A2(new_n333), .A3(G244), .A4(G1698), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G33), .A2(G116), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n274), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G250), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n279), .A2(new_n595), .A3(new_n500), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT82), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n299), .A2(new_n598), .A3(new_n500), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n598), .B1(new_n299), .B2(new_n500), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(G200), .B1(new_n594), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n299), .A2(new_n500), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT82), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n596), .B1(new_n605), .B2(new_n599), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n592), .B1(new_n588), .B2(new_n586), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(G190), .C1(new_n607), .C2(new_n274), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n584), .A2(new_n603), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n295), .B1(new_n594), .B2(new_n602), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n583), .B1(new_n490), .B2(new_n312), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n606), .B(new_n309), .C1(new_n607), .C2(new_n274), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n501), .A2(new_n274), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n331), .A2(new_n333), .A3(G257), .A4(G1698), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n331), .A2(new_n333), .A3(G250), .A4(new_n285), .ZN(new_n617));
  NAND2_X1  g0417(.A1(G33), .A2(G294), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AOI22_X1  g0419(.A1(G264), .A2(new_n615), .B1(new_n619), .B2(new_n279), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n620), .A2(KEYINPUT88), .A3(new_n292), .A4(new_n503), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT88), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n619), .A2(new_n279), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n501), .A2(G264), .A3(new_n274), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n503), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n622), .B1(new_n625), .B2(new_n320), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(G190), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n621), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n491), .A2(G107), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n264), .A2(G107), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n630), .B(KEYINPUT25), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n331), .A2(new_n333), .A3(new_n210), .A4(G87), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT22), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT22), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n283), .A2(new_n635), .A3(new_n210), .A4(G87), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n591), .A2(G20), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT23), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n210), .B2(G107), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n306), .A2(KEYINPUT23), .A3(G20), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT24), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT24), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n637), .A2(new_n645), .A3(new_n642), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n632), .B1(new_n647), .B2(new_n255), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n628), .A2(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n637), .A2(new_n645), .A3(new_n642), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n645), .B1(new_n637), .B2(new_n642), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n255), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n629), .A3(new_n631), .ZN(new_n653));
  INV_X1    g0453(.A(new_n503), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n620), .A2(G179), .ZN(new_n655));
  INV_X1    g0455(.A(new_n625), .ZN(new_n656));
  OAI22_X1  g0456(.A1(new_n654), .A2(new_n655), .B1(new_n656), .B2(new_n295), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT89), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n649), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n659), .B1(new_n649), .B2(new_n658), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n575), .B(new_n614), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n469), .A2(new_n534), .A3(new_n663), .ZN(G372));
  INV_X1    g0464(.A(new_n298), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n467), .A2(new_n318), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n421), .B1(new_n463), .B2(new_n666), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n408), .A2(new_n400), .A3(new_n409), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT18), .B1(new_n397), .B2(new_n350), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n665), .B1(new_n670), .B2(new_n294), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n568), .A2(new_n574), .A3(new_n614), .A4(new_n649), .ZN(new_n672));
  INV_X1    g0472(.A(new_n513), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT21), .B1(new_n528), .B2(new_n529), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n526), .A2(new_n531), .A3(new_n532), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n672), .B1(new_n676), .B2(new_n658), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n571), .A2(new_n573), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT26), .B1(new_n678), .B2(new_n614), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n609), .A2(new_n613), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n574), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n613), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n671), .B1(new_n469), .B2(new_n684), .ZN(G369));
  INV_X1    g0485(.A(G330), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n513), .B1(new_n530), .B2(new_n533), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT90), .Z(new_n690));
  INV_X1    g0490(.A(G213), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n688), .B2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n493), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT91), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n687), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT92), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT93), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n697), .B1(new_n534), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n700), .B2(new_n534), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n686), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n649), .A2(new_n658), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT89), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n660), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n653), .A2(new_n695), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT94), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT94), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n706), .A2(new_n710), .A3(new_n707), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n695), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n658), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n703), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n658), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n713), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n676), .A2(new_n695), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n709), .A2(new_n711), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n717), .A2(new_n719), .A3(new_n721), .ZN(G399));
  INV_X1    g0522(.A(new_n213), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(G87), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n206), .A2(new_n726), .A3(new_n473), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT95), .Z(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n725), .A2(G1), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n219), .B2(new_n725), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n713), .B1(new_n677), .B2(new_n683), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n736), .B(new_n713), .C1(new_n677), .C2(new_n683), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n568), .A2(new_n574), .A3(new_n614), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n739), .B1(new_n705), .B2(new_n660), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n740), .A2(new_n676), .A3(new_n527), .A4(new_n713), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n620), .A2(G179), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n536), .B1(new_n565), .B2(new_n279), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n594), .A2(new_n602), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n742), .A2(new_n743), .A3(new_n512), .A4(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n655), .A2(new_n594), .A3(new_n602), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n748), .A2(KEYINPUT30), .A3(new_n512), .A4(new_n743), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n625), .B(new_n309), .C1(new_n594), .C2(new_n602), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n529), .A2(new_n567), .A3(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(KEYINPUT31), .B(new_n695), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n537), .B1(new_n569), .B2(new_n570), .ZN(new_n755));
  INV_X1    g0555(.A(new_n751), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n526), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(new_n747), .A3(new_n749), .ZN(new_n758));
  AOI21_X1  g0558(.A(KEYINPUT31), .B1(new_n758), .B2(new_n695), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n686), .B1(new_n741), .B2(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n735), .A2(new_n738), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n732), .B1(new_n762), .B2(G1), .ZN(G364));
  AND2_X1   g0563(.A1(new_n210), .A2(G13), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n209), .B1(new_n764), .B2(G45), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n724), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n703), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n699), .A2(new_n686), .A3(new_n702), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT96), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n768), .A2(KEYINPUT96), .A3(new_n769), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n699), .A2(new_n702), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n767), .ZN(new_n779));
  AND3_X1   g0579(.A1(new_n213), .A2(G355), .A3(new_n283), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n723), .A2(new_n283), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(G45), .B2(new_n219), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(G45), .B2(new_n249), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n780), .B(new_n783), .C1(new_n473), .C2(new_n723), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n217), .B1(G20), .B2(new_n295), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n777), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n779), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n786), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n210), .A2(new_n292), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n309), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n210), .A2(G190), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G58), .A2(new_n793), .B1(new_n796), .B2(G77), .ZN(new_n797));
  NAND3_X1  g0597(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n292), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n797), .B1(new_n267), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT97), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n320), .A2(G179), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n794), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n306), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n790), .A2(new_n803), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n283), .B1(new_n806), .B2(new_n726), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G179), .A2(G200), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n794), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G159), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT32), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n210), .B1(new_n808), .B2(G190), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n798), .A2(G190), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n814), .A2(G97), .B1(G68), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n811), .A2(KEYINPUT32), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n812), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NOR4_X1   g0618(.A1(new_n802), .A2(new_n805), .A3(new_n807), .A4(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G311), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n795), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G322), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n792), .A2(new_n822), .B1(new_n804), .B2(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n821), .B(new_n824), .C1(G329), .C2(new_n810), .ZN(new_n825));
  INV_X1    g0625(.A(G294), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n363), .B1(new_n813), .B2(new_n826), .C1(new_n510), .C2(new_n806), .ZN(new_n827));
  INV_X1    g0627(.A(new_n815), .ZN(new_n828));
  XOR2_X1   g0628(.A(KEYINPUT33), .B(G317), .Z(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n827), .B(new_n830), .C1(G326), .C2(new_n799), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n819), .B1(new_n825), .B2(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n778), .B(new_n788), .C1(new_n789), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n774), .A2(new_n833), .ZN(G396));
  NOR2_X1   g0634(.A1(new_n318), .A2(new_n695), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n326), .B1(new_n319), .B2(new_n713), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(new_n318), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n733), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n713), .B(new_n837), .C1(new_n677), .C2(new_n683), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n761), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n767), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n842), .B2(new_n841), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n789), .A2(new_n776), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n767), .B1(G77), .B2(new_n845), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT98), .Z(new_n847));
  OAI221_X1 g0647(.A(new_n363), .B1(new_n813), .B2(new_n548), .C1(new_n306), .C2(new_n806), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n828), .A2(new_n823), .B1(new_n800), .B2(new_n510), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n792), .A2(new_n826), .B1(new_n804), .B2(new_n726), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n795), .A2(new_n473), .B1(new_n809), .B2(new_n820), .ZN(new_n851));
  NOR4_X1   g0651(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G143), .A2(new_n793), .B1(new_n796), .B2(G159), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n853), .B1(new_n800), .B2(new_n854), .C1(new_n258), .C2(new_n828), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT34), .ZN(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n283), .B1(new_n809), .B2(new_n857), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n806), .A2(new_n267), .B1(new_n804), .B2(new_n222), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n858), .B(new_n859), .C1(G58), .C2(new_n814), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n852), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n847), .B1(new_n789), .B2(new_n861), .C1(new_n837), .C2(new_n776), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n844), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G384));
  NOR2_X1   g0664(.A1(new_n764), .A2(new_n209), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n408), .A2(new_n415), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n406), .A2(KEYINPUT16), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n387), .B1(new_n867), .B2(new_n361), .ZN(new_n868));
  INV_X1    g0668(.A(new_n693), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n868), .B1(new_n350), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT37), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n397), .A2(new_n350), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n869), .B1(new_n380), .B2(new_n384), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n873), .A2(new_n874), .A3(new_n866), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n419), .A2(new_n420), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n669), .B1(KEYINPUT77), .B2(new_n385), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n878), .B1(new_n879), .B2(new_n399), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n868), .A2(new_n869), .ZN(new_n881));
  OAI211_X1 g0681(.A(KEYINPUT38), .B(new_n877), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n874), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n669), .A2(new_n668), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n883), .B1(new_n884), .B2(new_n878), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n873), .A2(new_n874), .A3(new_n866), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n876), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n882), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT40), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n838), .B1(new_n741), .B2(new_n760), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n458), .A2(new_n462), .ZN(new_n895));
  INV_X1    g0695(.A(new_n435), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n435), .A2(new_n713), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n897), .A2(new_n466), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n898), .B1(new_n463), .B2(new_n467), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n894), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n893), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n881), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n422), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n906), .B2(new_n877), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n881), .B1(new_n411), .B2(new_n421), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n872), .A2(new_n876), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n908), .A2(new_n890), .A3(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n902), .B(new_n894), .C1(new_n907), .C2(new_n910), .ZN(new_n911));
  XOR2_X1   g0711(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT102), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n911), .A2(KEYINPUT102), .A3(new_n912), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n904), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT103), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n469), .B1(new_n741), .B2(new_n760), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n686), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n918), .B2(new_n919), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n890), .B1(new_n908), .B2(new_n909), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n882), .A2(new_n922), .A3(KEYINPUT39), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT39), .B1(new_n882), .B2(new_n891), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n897), .A2(new_n695), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n835), .B(KEYINPUT100), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n840), .A2(new_n928), .B1(new_n900), .B2(new_n901), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n882), .A2(new_n922), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n929), .A2(new_n930), .B1(new_n884), .B2(new_n693), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n671), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n469), .B1(new_n734), .B2(new_n737), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n932), .B(new_n935), .Z(new_n936));
  AOI21_X1  g0736(.A(new_n865), .B1(new_n921), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n936), .B2(new_n921), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n555), .A2(KEYINPUT35), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n555), .A2(KEYINPUT35), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n939), .A2(G116), .A3(new_n218), .A4(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(KEYINPUT99), .B(KEYINPUT36), .Z(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n220), .B(G77), .C1(new_n357), .C2(new_n356), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n201), .A2(G68), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n209), .B(G13), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n938), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT104), .Z(G367));
  OAI21_X1  g0749(.A(new_n575), .B1(new_n558), .B2(new_n713), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n678), .A2(new_n695), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n717), .A2(KEYINPUT105), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(KEYINPUT105), .B1(new_n717), .B2(new_n953), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n713), .A2(new_n584), .ZN(new_n957));
  INV_X1    g0757(.A(new_n613), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n681), .B2(new_n957), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n956), .B1(KEYINPUT43), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n718), .A2(new_n568), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n695), .B1(new_n963), .B2(new_n574), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n721), .A2(new_n953), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n964), .B1(new_n965), .B2(KEYINPUT42), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(KEYINPUT42), .B2(new_n965), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n954), .A2(new_n968), .A3(new_n955), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n961), .A2(new_n962), .A3(new_n967), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n961), .A2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n967), .A2(new_n962), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n724), .B(KEYINPUT41), .Z(new_n974));
  NAND3_X1  g0774(.A1(new_n721), .A2(new_n719), .A3(new_n952), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT45), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n721), .A2(new_n719), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n953), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT44), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n980), .A2(KEYINPUT44), .A3(new_n953), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n979), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n986), .A2(KEYINPUT106), .A3(new_n703), .A4(new_n716), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n977), .A2(new_n978), .B1(new_n983), .B2(new_n984), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT106), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n717), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n762), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n716), .A2(new_n720), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n721), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n703), .ZN(new_n994));
  INV_X1    g0794(.A(new_n703), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n992), .A2(new_n995), .A3(new_n721), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n991), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n987), .A2(new_n990), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n974), .B1(new_n998), .B2(new_n762), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n970), .B(new_n973), .C1(new_n999), .C2(new_n766), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n787), .B1(new_n213), .B2(new_n312), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n781), .B2(new_n245), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n800), .A2(new_n820), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n283), .B(new_n1003), .C1(G317), .C2(new_n810), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n806), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(G116), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT46), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n814), .A2(G107), .B1(G294), .B2(new_n815), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n792), .A2(new_n510), .B1(new_n795), .B2(new_n823), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n804), .A2(new_n548), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1004), .A2(new_n1007), .A3(new_n1008), .A4(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n813), .A2(new_n222), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G150), .B2(new_n793), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT107), .Z(new_n1015));
  OAI21_X1  g0815(.A(new_n283), .B1(new_n795), .B2(new_n201), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G143), .B2(new_n799), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n804), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(G77), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G58), .A2(new_n1005), .B1(new_n810), .B2(G137), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n815), .A2(G159), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1012), .B1(new_n1015), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT47), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n779), .B(new_n1002), .C1(new_n1024), .C2(new_n786), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n777), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1025), .B1(new_n960), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1000), .A2(new_n1027), .ZN(G387));
  NAND2_X1  g0828(.A1(new_n994), .A2(new_n996), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n762), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n994), .A2(new_n991), .A3(new_n996), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n724), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n712), .A2(new_n715), .A3(new_n777), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n806), .A2(new_n826), .B1(new_n813), .B2(new_n823), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G317), .A2(new_n793), .B1(new_n796), .B2(G303), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n800), .B2(new_n822), .C1(new_n820), .C2(new_n828), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT48), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n1037), .B2(new_n1036), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT49), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n804), .A2(new_n473), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n283), .B(new_n1043), .C1(G326), .C2(new_n810), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n806), .A2(new_n425), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n792), .A2(new_n267), .B1(new_n795), .B2(new_n222), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(G150), .C2(new_n810), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n363), .B(new_n1010), .C1(new_n382), .C2(new_n815), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n813), .A2(new_n312), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n799), .A2(G159), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n789), .B1(new_n1045), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n728), .A2(new_n213), .A3(new_n283), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n729), .B(new_n499), .C1(new_n222), .C2(new_n425), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT108), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n382), .A2(new_n267), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT50), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n242), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n781), .B1(new_n1060), .B2(new_n499), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1054), .B1(G107), .B2(new_n213), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n779), .B(new_n1053), .C1(new_n787), .C2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1029), .A2(new_n766), .B1(new_n1033), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1032), .A2(new_n1064), .ZN(G393));
  INV_X1    g0865(.A(new_n781), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n787), .B1(new_n548), .B2(new_n213), .C1(new_n1066), .C2(new_n252), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1067), .A2(new_n767), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n813), .A2(new_n425), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n256), .B2(new_n795), .C1(new_n828), .C2(new_n201), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT109), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n800), .A2(new_n258), .B1(new_n792), .B2(new_n389), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n363), .B1(new_n1018), .B2(G87), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n226), .A2(new_n1005), .B1(new_n810), .B2(G143), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n793), .A2(G311), .B1(G317), .B2(new_n799), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT52), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n806), .A2(new_n823), .B1(new_n809), .B2(new_n822), .ZN(new_n1080));
  NOR4_X1   g0880(.A1(new_n1079), .A2(new_n283), .A3(new_n805), .A4(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n795), .A2(new_n826), .B1(new_n813), .B2(new_n473), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G303), .B2(new_n815), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT110), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1072), .A2(new_n1077), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1068), .B1(new_n789), .B2(new_n1085), .C1(new_n952), .C2(new_n1026), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n988), .B(new_n717), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1086), .B1(new_n1087), .B2(new_n765), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n725), .B1(new_n1087), .B2(new_n1030), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1088), .B1(new_n998), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(G390));
  INV_X1    g0891(.A(KEYINPUT114), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n894), .A2(new_n902), .A3(G330), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n926), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n840), .A2(new_n928), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n902), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT39), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT38), .B1(new_n885), .B2(new_n888), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1098), .B1(new_n910), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n882), .A2(new_n922), .A3(KEYINPUT39), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1095), .A2(new_n1097), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n910), .A2(new_n1099), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n929), .A2(new_n1103), .A3(new_n926), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1094), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n923), .A2(new_n924), .B1(new_n929), .B2(new_n926), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1097), .A2(new_n1095), .A3(new_n892), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n1093), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1092), .B1(new_n1109), .B2(new_n765), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1105), .A2(KEYINPUT114), .A3(new_n766), .A4(new_n1108), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n767), .B1(new_n382), .B2(new_n845), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n804), .A2(new_n222), .B1(new_n809), .B2(new_n826), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT116), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1070), .B1(new_n800), .B2(new_n823), .C1(new_n306), .C2(new_n828), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n363), .B1(new_n806), .B2(new_n726), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n792), .A2(new_n473), .B1(new_n795), .B2(new_n548), .ZN(new_n1118));
  OR4_X1    g0918(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(G128), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n828), .A2(new_n854), .B1(new_n800), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G159), .B2(new_n814), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1005), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT53), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n806), .B2(new_n258), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n283), .B1(new_n804), .B2(new_n201), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1123), .A2(new_n1125), .B1(KEYINPUT115), .B2(new_n1126), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n1126), .A2(KEYINPUT115), .ZN(new_n1128));
  INV_X1    g0928(.A(G125), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n792), .A2(new_n857), .B1(new_n809), .B2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1130), .B1(new_n796), .B2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1122), .A2(new_n1127), .A3(new_n1128), .A4(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1119), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1113), .B1(new_n1135), .B2(new_n786), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n925), .B2(new_n776), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1112), .A2(new_n1137), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1106), .A2(new_n1093), .A3(new_n1107), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1093), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(KEYINPUT111), .B1(new_n842), .B2(new_n469), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n469), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT111), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1143), .A2(new_n1144), .A3(new_n761), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n663), .A2(new_n534), .A3(new_n695), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n758), .A2(new_n695), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT31), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n753), .ZN(new_n1151));
  OAI211_X1 g0951(.A(G330), .B(new_n837), .C1(new_n1147), .C2(new_n1151), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n900), .A2(new_n901), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1096), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1154), .A2(new_n1155), .A3(new_n1093), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1154), .B2(new_n1093), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n935), .B(new_n1146), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT112), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1141), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(KEYINPUT112), .B1(new_n1109), .B2(new_n1158), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1109), .A2(KEYINPUT113), .A3(new_n1158), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n724), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT113), .B1(new_n1109), .B2(new_n1158), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1138), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(G378));
  NAND2_X1  g0969(.A1(new_n294), .A2(new_n297), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n869), .A2(new_n270), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1170), .B(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1172), .B(new_n1173), .Z(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n917), .A2(G330), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n904), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n911), .A2(KEYINPUT102), .A3(new_n912), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT102), .B1(new_n911), .B2(new_n912), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1177), .B(G330), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n1174), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n932), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1176), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1182), .B1(new_n1176), .B2(new_n1181), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n766), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1174), .A2(new_n775), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n767), .B1(new_n202), .B2(new_n845), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n283), .A2(G41), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1190), .A2(new_n1046), .A3(new_n1013), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n548), .B2(new_n828), .C1(new_n473), .C2(new_n800), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n792), .A2(new_n306), .B1(new_n809), .B2(new_n823), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n312), .A2(new_n795), .B1(new_n804), .B2(new_n357), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1190), .B(new_n267), .C1(G33), .C2(G41), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n806), .A2(new_n1131), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n792), .A2(new_n1120), .B1(new_n795), .B2(new_n854), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(G132), .C2(new_n815), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n800), .A2(new_n1129), .B1(new_n813), .B2(new_n258), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT118), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1018), .A2(G159), .ZN(new_n1209));
  AOI211_X1 g1009(.A(G33), .B(G41), .C1(new_n810), .C2(G124), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1200), .B1(new_n1207), .B2(new_n1211), .C1(new_n1197), .C2(new_n1195), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1188), .B1(new_n1212), .B2(new_n786), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1187), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1186), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1175), .B1(new_n917), .B2(G330), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1180), .A2(new_n1174), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n932), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n1183), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n934), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n842), .A2(new_n469), .A3(KEYINPUT111), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1144), .B1(new_n1143), .B2(new_n761), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n671), .B(new_n1220), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1160), .B1(new_n1141), .B2(new_n1159), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1109), .A2(KEYINPUT112), .A3(new_n1158), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1219), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT57), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n725), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT119), .B1(new_n1218), .B2(new_n1183), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1183), .A2(KEYINPUT119), .ZN(new_n1232));
  OAI211_X1 g1032(.A(KEYINPUT57), .B(new_n1227), .C1(new_n1231), .C2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1215), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(G375));
  INV_X1    g1035(.A(new_n1157), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1154), .A2(new_n1155), .A3(new_n1093), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1153), .A2(new_n775), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n767), .B1(G68), .B2(new_n845), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n806), .A2(new_n548), .B1(new_n809), .B2(new_n510), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT120), .Z(new_n1242));
  OAI221_X1 g1042(.A(new_n1050), .B1(new_n800), .B2(new_n826), .C1(new_n473), .C2(new_n828), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1019), .A2(new_n363), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n792), .A2(new_n823), .B1(new_n795), .B2(new_n306), .ZN(new_n1245));
  OR3_X1    g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n795), .A2(new_n258), .B1(new_n809), .B2(new_n1120), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n283), .B1(new_n804), .B2(new_n357), .C1(new_n828), .C2(new_n1131), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n854), .A2(new_n792), .B1(new_n806), .B2(new_n389), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n813), .A2(new_n267), .ZN(new_n1250));
  OR4_X1    g1050(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n799), .A2(G132), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT121), .Z(new_n1253));
  OAI22_X1  g1053(.A1(new_n1242), .A2(new_n1246), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1240), .B1(new_n1254), .B2(new_n786), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1238), .A2(new_n766), .B1(new_n1239), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n974), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1158), .A2(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1224), .A2(new_n1238), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1256), .B1(new_n1258), .B2(new_n1259), .ZN(G381));
  NAND3_X1  g1060(.A1(new_n1000), .A2(new_n1090), .A3(new_n1027), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(G396), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1032), .A2(new_n1263), .A3(new_n1064), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1264), .A2(G384), .A3(G381), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1234), .A2(new_n1168), .A3(new_n1262), .A4(new_n1265), .ZN(G407));
  NOR2_X1   g1066(.A1(new_n691), .A2(G343), .ZN(new_n1267));
  XOR2_X1   g1067(.A(new_n1267), .B(KEYINPUT122), .Z(new_n1268));
  NAND3_X1  g1068(.A1(new_n1234), .A2(new_n1168), .A3(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(G407), .A2(G213), .A3(new_n1269), .ZN(G409));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1090), .B1(new_n1000), .B2(new_n1027), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1264), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1263), .B1(new_n1032), .B2(new_n1064), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT123), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G393), .A2(G396), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT123), .B1(new_n1277), .B2(new_n1264), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1262), .A2(new_n1272), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G387), .A2(G390), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1276), .B1(new_n1281), .B2(new_n1261), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1271), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1267), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1168), .B(new_n1215), .C1(new_n1230), .C2(new_n1233), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1214), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1219), .A2(new_n1227), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(new_n1287), .B2(new_n1257), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n766), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G378), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1284), .B1(new_n1285), .B2(new_n1290), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1158), .A2(KEYINPUT60), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n725), .B1(new_n1292), .B2(new_n1259), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(new_n1259), .B2(new_n1292), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1256), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n863), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(G384), .A3(new_n1256), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(G2897), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1284), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n1296), .A2(new_n1297), .B1(G2897), .B2(new_n1268), .ZN(new_n1301));
  OR2_X1    g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1283), .B1(new_n1291), .B2(new_n1302), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1284), .B(new_n1304), .C1(new_n1285), .C2(new_n1290), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT63), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1168), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1234), .A2(G378), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1268), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT124), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1298), .A2(new_n1306), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1312), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1303), .B(new_n1307), .C1(new_n1314), .C2(new_n1315), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1317), .B1(new_n1311), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1298), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1268), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1321), .B(new_n1322), .C1(new_n1285), .C2(new_n1290), .ZN(new_n1323));
  AOI22_X1  g1123(.A1(KEYINPUT126), .A2(new_n1323), .B1(new_n1305), .B2(new_n1320), .ZN(new_n1324));
  OR2_X1    g1124(.A1(new_n1323), .A2(KEYINPUT126), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1319), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1281), .B(new_n1261), .C1(new_n1276), .C2(new_n1278), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT127), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1262), .A2(new_n1272), .ZN(new_n1329));
  OAI211_X1 g1129(.A(new_n1327), .B(new_n1328), .C1(new_n1329), .C2(new_n1276), .ZN(new_n1330));
  OAI21_X1  g1130(.A(KEYINPUT127), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1316), .B1(new_n1326), .B2(new_n1332), .ZN(G405));
  NOR2_X1   g1133(.A1(new_n1234), .A2(G378), .ZN(new_n1334));
  OR3_X1    g1134(.A1(new_n1334), .A2(new_n1285), .A3(new_n1304), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1304), .B1(new_n1334), .B2(new_n1285), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  XOR2_X1   g1137(.A(new_n1337), .B(new_n1332), .Z(G402));
endmodule


