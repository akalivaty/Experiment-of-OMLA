

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575;

  NOR2_X1 U318 ( .A1(n441), .A2(n520), .ZN(n557) );
  AND2_X1 U319 ( .A1(G230GAT), .A2(G233GAT), .ZN(n286) );
  XNOR2_X1 U320 ( .A(n365), .B(n286), .ZN(n322) );
  XOR2_X1 U321 ( .A(G57GAT), .B(KEYINPUT13), .Z(n342) );
  XNOR2_X1 U322 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U323 ( .A(n328), .B(n414), .ZN(n329) );
  XNOR2_X1 U324 ( .A(n330), .B(n329), .ZN(n332) );
  INV_X1 U325 ( .A(KEYINPUT123), .ZN(n442) );
  XOR2_X1 U326 ( .A(n440), .B(n439), .Z(n520) );
  XNOR2_X1 U327 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U328 ( .A(n445), .B(n444), .ZN(G1348GAT) );
  XOR2_X1 U329 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n288) );
  NAND2_X1 U330 ( .A1(G229GAT), .A2(G233GAT), .ZN(n287) );
  XNOR2_X1 U331 ( .A(n288), .B(n287), .ZN(n289) );
  XOR2_X1 U332 ( .A(n289), .B(KEYINPUT68), .Z(n297) );
  XOR2_X1 U333 ( .A(G113GAT), .B(G50GAT), .Z(n291) );
  XNOR2_X1 U334 ( .A(G169GAT), .B(G43GAT), .ZN(n290) );
  XNOR2_X1 U335 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U336 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n293) );
  XNOR2_X1 U337 ( .A(G197GAT), .B(G141GAT), .ZN(n292) );
  XNOR2_X1 U338 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n303) );
  XOR2_X1 U341 ( .A(G29GAT), .B(G36GAT), .Z(n299) );
  XNOR2_X1 U342 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n299), .B(n298), .ZN(n361) );
  XOR2_X1 U344 ( .A(G1GAT), .B(G8GAT), .Z(n301) );
  XNOR2_X1 U345 ( .A(G15GAT), .B(G22GAT), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n343) );
  XOR2_X1 U347 ( .A(n361), .B(n343), .Z(n302) );
  XOR2_X1 U348 ( .A(n303), .B(n302), .Z(n523) );
  INV_X1 U349 ( .A(n523), .ZN(n563) );
  XOR2_X1 U350 ( .A(G92GAT), .B(G8GAT), .Z(n305) );
  NAND2_X1 U351 ( .A1(G226GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n307) );
  XNOR2_X1 U353 ( .A(G176GAT), .B(G204GAT), .ZN(n306) );
  XOR2_X1 U354 ( .A(n306), .B(G64GAT), .Z(n331) );
  XNOR2_X1 U355 ( .A(n307), .B(n331), .ZN(n313) );
  XNOR2_X1 U356 ( .A(G211GAT), .B(KEYINPUT87), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n308), .B(KEYINPUT21), .ZN(n309) );
  XOR2_X1 U358 ( .A(n309), .B(KEYINPUT88), .Z(n311) );
  XNOR2_X1 U359 ( .A(G197GAT), .B(G218GAT), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n423) );
  XNOR2_X1 U361 ( .A(G36GAT), .B(n423), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n320) );
  XOR2_X1 U363 ( .A(G183GAT), .B(KEYINPUT81), .Z(n315) );
  XNOR2_X1 U364 ( .A(G169GAT), .B(KEYINPUT80), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U366 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n317) );
  XNOR2_X1 U367 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U369 ( .A(n319), .B(n318), .ZN(n440) );
  XNOR2_X1 U370 ( .A(n320), .B(n440), .ZN(n510) );
  XOR2_X1 U371 ( .A(KEYINPUT46), .B(KEYINPUT116), .Z(n339) );
  XNOR2_X1 U372 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n333) );
  XNOR2_X1 U373 ( .A(n342), .B(KEYINPUT32), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n321), .B(KEYINPUT31), .ZN(n323) );
  XOR2_X1 U375 ( .A(G85GAT), .B(G92GAT), .Z(n365) );
  XOR2_X1 U376 ( .A(n324), .B(KEYINPUT33), .Z(n330) );
  XNOR2_X1 U377 ( .A(G99GAT), .B(G71GAT), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n325), .B(G120GAT), .ZN(n436) );
  XNOR2_X1 U379 ( .A(n436), .B(KEYINPUT71), .ZN(n328) );
  XOR2_X1 U380 ( .A(G78GAT), .B(G148GAT), .Z(n327) );
  XNOR2_X1 U381 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n414) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n334) );
  NAND2_X1 U384 ( .A1(n333), .A2(n334), .ZN(n337) );
  INV_X1 U385 ( .A(n333), .ZN(n335) );
  INV_X1 U386 ( .A(n334), .ZN(n377) );
  NAND2_X1 U387 ( .A1(n335), .A2(n377), .ZN(n336) );
  NAND2_X1 U388 ( .A1(n337), .A2(n336), .ZN(n541) );
  NAND2_X1 U389 ( .A1(n541), .A2(n563), .ZN(n338) );
  XNOR2_X1 U390 ( .A(n339), .B(n338), .ZN(n357) );
  XOR2_X1 U391 ( .A(G78GAT), .B(G155GAT), .Z(n341) );
  XNOR2_X1 U392 ( .A(G127GAT), .B(G211GAT), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n356) );
  XOR2_X1 U394 ( .A(n342), .B(G71GAT), .Z(n345) );
  XNOR2_X1 U395 ( .A(n343), .B(G183GAT), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U397 ( .A(KEYINPUT15), .B(KEYINPUT75), .Z(n347) );
  NAND2_X1 U398 ( .A1(G231GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U400 ( .A(n349), .B(n348), .Z(n354) );
  XOR2_X1 U401 ( .A(KEYINPUT14), .B(KEYINPUT74), .Z(n351) );
  XNOR2_X1 U402 ( .A(G64GAT), .B(KEYINPUT73), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U404 ( .A(n352), .B(KEYINPUT12), .ZN(n353) );
  XNOR2_X1 U405 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U406 ( .A(n356), .B(n355), .Z(n375) );
  INV_X1 U407 ( .A(n375), .ZN(n570) );
  NOR2_X1 U408 ( .A1(n357), .A2(n570), .ZN(n373) );
  XOR2_X1 U409 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n359) );
  XNOR2_X1 U410 ( .A(G99GAT), .B(KEYINPUT9), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U412 ( .A(G50GAT), .B(G162GAT), .Z(n415) );
  XOR2_X1 U413 ( .A(n360), .B(n415), .Z(n363) );
  XOR2_X1 U414 ( .A(G43GAT), .B(G134GAT), .Z(n428) );
  XNOR2_X1 U415 ( .A(n361), .B(n428), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U417 ( .A(n364), .B(KEYINPUT72), .Z(n367) );
  XNOR2_X1 U418 ( .A(G218GAT), .B(n365), .ZN(n366) );
  XNOR2_X1 U419 ( .A(n367), .B(n366), .ZN(n372) );
  XOR2_X1 U420 ( .A(G106GAT), .B(KEYINPUT66), .Z(n369) );
  NAND2_X1 U421 ( .A1(G232GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U423 ( .A(G190GAT), .B(n370), .Z(n371) );
  XOR2_X1 U424 ( .A(n372), .B(n371), .Z(n558) );
  INV_X1 U425 ( .A(n558), .ZN(n461) );
  NAND2_X1 U426 ( .A1(n373), .A2(n461), .ZN(n374) );
  XNOR2_X1 U427 ( .A(KEYINPUT47), .B(n374), .ZN(n381) );
  XOR2_X1 U428 ( .A(KEYINPUT36), .B(n558), .Z(n573) );
  NOR2_X1 U429 ( .A1(n573), .A2(n375), .ZN(n376) );
  XNOR2_X1 U430 ( .A(KEYINPUT45), .B(n376), .ZN(n378) );
  NAND2_X1 U431 ( .A1(n378), .A2(n334), .ZN(n379) );
  NOR2_X1 U432 ( .A1(n563), .A2(n379), .ZN(n380) );
  NOR2_X1 U433 ( .A1(n381), .A2(n380), .ZN(n382) );
  XNOR2_X1 U434 ( .A(KEYINPUT48), .B(n382), .ZN(n539) );
  NOR2_X1 U435 ( .A1(n510), .A2(n539), .ZN(n383) );
  XNOR2_X1 U436 ( .A(n383), .B(KEYINPUT54), .ZN(n407) );
  XOR2_X1 U437 ( .A(G57GAT), .B(G148GAT), .Z(n385) );
  XNOR2_X1 U438 ( .A(G1GAT), .B(G120GAT), .ZN(n384) );
  XNOR2_X1 U439 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U440 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n387) );
  XNOR2_X1 U441 ( .A(KEYINPUT6), .B(KEYINPUT92), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U443 ( .A(n389), .B(n388), .Z(n394) );
  XOR2_X1 U444 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n391) );
  NAND2_X1 U445 ( .A1(G225GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U447 ( .A(KEYINPUT5), .B(n392), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n400) );
  XOR2_X1 U449 ( .A(G85GAT), .B(G162GAT), .Z(n398) );
  XOR2_X1 U450 ( .A(G127GAT), .B(KEYINPUT0), .Z(n396) );
  XNOR2_X1 U451 ( .A(G113GAT), .B(KEYINPUT77), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n396), .B(n395), .ZN(n435) );
  XNOR2_X1 U453 ( .A(n435), .B(G134GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U455 ( .A(n400), .B(n399), .Z(n406) );
  XNOR2_X1 U456 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n401), .B(KEYINPUT89), .ZN(n402) );
  XOR2_X1 U458 ( .A(n402), .B(KEYINPUT90), .Z(n404) );
  XNOR2_X1 U459 ( .A(G141GAT), .B(G155GAT), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n419) );
  XNOR2_X1 U461 ( .A(G29GAT), .B(n419), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n508) );
  NAND2_X1 U463 ( .A1(n407), .A2(n508), .ZN(n561) );
  XOR2_X1 U464 ( .A(KEYINPUT24), .B(KEYINPUT86), .Z(n409) );
  XNOR2_X1 U465 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U467 ( .A(KEYINPUT85), .B(KEYINPUT91), .Z(n411) );
  XNOR2_X1 U468 ( .A(G22GAT), .B(G204GAT), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U470 ( .A(n413), .B(n412), .Z(n421) );
  XOR2_X1 U471 ( .A(n415), .B(n414), .Z(n417) );
  NAND2_X1 U472 ( .A1(G228GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n452) );
  NOR2_X1 U477 ( .A1(n561), .A2(n452), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n424), .B(KEYINPUT55), .ZN(n441) );
  XOR2_X1 U479 ( .A(KEYINPUT83), .B(KEYINPUT78), .Z(n426) );
  XNOR2_X1 U480 ( .A(G15GAT), .B(KEYINPUT82), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U482 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U483 ( .A1(G227GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U485 ( .A(G176GAT), .B(KEYINPUT20), .Z(n432) );
  XNOR2_X1 U486 ( .A(KEYINPUT65), .B(KEYINPUT79), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U488 ( .A(n434), .B(n433), .Z(n438) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n439) );
  NAND2_X1 U491 ( .A1(n563), .A2(n557), .ZN(n445) );
  XNOR2_X1 U492 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n443) );
  XOR2_X1 U493 ( .A(n510), .B(KEYINPUT95), .Z(n446) );
  XNOR2_X1 U494 ( .A(KEYINPUT27), .B(n446), .ZN(n454) );
  NOR2_X1 U495 ( .A1(n508), .A2(n454), .ZN(n447) );
  XOR2_X1 U496 ( .A(KEYINPUT96), .B(n447), .Z(n537) );
  XOR2_X1 U497 ( .A(KEYINPUT28), .B(n452), .Z(n516) );
  INV_X1 U498 ( .A(n516), .ZN(n448) );
  NOR2_X1 U499 ( .A1(n537), .A2(n448), .ZN(n522) );
  XNOR2_X1 U500 ( .A(KEYINPUT84), .B(n520), .ZN(n449) );
  NAND2_X1 U501 ( .A1(n522), .A2(n449), .ZN(n460) );
  NOR2_X1 U502 ( .A1(n510), .A2(n520), .ZN(n450) );
  NOR2_X1 U503 ( .A1(n452), .A2(n450), .ZN(n451) );
  XNOR2_X1 U504 ( .A(KEYINPUT25), .B(n451), .ZN(n457) );
  NAND2_X1 U505 ( .A1(n452), .A2(n520), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n453), .B(KEYINPUT26), .ZN(n562) );
  NOR2_X1 U507 ( .A1(n562), .A2(n454), .ZN(n455) );
  XNOR2_X1 U508 ( .A(KEYINPUT97), .B(n455), .ZN(n456) );
  NAND2_X1 U509 ( .A1(n457), .A2(n456), .ZN(n458) );
  NAND2_X1 U510 ( .A1(n508), .A2(n458), .ZN(n459) );
  NAND2_X1 U511 ( .A1(n460), .A2(n459), .ZN(n477) );
  XOR2_X1 U512 ( .A(KEYINPUT76), .B(KEYINPUT16), .Z(n463) );
  NAND2_X1 U513 ( .A1(n570), .A2(n461), .ZN(n462) );
  XNOR2_X1 U514 ( .A(n463), .B(n462), .ZN(n464) );
  NAND2_X1 U515 ( .A1(n477), .A2(n464), .ZN(n465) );
  XNOR2_X1 U516 ( .A(n465), .B(KEYINPUT98), .ZN(n493) );
  NAND2_X1 U517 ( .A1(n563), .A2(n334), .ZN(n481) );
  OR2_X1 U518 ( .A1(n493), .A2(n481), .ZN(n474) );
  NOR2_X1 U519 ( .A1(n508), .A2(n474), .ZN(n467) );
  XNOR2_X1 U520 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U522 ( .A(G1GAT), .B(n468), .ZN(G1324GAT) );
  NOR2_X1 U523 ( .A1(n510), .A2(n474), .ZN(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT100), .B(n469), .Z(n470) );
  XNOR2_X1 U525 ( .A(G8GAT), .B(n470), .ZN(G1325GAT) );
  NOR2_X1 U526 ( .A1(n520), .A2(n474), .ZN(n472) );
  XNOR2_X1 U527 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n471) );
  XNOR2_X1 U528 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U529 ( .A(G15GAT), .B(n473), .Z(G1326GAT) );
  NOR2_X1 U530 ( .A1(n516), .A2(n474), .ZN(n475) );
  XOR2_X1 U531 ( .A(KEYINPUT102), .B(n475), .Z(n476) );
  XNOR2_X1 U532 ( .A(G22GAT), .B(n476), .ZN(G1327GAT) );
  XNOR2_X1 U533 ( .A(KEYINPUT37), .B(KEYINPUT103), .ZN(n480) );
  NOR2_X1 U534 ( .A1(n573), .A2(n570), .ZN(n478) );
  NAND2_X1 U535 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U536 ( .A(n480), .B(n479), .ZN(n507) );
  NOR2_X1 U537 ( .A1(n507), .A2(n481), .ZN(n482) );
  XOR2_X1 U538 ( .A(KEYINPUT38), .B(n482), .Z(n483) );
  XNOR2_X1 U539 ( .A(KEYINPUT104), .B(n483), .ZN(n491) );
  NOR2_X1 U540 ( .A1(n508), .A2(n491), .ZN(n485) );
  XNOR2_X1 U541 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n485), .B(n484), .ZN(G1328GAT) );
  NOR2_X1 U543 ( .A1(n510), .A2(n491), .ZN(n487) );
  XNOR2_X1 U544 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(G1329GAT) );
  NOR2_X1 U546 ( .A1(n520), .A2(n491), .ZN(n489) );
  XNOR2_X1 U547 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U549 ( .A(G43GAT), .B(n490), .Z(G1330GAT) );
  NOR2_X1 U550 ( .A1(n516), .A2(n491), .ZN(n492) );
  XOR2_X1 U551 ( .A(G50GAT), .B(n492), .Z(G1331GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT107), .B(n541), .Z(n552) );
  NAND2_X1 U553 ( .A1(n523), .A2(n552), .ZN(n506) );
  OR2_X1 U554 ( .A1(n493), .A2(n506), .ZN(n502) );
  NOR2_X1 U555 ( .A1(n508), .A2(n502), .ZN(n495) );
  XNOR2_X1 U556 ( .A(KEYINPUT42), .B(KEYINPUT108), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U558 ( .A(G57GAT), .B(n496), .Z(G1332GAT) );
  NOR2_X1 U559 ( .A1(n510), .A2(n502), .ZN(n498) );
  XNOR2_X1 U560 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U562 ( .A(G64GAT), .B(n499), .ZN(G1333GAT) );
  NOR2_X1 U563 ( .A1(n520), .A2(n502), .ZN(n501) );
  XNOR2_X1 U564 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n501), .B(n500), .ZN(G1334GAT) );
  NOR2_X1 U566 ( .A1(n516), .A2(n502), .ZN(n504) );
  XNOR2_X1 U567 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U569 ( .A(G78GAT), .B(n505), .ZN(G1335GAT) );
  OR2_X1 U570 ( .A1(n507), .A2(n506), .ZN(n515) );
  NOR2_X1 U571 ( .A1(n508), .A2(n515), .ZN(n509) );
  XOR2_X1 U572 ( .A(G85GAT), .B(n509), .Z(G1336GAT) );
  NOR2_X1 U573 ( .A1(n510), .A2(n515), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G92GAT), .B(KEYINPUT113), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(G1337GAT) );
  NOR2_X1 U576 ( .A1(n520), .A2(n515), .ZN(n513) );
  XOR2_X1 U577 ( .A(KEYINPUT114), .B(n513), .Z(n514) );
  XNOR2_X1 U578 ( .A(G99GAT), .B(n514), .ZN(G1338GAT) );
  NOR2_X1 U579 ( .A1(n516), .A2(n515), .ZN(n518) );
  XNOR2_X1 U580 ( .A(KEYINPUT44), .B(KEYINPUT115), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U582 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  NOR2_X1 U583 ( .A1(n520), .A2(n539), .ZN(n521) );
  NAND2_X1 U584 ( .A1(n522), .A2(n521), .ZN(n526) );
  NOR2_X1 U585 ( .A1(n523), .A2(n526), .ZN(n525) );
  XNOR2_X1 U586 ( .A(G113GAT), .B(KEYINPUT117), .ZN(n524) );
  XNOR2_X1 U587 ( .A(n525), .B(n524), .ZN(G1340GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n528) );
  INV_X1 U589 ( .A(n526), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n533), .A2(n552), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U592 ( .A(G120GAT), .B(n529), .ZN(G1341GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n531) );
  NAND2_X1 U594 ( .A1(n533), .A2(n570), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(n532), .ZN(G1342GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n535) );
  NAND2_X1 U598 ( .A1(n533), .A2(n558), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G134GAT), .B(n536), .ZN(G1343GAT) );
  OR2_X1 U601 ( .A1(n562), .A2(n537), .ZN(n538) );
  NOR2_X1 U602 ( .A1(n539), .A2(n538), .ZN(n547) );
  AND2_X1 U603 ( .A1(n563), .A2(n547), .ZN(n540) );
  XOR2_X1 U604 ( .A(G141GAT), .B(n540), .Z(G1344GAT) );
  XOR2_X1 U605 ( .A(G148GAT), .B(KEYINPUT53), .Z(n543) );
  NAND2_X1 U606 ( .A1(n547), .A2(n541), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(n545) );
  XOR2_X1 U608 ( .A(KEYINPUT52), .B(KEYINPUT121), .Z(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1345GAT) );
  NAND2_X1 U610 ( .A1(n570), .A2(n547), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n546), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U612 ( .A1(n547), .A2(n558), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n548), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n550) );
  XNOR2_X1 U615 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U617 ( .A(KEYINPUT56), .B(n551), .Z(n554) );
  NAND2_X1 U618 ( .A1(n557), .A2(n552), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1349GAT) );
  NAND2_X1 U620 ( .A1(n570), .A2(n557), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(KEYINPUT126), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G183GAT), .B(n556), .ZN(G1350GAT) );
  XNOR2_X1 U623 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n560) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1351GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n565) );
  NOR2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n569), .A2(n563), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(n566), .ZN(G1352GAT) );
  XOR2_X1 U631 ( .A(G204GAT), .B(KEYINPUT61), .Z(n568) );
  INV_X1 U632 ( .A(n569), .ZN(n572) );
  OR2_X1 U633 ( .A1(n572), .A2(n334), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1353GAT) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT62), .B(n574), .Z(n575) );
  XNOR2_X1 U639 ( .A(G218GAT), .B(n575), .ZN(G1355GAT) );
endmodule

