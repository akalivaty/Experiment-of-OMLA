//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n203));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  NOR2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n205), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT24), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(G183gat), .A3(G190gat), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n213), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n203), .B1(new_n211), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(new_n215), .ZN(new_n220));
  XOR2_X1   g019(.A(KEYINPUT66), .B(G183gat), .Z(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n206), .A2(KEYINPUT65), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(KEYINPUT23), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n203), .B1(new_n207), .B2(new_n208), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n222), .A2(new_n226), .A3(new_n205), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n219), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT26), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n223), .A2(new_n230), .A3(new_n225), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n205), .B(new_n231), .C1(new_n230), .C2(new_n206), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(new_n233), .A3(new_n212), .ZN(new_n234));
  OR2_X1    g033(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n236));
  NAND2_X1  g035(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n236), .B1(new_n235), .B2(new_n237), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT28), .B1(new_n240), .B2(G190gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n221), .A2(KEYINPUT27), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n235), .ZN(new_n243));
  NOR2_X1   g042(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n234), .A2(new_n241), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n233), .B1(new_n232), .B2(new_n212), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n229), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(G226gat), .A2(G233gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n212), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT68), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n252), .A2(new_n234), .A3(new_n245), .A4(new_n241), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT29), .B1(new_n253), .B2(new_n229), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n250), .B1(new_n254), .B2(new_n249), .ZN(new_n255));
  XNOR2_X1  g054(.A(G197gat), .B(G204gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT22), .ZN(new_n257));
  INV_X1    g056(.A(G211gat), .ZN(new_n258));
  INV_X1    g057(.A(G218gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G211gat), .B(G218gat), .Z(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n255), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n250), .B(new_n263), .C1(new_n254), .C2(new_n249), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G8gat), .B(G36gat), .Z(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT73), .ZN(new_n269));
  XNOR2_X1  g068(.A(G64gat), .B(G92gat), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n269), .B(new_n270), .Z(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n202), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT30), .A4(new_n271), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n267), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT72), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n275), .B1(new_n272), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G15gat), .B(G43gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(G71gat), .B(G99gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G227gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G113gat), .B(G120gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(KEYINPUT1), .ZN(new_n287));
  XOR2_X1   g086(.A(G127gat), .B(G134gat), .Z(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n289), .B(new_n229), .C1(new_n246), .C2(new_n247), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n289), .B1(new_n253), .B2(new_n229), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n285), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n283), .B1(new_n293), .B2(KEYINPUT32), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT33), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n298));
  INV_X1    g097(.A(new_n289), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n248), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n284), .B1(new_n300), .B2(new_n290), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n283), .A2(new_n295), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n298), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n293), .A2(new_n298), .A3(KEYINPUT32), .A4(new_n305), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n297), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n300), .A2(new_n284), .A3(new_n290), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n312), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G78gat), .B(G106gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT31), .B(G50gat), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n317), .B(new_n318), .Z(new_n319));
  XOR2_X1   g118(.A(new_n319), .B(KEYINPUT80), .Z(new_n320));
  NAND2_X1  g119(.A1(G228gat), .A2(G233gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322));
  XNOR2_X1  g121(.A(G141gat), .B(G148gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(KEYINPUT2), .ZN(new_n324));
  INV_X1    g123(.A(G155gat), .ZN(new_n325));
  INV_X1    g124(.A(G162gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n324), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n327), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT2), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  OR2_X1    g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n336));
  NAND2_X1  g135(.A1(G141gat), .A2(G148gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n336), .B1(new_n335), .B2(new_n337), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n334), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(KEYINPUT75), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n323), .A2(KEYINPUT74), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n338), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n343), .B1(new_n345), .B2(new_n334), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n322), .B(new_n330), .C1(new_n342), .C2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n263), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT81), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n321), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n341), .A2(KEYINPUT75), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n345), .A2(new_n343), .A3(new_n334), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n329), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT3), .B1(new_n263), .B2(new_n348), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n347), .A2(new_n348), .ZN(new_n359));
  AOI221_X4 g158(.A(new_n356), .B1(new_n350), .B2(new_n321), .C1(new_n359), .C2(new_n264), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n358), .A2(new_n360), .A3(G22gat), .ZN(new_n361));
  INV_X1    g160(.A(G22gat), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT29), .B1(new_n354), .B2(new_n322), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT81), .B1(new_n363), .B2(new_n263), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n364), .B(new_n321), .C1(new_n349), .C2(new_n356), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n351), .A2(new_n357), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n320), .B1(new_n361), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n369), .B(G22gat), .C1(new_n358), .C2(new_n360), .ZN(new_n370));
  INV_X1    g169(.A(new_n319), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n365), .B(new_n366), .C1(KEYINPUT82), .C2(new_n362), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n293), .A2(KEYINPUT32), .A3(new_n305), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT69), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n376), .A2(new_n307), .B1(new_n296), .B2(new_n294), .ZN(new_n377));
  INV_X1    g176(.A(new_n315), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n316), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n354), .A2(new_n289), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n354), .A2(KEYINPUT4), .A3(new_n289), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT77), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n299), .B1(new_n354), .B2(new_n322), .ZN(new_n389));
  INV_X1    g188(.A(new_n347), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT76), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n330), .B1(new_n342), .B2(new_n346), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n289), .B1(new_n393), .B2(KEYINPUT3), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT76), .B1(new_n394), .B2(new_n347), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n385), .B(new_n388), .C1(new_n392), .C2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT5), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n393), .A2(new_n299), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n381), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n397), .B1(new_n399), .B2(new_n387), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n384), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n391), .B1(new_n389), .B2(new_n390), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n394), .A2(KEYINPUT76), .A3(new_n347), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(new_n397), .A3(new_n388), .ZN(new_n406));
  XOR2_X1   g205(.A(G1gat), .B(G29gat), .Z(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G57gat), .B(G85gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n401), .A2(new_n406), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n413), .A2(KEYINPUT79), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT79), .B1(new_n413), .B2(new_n414), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n412), .B1(new_n401), .B2(new_n406), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(KEYINPUT6), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n280), .B(new_n380), .C1(new_n418), .C2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT35), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n413), .A2(new_n414), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n419), .B1(new_n423), .B2(new_n417), .ZN(new_n424));
  AND4_X1   g223(.A1(new_n422), .A2(new_n280), .A3(new_n424), .A4(new_n374), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT71), .B1(new_n316), .B2(new_n379), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT71), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n427), .B1(new_n377), .B2(new_n378), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n421), .A2(KEYINPUT35), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n279), .A2(new_n272), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(new_n273), .A3(new_n274), .ZN(new_n432));
  OR3_X1    g231(.A1(new_n405), .A2(KEYINPUT39), .A3(new_n388), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n398), .A2(new_n388), .A3(new_n381), .ZN(new_n434));
  OAI211_X1 g233(.A(KEYINPUT39), .B(new_n434), .C1(new_n405), .C2(new_n388), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n412), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT40), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n417), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n437), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n432), .A2(new_n438), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT84), .B(KEYINPUT38), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT37), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n443), .B1(new_n277), .B2(new_n278), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n272), .B1(new_n267), .B2(KEYINPUT37), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n439), .A2(new_n414), .A3(new_n413), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n267), .A2(new_n272), .ZN(new_n448));
  INV_X1    g247(.A(new_n445), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n442), .B1(new_n267), .B2(KEYINPUT37), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n446), .A2(new_n447), .A3(new_n451), .A4(new_n419), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n441), .A2(new_n452), .A3(new_n374), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT36), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n455), .B1(new_n426), .B2(new_n428), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n316), .A2(new_n379), .A3(KEYINPUT36), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n374), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT79), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n417), .B1(new_n423), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n413), .A2(KEYINPUT79), .A3(new_n414), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n420), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n459), .B1(new_n463), .B2(new_n432), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n454), .B1(new_n465), .B2(KEYINPUT83), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT83), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n458), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n430), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NOR3_X1   g270(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n472));
  INV_X1    g271(.A(G29gat), .ZN(new_n473));
  INV_X1    g272(.A(G36gat), .ZN(new_n474));
  OAI22_X1  g273(.A1(new_n471), .A2(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G43gat), .B(G50gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(KEYINPUT15), .A3(new_n476), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n476), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(KEYINPUT15), .B2(new_n476), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT86), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n472), .A2(new_n480), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n471), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n477), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT17), .ZN(new_n485));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT16), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n486), .B1(new_n487), .B2(G1gat), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(G1gat), .B2(new_n486), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(G8gat), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G229gat), .A2(G233gat), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n493), .B(KEYINPUT87), .Z(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(new_n484), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT18), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n490), .B(new_n484), .ZN(new_n499));
  XOR2_X1   g298(.A(new_n494), .B(KEYINPUT13), .Z(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n496), .A2(new_n497), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G113gat), .B(G141gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT85), .B(G197gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(KEYINPUT11), .B(G169gat), .Z(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT12), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n498), .A2(new_n501), .A3(new_n502), .A4(new_n509), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n469), .A2(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(G120gat), .B(G148gat), .Z(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT97), .ZN(new_n517));
  XNOR2_X1  g316(.A(G176gat), .B(G204gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G230gat), .A2(G233gat), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT89), .ZN(new_n523));
  XNOR2_X1  g322(.A(G71gat), .B(G78gat), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n526));
  INV_X1    g325(.A(G57gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(G64gat), .ZN(new_n528));
  INV_X1    g327(.A(G64gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(G57gat), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n526), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT88), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n523), .B(new_n525), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G71gat), .A2(G78gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n529), .A2(G57gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n527), .A2(G64gat), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT89), .B1(new_n539), .B2(KEYINPUT88), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n524), .B1(new_n531), .B2(new_n523), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n533), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT91), .ZN(new_n544));
  INV_X1    g343(.A(G92gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G85gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(KEYINPUT91), .A2(G92gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(G99gat), .ZN(new_n550));
  INV_X1    g349(.A(G106gat), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT8), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(KEYINPUT90), .A2(G85gat), .A3(G92gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT7), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(KEYINPUT90), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n549), .A2(new_n552), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G99gat), .B(G106gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(KEYINPUT92), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n559), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n555), .A2(new_n556), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n562), .A2(new_n558), .A3(new_n552), .A4(new_n549), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n543), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT95), .B(KEYINPUT10), .Z(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n569));
  AND4_X1   g368(.A1(new_n569), .A2(new_n542), .A3(new_n561), .A4(new_n563), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n561), .A2(new_n563), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n569), .B1(new_n571), .B2(new_n542), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n566), .B(new_n568), .C1(new_n570), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n565), .A2(new_n560), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(KEYINPUT10), .A3(new_n542), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n522), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n566), .B1(new_n570), .B2(new_n572), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n577), .A2(new_n522), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n520), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT98), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT99), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT96), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n577), .A2(new_n583), .A3(new_n522), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n519), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n583), .B1(new_n577), .B2(new_n522), .ZN(new_n586));
  NOR3_X1   g385(.A1(new_n585), .A2(new_n576), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n581), .A2(new_n582), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n582), .B1(new_n581), .B2(new_n588), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n542), .A2(KEYINPUT21), .ZN(new_n593));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G127gat), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n490), .B1(KEYINPUT21), .B2(new_n542), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G155gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(G183gat), .B(G211gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n485), .A2(new_n560), .A3(new_n565), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n574), .A2(new_n484), .ZN(new_n607));
  NAND3_X1  g406(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G190gat), .B(G218gat), .Z(new_n610));
  AND2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  XOR2_X1   g411(.A(G134gat), .B(G162gat), .Z(new_n613));
  AOI21_X1  g412(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(KEYINPUT93), .Z(new_n616));
  OR3_X1    g415(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(KEYINPUT93), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(new_n611), .B2(new_n612), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n592), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n515), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n461), .A2(new_n462), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n419), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT100), .B(G1gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(G1324gat));
  NAND3_X1  g428(.A1(new_n515), .A2(new_n432), .A3(new_n623), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n630), .A2(G8gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT101), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G8gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT42), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(KEYINPUT42), .B2(new_n634), .ZN(G1325gat));
  OAI21_X1  g435(.A(G15gat), .B1(new_n624), .B2(new_n458), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n376), .A2(new_n307), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n638), .A2(new_n378), .A3(new_n297), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n378), .B1(new_n638), .B2(new_n297), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n427), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n428), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n643), .A2(G15gat), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n637), .B1(new_n624), .B2(new_n644), .ZN(G1326gat));
  NAND2_X1  g444(.A1(new_n515), .A2(new_n459), .ZN(new_n646));
  INV_X1    g445(.A(new_n623), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT43), .B(G22gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(G1327gat));
  NOR2_X1   g449(.A1(new_n469), .A2(new_n621), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n592), .A2(new_n605), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n514), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n655), .A2(new_n473), .A3(new_n463), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT45), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT44), .B1(new_n469), .B2(new_n621), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n421), .A2(KEYINPUT35), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n425), .A2(new_n429), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n458), .A2(new_n464), .A3(new_n453), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n659), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n662), .A2(new_n659), .A3(new_n663), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n665), .A2(new_n666), .A3(new_n620), .A4(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n658), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n654), .ZN(new_n670));
  OAI21_X1  g469(.A(G29gat), .B1(new_n670), .B2(new_n626), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n657), .A2(new_n671), .ZN(G1328gat));
  NAND3_X1  g471(.A1(new_n655), .A2(new_n474), .A3(new_n432), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(KEYINPUT46), .Z(new_n674));
  OAI21_X1  g473(.A(G36gat), .B1(new_n670), .B2(new_n280), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(G1329gat));
  NOR2_X1   g475(.A1(new_n643), .A2(G43gat), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n651), .A2(new_n654), .A3(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(KEYINPUT103), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(KEYINPUT103), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT47), .ZN(new_n681));
  AOI22_X1  g480(.A1(new_n679), .A2(new_n680), .B1(KEYINPUT104), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n681), .A2(KEYINPUT104), .ZN(new_n683));
  OAI21_X1  g482(.A(G43gat), .B1(new_n670), .B2(new_n458), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n683), .B1(new_n682), .B2(new_n684), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(G1330gat));
  OAI21_X1  g486(.A(G50gat), .B1(new_n670), .B2(new_n374), .ZN(new_n688));
  OR3_X1    g487(.A1(new_n653), .A2(G50gat), .A3(new_n621), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n688), .B1(new_n646), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT48), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1331gat));
  INV_X1    g491(.A(new_n667), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n664), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n622), .A2(new_n513), .A3(new_n591), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n463), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT105), .B(G57gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1332gat));
  INV_X1    g498(.A(new_n696), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n280), .ZN(new_n701));
  NOR2_X1   g500(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n702));
  AND2_X1   g501(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n701), .B2(new_n702), .ZN(G1333gat));
  INV_X1    g504(.A(new_n457), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n643), .B2(new_n455), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n696), .A2(G71gat), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n429), .B(KEYINPUT107), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n700), .A2(new_n713), .ZN(new_n714));
  OAI22_X1  g513(.A1(new_n710), .A2(new_n711), .B1(G71gat), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g515(.A1(new_n696), .A2(new_n459), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g517(.A1(new_n605), .A2(new_n513), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n591), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n658), .B2(new_n668), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(G85gat), .B1(new_n724), .B2(new_n626), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n280), .B1(new_n418), .B2(new_n420), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n726), .A2(new_n459), .B1(new_n456), .B2(new_n457), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n727), .A2(new_n453), .B1(new_n660), .B2(new_n661), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n720), .A2(new_n621), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT51), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n662), .A2(new_n663), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT51), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n732), .A2(new_n733), .A3(new_n729), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n731), .A2(new_n592), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n735), .A2(new_n547), .A3(new_n463), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n725), .A2(new_n736), .ZN(G1336gat));
  AOI22_X1  g536(.A1(new_n723), .A2(new_n432), .B1(new_n546), .B2(new_n548), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n735), .A2(new_n545), .A3(new_n432), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT52), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n724), .B2(new_n280), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n546), .A2(new_n548), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n723), .A2(KEYINPUT108), .A3(new_n432), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n739), .A2(KEYINPUT52), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n740), .B1(new_n745), .B2(new_n746), .ZN(G1337gat));
  NAND3_X1  g546(.A1(new_n723), .A2(G99gat), .A3(new_n707), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n735), .A2(new_n429), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(G99gat), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT109), .ZN(G1338gat));
  AOI21_X1  g550(.A(new_n551), .B1(new_n723), .B2(new_n459), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n374), .A2(G106gat), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n731), .A2(new_n734), .A3(new_n592), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT110), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT53), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n374), .B1(new_n626), .B2(new_n280), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT83), .B1(new_n758), .B2(new_n707), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(new_n468), .A3(new_n453), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n662), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n666), .B1(new_n761), .B2(new_n620), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n620), .A2(new_n666), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n693), .A2(new_n664), .A3(new_n763), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n459), .B(new_n721), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G106gat), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n754), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n757), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  AOI211_X1 g569(.A(KEYINPUT111), .B(new_n768), .C1(new_n765), .C2(G106gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n756), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n756), .B(KEYINPUT112), .C1(new_n770), .C2(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(G1339gat));
  NOR2_X1   g575(.A1(new_n647), .A2(new_n513), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n605), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n576), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n573), .A2(new_n522), .A3(new_n575), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI211_X1 g584(.A(KEYINPUT54), .B(new_n522), .C1(new_n573), .C2(new_n575), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n786), .A2(new_n787), .A3(new_n519), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n573), .A2(new_n575), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(new_n782), .A3(new_n521), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT113), .B1(new_n790), .B2(new_n520), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n785), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n588), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n787), .B1(new_n786), .B2(new_n519), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n790), .A2(KEYINPUT113), .A3(new_n520), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n783), .A2(new_n784), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT55), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n780), .B1(new_n793), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n494), .B1(new_n492), .B2(new_n495), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n499), .A2(new_n500), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n508), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n512), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n617), .B2(new_n619), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n797), .B1(new_n788), .B2(new_n791), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n781), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n587), .B1(new_n796), .B2(new_n785), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n807), .A3(KEYINPUT114), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n799), .A2(new_n804), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n799), .A2(new_n513), .A3(new_n808), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n512), .B(new_n802), .C1(new_n589), .C2(new_n590), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n809), .B1(new_n812), .B2(new_n621), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n779), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI211_X1 g614(.A(KEYINPUT115), .B(new_n809), .C1(new_n812), .C2(new_n621), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n778), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n459), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n626), .A2(new_n432), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n429), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(G113gat), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n821), .A2(new_n822), .A3(new_n514), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n817), .A2(new_n463), .A3(new_n380), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n432), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n817), .A2(KEYINPUT116), .A3(new_n463), .A4(new_n380), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n513), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n823), .B1(new_n829), .B2(new_n822), .ZN(G1340gat));
  INV_X1    g629(.A(G120gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n831), .A3(new_n592), .ZN(new_n832));
  OAI21_X1  g631(.A(G120gat), .B1(new_n821), .B2(new_n591), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n832), .B1(new_n835), .B2(new_n836), .ZN(G1341gat));
  INV_X1    g636(.A(G127gat), .ZN(new_n838));
  OR3_X1    g637(.A1(new_n821), .A2(new_n838), .A3(new_n779), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n825), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n840), .A2(new_n280), .A3(new_n605), .A4(new_n827), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(KEYINPUT118), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n826), .A2(new_n843), .A3(new_n605), .A4(new_n827), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n838), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n839), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g647(.A(KEYINPUT119), .B(new_n839), .C1(new_n842), .C2(new_n845), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(G1342gat));
  INV_X1    g649(.A(G134gat), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n828), .A2(new_n851), .A3(new_n620), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n853));
  OAI21_X1  g652(.A(G134gat), .B1(new_n821), .B2(new_n621), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(G1343gat));
  AND2_X1   g655(.A1(new_n458), .A2(new_n820), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n459), .A2(KEYINPUT57), .ZN(new_n858));
  INV_X1    g657(.A(new_n805), .ZN(new_n859));
  XNOR2_X1  g658(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n513), .B(new_n807), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n620), .B1(new_n811), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n809), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n605), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(KEYINPUT121), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n777), .B1(new_n864), .B2(KEYINPUT121), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n858), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT57), .B1(new_n817), .B2(new_n459), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n857), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G141gat), .B1(new_n869), .B2(new_n514), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n458), .A2(new_n459), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(new_n432), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n817), .A2(new_n463), .A3(new_n872), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n514), .A2(G141gat), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g675(.A(new_n858), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n817), .A2(new_n877), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n804), .A2(new_n807), .A3(new_n806), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n779), .B1(new_n862), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n778), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n881), .B2(new_n459), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n857), .A2(new_n592), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT59), .B(G148gat), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT59), .B1(new_n873), .B2(new_n591), .ZN(new_n886));
  INV_X1    g685(.A(G148gat), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n591), .A2(KEYINPUT59), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n885), .B(new_n888), .C1(new_n869), .C2(new_n889), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT122), .ZN(G1345gat));
  OAI21_X1  g690(.A(G155gat), .B1(new_n869), .B2(new_n779), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n605), .A2(new_n325), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n873), .B2(new_n893), .ZN(G1346gat));
  OAI21_X1  g693(.A(new_n326), .B1(new_n873), .B2(new_n621), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n621), .A2(new_n326), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n895), .B1(new_n869), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT123), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n818), .A2(new_n463), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n900), .A2(new_n432), .A3(new_n380), .ZN(new_n901));
  AOI21_X1  g700(.A(G169gat), .B1(new_n901), .B2(new_n513), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n463), .A2(new_n280), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n819), .A2(new_n712), .A3(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(G169gat), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n904), .A2(new_n905), .A3(new_n514), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n902), .A2(new_n906), .ZN(G1348gat));
  INV_X1    g706(.A(G176gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n901), .A2(new_n908), .A3(new_n592), .ZN(new_n909));
  OAI21_X1  g708(.A(G176gat), .B1(new_n904), .B2(new_n591), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n911), .B(new_n912), .ZN(G1349gat));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(KEYINPUT60), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n914), .A2(KEYINPUT60), .ZN(new_n916));
  INV_X1    g715(.A(new_n240), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n917), .A3(new_n605), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n221), .B1(new_n904), .B2(new_n779), .ZN(new_n919));
  AOI211_X1 g718(.A(new_n915), .B(new_n916), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  AND4_X1   g719(.A1(new_n914), .A2(new_n918), .A3(KEYINPUT60), .A4(new_n919), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(G1350gat));
  NAND3_X1  g721(.A1(new_n901), .A2(new_n217), .A3(new_n620), .ZN(new_n923));
  OAI21_X1  g722(.A(G190gat), .B1(new_n904), .B2(new_n621), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n924), .A2(KEYINPUT61), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(KEYINPUT61), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1351gat));
  NOR2_X1   g726(.A1(new_n871), .A2(new_n280), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n900), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n929), .A2(G197gat), .A3(new_n514), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT126), .Z(new_n931));
  AND2_X1   g730(.A1(new_n458), .A2(new_n903), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n932), .B1(new_n878), .B2(new_n882), .ZN(new_n933));
  OAI21_X1  g732(.A(G197gat), .B1(new_n933), .B2(new_n514), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n931), .A2(new_n934), .ZN(G1352gat));
  NOR3_X1   g734(.A1(new_n929), .A2(G204gat), .A3(new_n591), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  OAI21_X1  g738(.A(G204gat), .B1(new_n933), .B2(new_n591), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G1353gat));
  OAI211_X1 g740(.A(new_n605), .B(new_n932), .C1(new_n878), .C2(new_n882), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943));
  OAI21_X1  g742(.A(G211gat), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n942), .A2(new_n943), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT63), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n946), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n948), .A2(new_n944), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n605), .A2(new_n258), .ZN(new_n951));
  OAI22_X1  g750(.A1(new_n947), .A2(new_n950), .B1(new_n929), .B2(new_n951), .ZN(G1354gat));
  OAI21_X1  g751(.A(G218gat), .B1(new_n933), .B2(new_n621), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n620), .A2(new_n259), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n929), .B2(new_n954), .ZN(G1355gat));
endmodule


