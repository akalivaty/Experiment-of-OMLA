//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n602,
    new_n605, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT67), .Z(new_n451));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  AND2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(G319));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(KEYINPUT3), .A3(new_n463), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n469), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  OR2_X1    g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n468), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n467), .A2(KEYINPUT70), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n478), .B1(new_n466), .B2(G2105), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n464), .A2(G2105), .A3(new_n465), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  OR2_X1    g058(.A1(new_n471), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n483), .A2(G124), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OR2_X1    g064(.A1(new_n471), .A2(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n482), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n471), .A2(G138), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n497));
  OR2_X1    g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n469), .A2(new_n496), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n464), .A2(new_n465), .A3(new_n496), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n502), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n495), .B1(new_n505), .B2(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n508), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n512));
  XOR2_X1   g087(.A(KEYINPUT6), .B(G651), .Z(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n511), .A2(new_n514), .ZN(G166));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  XOR2_X1   g092(.A(KEYINPUT5), .B(G543), .Z(new_n518));
  NOR2_X1   g093(.A1(new_n518), .A2(new_n513), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G89), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT74), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n513), .A2(KEYINPUT73), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n524), .A2(G543), .A3(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n528), .A2(G51), .B1(new_n508), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n523), .A2(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND2_X1  g107(.A1(new_n528), .A2(G52), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n510), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n519), .A2(G90), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  XOR2_X1   g113(.A(KEYINPUT75), .B(G81), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n519), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n524), .A2(G543), .A3(new_n527), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n543), .B(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n510), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND4_X1  g128(.A1(new_n524), .A2(G53), .A3(G543), .A4(new_n527), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n518), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G651), .B1(new_n519), .B2(G91), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G166), .ZN(G303));
  NAND2_X1  g136(.A1(new_n528), .A2(G49), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n519), .A2(G87), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(G288));
  AOI22_X1  g140(.A1(new_n508), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(new_n513), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n508), .A2(G61), .ZN(new_n569));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n510), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(KEYINPUT77), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n573));
  AOI211_X1 g148(.A(new_n573), .B(new_n510), .C1(new_n569), .C2(new_n570), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n568), .B1(new_n572), .B2(new_n574), .ZN(G305));
  AOI22_X1  g150(.A1(new_n528), .A2(G47), .B1(G85), .B2(new_n519), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT79), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n510), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n576), .A2(KEYINPUT79), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(KEYINPUT80), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n508), .A2(new_n525), .A3(G92), .ZN(new_n588));
  XOR2_X1   g163(.A(new_n588), .B(KEYINPUT10), .Z(new_n589));
  AOI22_X1  g164(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n510), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n528), .A2(G54), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n586), .A2(KEYINPUT80), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n587), .B1(new_n596), .B2(new_n597), .ZN(G284));
  AOI21_X1  g173(.A(new_n587), .B1(new_n596), .B2(new_n597), .ZN(G321));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n600));
  NOR2_X1   g175(.A1(G168), .A2(new_n595), .ZN(new_n601));
  AOI211_X1 g176(.A(new_n600), .B(new_n601), .C1(new_n595), .C2(G299), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(new_n600), .B2(new_n601), .ZN(G297));
  AOI21_X1  g178(.A(new_n602), .B1(new_n600), .B2(new_n601), .ZN(G280));
  INV_X1    g179(.A(new_n594), .ZN(new_n605));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n473), .A2(new_n469), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n480), .A2(G135), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n471), .A2(G111), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n483), .A2(G123), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n621), .A2(G2096), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(G2096), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n615), .A2(new_n622), .A3(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT83), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2427), .B(G2430), .Z(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n633), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  NOR2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT84), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  AND3_X1   g216(.A1(new_n640), .A2(G14), .A3(new_n641), .ZN(G401));
  XNOR2_X1  g217(.A(G2072), .B(G2078), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT17), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT85), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n644), .A2(new_n645), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n650), .B(new_n647), .C1(new_n643), .C2(new_n645), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n646), .A2(new_n643), .A3(new_n645), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT18), .Z(new_n653));
  NAND3_X1  g228(.A1(new_n649), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT86), .Z(new_n664));
  OR2_X1    g239(.A1(new_n664), .A2(KEYINPUT20), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(KEYINPUT20), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n659), .A2(KEYINPUT87), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n660), .A2(new_n661), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n658), .B2(new_n662), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n667), .B(new_n669), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n665), .A2(new_n666), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G229));
  NOR2_X1   g253(.A1(G16), .A2(G24), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n584), .B(KEYINPUT88), .Z(new_n680));
  AOI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(G16), .ZN(new_n681));
  INV_X1    g256(.A(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n483), .A2(G119), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n471), .A2(G107), .ZN(new_n685));
  OAI21_X1  g260(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n477), .A2(new_n479), .ZN(new_n687));
  INV_X1    g262(.A(G131), .ZN(new_n688));
  OAI221_X1 g263(.A(new_n684), .B1(new_n685), .B2(new_n686), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  MUX2_X1   g264(.A(G25), .B(new_n689), .S(G29), .Z(new_n690));
  XOR2_X1   g265(.A(KEYINPUT35), .B(G1991), .Z(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G288), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n695), .B2(G23), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT33), .B(G1976), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n697), .A2(new_n699), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n695), .A2(G22), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n695), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1971), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n695), .A2(G6), .ZN(new_n705));
  INV_X1    g280(.A(G305), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n695), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT32), .B(G1981), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NOR4_X1   g284(.A1(new_n700), .A2(new_n701), .A3(new_n704), .A4(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n693), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n683), .B(new_n712), .C1(new_n711), .C2(new_n710), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT36), .Z(new_n714));
  NAND3_X1  g289(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT25), .Z(new_n716));
  AOI22_X1  g291(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n717));
  INV_X1    g292(.A(G139), .ZN(new_n718));
  OAI221_X1 g293(.A(new_n716), .B1(new_n471), .B2(new_n717), .C1(new_n687), .C2(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G33), .B(new_n719), .S(G29), .Z(new_n720));
  NOR2_X1   g295(.A1(new_n720), .A2(G2072), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT90), .ZN(new_n722));
  INV_X1    g297(.A(G2090), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G35), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G162), .B2(new_n724), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT29), .Z(new_n727));
  OAI21_X1  g302(.A(new_n722), .B1(new_n723), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n723), .B2(new_n727), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n483), .A2(G129), .B1(G105), .B2(new_n473), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT91), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT26), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n480), .B2(G141), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(new_n724), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n724), .B2(G32), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT27), .B(G1996), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT92), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n695), .A2(G5), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G171), .B2(new_n695), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT93), .ZN(new_n744));
  INV_X1    g319(.A(G1961), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n738), .A2(new_n740), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n741), .A2(new_n746), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n695), .A2(G4), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n605), .B2(new_n695), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1348), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n695), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n695), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1966), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n720), .A2(G2072), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n757), .A2(G28), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n724), .B1(new_n757), .B2(G28), .ZN(new_n759));
  AND2_X1   g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  NOR2_X1   g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT24), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G34), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(G34), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n475), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(G2084), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n762), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n616), .A2(G29), .A3(new_n620), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n767), .A2(new_n768), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n756), .A2(new_n769), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n749), .A2(new_n752), .A3(new_n755), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n695), .A2(G20), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT23), .Z(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G299), .B2(G16), .ZN(new_n776));
  INV_X1    g351(.A(G1956), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n724), .A2(G26), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT28), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n483), .A2(G128), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n471), .A2(G116), .ZN(new_n782));
  OAI21_X1  g357(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n783));
  INV_X1    g358(.A(G140), .ZN(new_n784));
  OAI221_X1 g359(.A(new_n781), .B1(new_n782), .B2(new_n783), .C1(new_n687), .C2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n780), .B1(new_n785), .B2(G29), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2067), .ZN(new_n787));
  NOR2_X1   g362(.A1(G27), .A2(G29), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G164), .B2(G29), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n787), .B1(G2078), .B2(new_n789), .ZN(new_n790));
  AOI211_X1 g365(.A(new_n778), .B(new_n790), .C1(G2078), .C2(new_n789), .ZN(new_n791));
  NOR2_X1   g366(.A1(G16), .A2(G19), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n548), .B2(G16), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT89), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G1341), .Z(new_n795));
  NAND4_X1  g370(.A1(new_n729), .A2(new_n773), .A3(new_n791), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n714), .A2(new_n796), .ZN(G311));
  INV_X1    g372(.A(G311), .ZN(G150));
  AOI22_X1  g373(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(new_n510), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G93), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n520), .ZN(new_n804));
  INV_X1    g379(.A(G55), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n800), .A2(new_n801), .B1(new_n541), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G860), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT37), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n594), .A2(new_n606), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n548), .A2(new_n807), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n545), .A2(new_n547), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n804), .B2(new_n806), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n813), .B(new_n817), .Z(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n808), .B1(new_n819), .B2(KEYINPUT39), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n810), .B1(new_n820), .B2(new_n821), .ZN(G145));
  INV_X1    g397(.A(G37), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n503), .A2(new_n504), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n824), .A2(new_n506), .A3(new_n500), .ZN(new_n825));
  INV_X1    g400(.A(new_n495), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n785), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n735), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n719), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT96), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G118), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n831), .A2(new_n832), .B1(new_n834), .B2(G2105), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n483), .A2(G130), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G142), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n687), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n613), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n689), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT97), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n830), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n621), .B(new_n475), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n488), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n840), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n842), .B(new_n845), .C1(new_n830), .C2(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n830), .A2(new_n841), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(new_n842), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n823), .B(new_n847), .C1(new_n849), .C2(new_n845), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g426(.A1(new_n594), .A2(G299), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n594), .A2(G299), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT41), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT41), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n852), .A2(new_n857), .A3(new_n853), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n854), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(KEYINPUT98), .A3(new_n857), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n817), .B(new_n608), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n860), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(KEYINPUT100), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT100), .B1(new_n864), .B2(new_n865), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT42), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n584), .B(new_n706), .ZN(new_n869));
  XNOR2_X1  g444(.A(G288), .B(G166), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n869), .B(new_n870), .Z(new_n871));
  OAI21_X1  g446(.A(new_n868), .B1(new_n871), .B2(KEYINPUT99), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n869), .B(new_n870), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT42), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n866), .B1(new_n867), .B2(new_n876), .ZN(new_n877));
  MUX2_X1   g452(.A(new_n862), .B(new_n854), .S(new_n863), .Z(new_n878));
  NAND4_X1  g453(.A1(new_n878), .A2(KEYINPUT100), .A3(new_n872), .A4(new_n875), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(G868), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n807), .A2(G868), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n595), .B1(new_n877), .B2(new_n879), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT101), .B1(new_n886), .B2(new_n883), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(G295));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n881), .A2(new_n889), .A3(new_n884), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT102), .B1(new_n886), .B2(new_n883), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(G331));
  XOR2_X1   g467(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n893));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n814), .A2(G301), .A3(new_n816), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(G301), .B1(new_n814), .B2(new_n816), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n896), .A2(new_n897), .A3(G286), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n817), .A2(G171), .ZN(new_n899));
  AOI21_X1  g474(.A(G168), .B1(new_n899), .B2(new_n895), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n860), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(G286), .B1(new_n896), .B2(new_n897), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(G168), .A3(new_n895), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n902), .A2(new_n903), .A3(new_n861), .A4(new_n859), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n871), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n823), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n871), .B1(new_n901), .B2(new_n904), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n854), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n855), .A2(new_n910), .A3(new_n858), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n902), .A2(new_n903), .A3(new_n909), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n901), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n873), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n914), .A2(new_n915), .A3(new_n823), .A4(new_n905), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n894), .B1(new_n908), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n907), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n918), .A2(new_n823), .A3(new_n905), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT104), .B1(new_n919), .B2(KEYINPUT43), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n893), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n914), .A2(new_n823), .A3(new_n905), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT106), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n914), .A2(new_n924), .A3(new_n823), .A4(new_n905), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(KEYINPUT43), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n906), .A2(new_n907), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(new_n915), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n921), .A2(new_n930), .ZN(G397));
  AOI21_X1  g506(.A(G1384), .B1(new_n825), .B2(new_n826), .ZN(new_n932));
  XOR2_X1   g507(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n468), .A2(new_n472), .A3(G40), .A4(new_n474), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT109), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n785), .B(G2067), .Z(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n735), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT127), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n938), .A2(G1996), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(KEYINPUT46), .Z(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT47), .ZN(new_n947));
  INV_X1    g522(.A(G1996), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n940), .B1(new_n948), .B2(new_n735), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n939), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n944), .A2(new_n735), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n689), .B(new_n692), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n952), .B1(new_n939), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n584), .A2(new_n682), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(new_n938), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT48), .Z(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n947), .A2(new_n958), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n689), .A2(new_n692), .ZN(new_n960));
  OAI22_X1  g535(.A1(new_n952), .A2(new_n960), .B1(G2067), .B2(new_n785), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT126), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n959), .B1(new_n939), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n933), .B1(G164), .B2(G1384), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n502), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT71), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n966), .A2(new_n967), .A3(new_n501), .ZN(new_n968));
  OAI211_X1 g543(.A(KEYINPUT45), .B(new_n965), .C1(new_n968), .C2(new_n495), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n964), .A2(new_n969), .A3(new_n937), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT110), .ZN(new_n971));
  INV_X1    g546(.A(G1971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n964), .A2(new_n969), .A3(new_n973), .A4(new_n937), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n965), .B1(new_n968), .B2(new_n495), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n936), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT111), .B1(new_n932), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n980));
  NOR4_X1   g555(.A1(G164), .A2(new_n980), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n977), .B(new_n723), .C1(new_n979), .C2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n975), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G8), .ZN(new_n984));
  NOR2_X1   g559(.A1(G166), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT55), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n986), .B(KEYINPUT112), .Z(new_n987));
  NAND3_X1  g562(.A1(new_n983), .A2(G8), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1981), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n990), .B(new_n568), .C1(new_n572), .C2(new_n574), .ZN(new_n991));
  OAI21_X1  g566(.A(G1981), .B1(new_n567), .B2(new_n571), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n993), .A2(KEYINPUT49), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n984), .B1(new_n932), .B2(new_n937), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n991), .A2(KEYINPUT49), .A3(new_n992), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n996), .A2(KEYINPUT113), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(KEYINPUT113), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n994), .B(new_n995), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n694), .A2(G1976), .ZN(new_n1000));
  INV_X1    g575(.A(G1976), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT52), .B1(G288), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n995), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n995), .A2(new_n1000), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT52), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n999), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n989), .A2(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n999), .A2(new_n1001), .A3(new_n694), .ZN(new_n1008));
  INV_X1    g583(.A(new_n991), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n995), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n984), .B1(new_n975), .B2(new_n982), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1006), .B1(new_n1012), .B2(new_n986), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT115), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1006), .B(new_n1015), .C1(new_n1012), .C2(new_n986), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT63), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n827), .A2(new_n965), .A3(new_n934), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(G164), .B2(G1384), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(new_n1021), .A3(new_n937), .ZN(new_n1022));
  INV_X1    g597(.A(G1966), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n977), .B(new_n768), .C1(new_n979), .C2(new_n981), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n937), .B1(new_n932), .B2(KEYINPUT45), .ZN(new_n1028));
  NOR3_X1   g603(.A1(G164), .A2(G1384), .A3(new_n933), .ZN(new_n1029));
  OAI211_X1 g604(.A(KEYINPUT114), .B(new_n1023), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(G8), .A3(G168), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n989), .A2(new_n1018), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1017), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n932), .A2(new_n978), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n977), .A2(new_n723), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n984), .B1(new_n975), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n988), .B(new_n1006), .C1(new_n986), .C2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1018), .B1(new_n1038), .B2(new_n1032), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1011), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT122), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT114), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1026), .A2(KEYINPUT122), .A3(new_n1027), .A4(new_n1030), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(G168), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(new_n984), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(G286), .A2(G8), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1047), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1051), .B1(new_n1031), .B2(G8), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT62), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1050), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n979), .A2(new_n981), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1961), .B1(new_n1059), .B2(new_n977), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1022), .A2(new_n1061), .A3(G2078), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n971), .A2(new_n974), .ZN(new_n1063));
  INV_X1    g638(.A(G2078), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(KEYINPUT124), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n1068));
  AOI21_X1  g643(.A(G2078), .B1(new_n971), .B2(new_n974), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1066), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI211_X1 g646(.A(new_n1060), .B(new_n1062), .C1(new_n1067), .C2(new_n1071), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1072), .A2(new_n1038), .A3(G301), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1052), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT62), .B1(new_n1074), .B2(new_n1056), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1058), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1040), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1956), .B1(new_n977), .B2(new_n1035), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT56), .B(G2072), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n970), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n555), .A2(new_n1084), .A3(new_n559), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1084), .B1(new_n555), .B2(new_n559), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT116), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1087), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(new_n1085), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1078), .B1(new_n1083), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n970), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n1080), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1096), .A2(new_n937), .A3(new_n1035), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n777), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1092), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1099), .A2(new_n1100), .A3(KEYINPUT117), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1093), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1348), .B1(new_n1059), .B2(new_n977), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n932), .A2(new_n937), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(G2067), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1102), .B1(new_n594), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1095), .A2(new_n1098), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT58), .B(G1341), .Z(new_n1111));
  NAND2_X1  g686(.A1(new_n1104), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n970), .B2(G1996), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1113), .A2(new_n1114), .A3(new_n548), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1114), .B1(new_n1113), .B2(new_n548), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1109), .A2(KEYINPUT61), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n1102), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1108), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT61), .B1(new_n1120), .B2(KEYINPUT118), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n1122));
  OAI22_X1  g697(.A1(new_n1079), .A2(new_n1082), .B1(new_n1087), .B2(new_n1086), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT118), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n1109), .A3(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1121), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1122), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1119), .B(KEYINPUT120), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1106), .A2(KEYINPUT60), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT60), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1131), .A2(KEYINPUT121), .A3(new_n605), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT121), .B1(new_n1131), .B2(new_n605), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1129), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1134), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1136), .A2(KEYINPUT60), .A3(new_n1106), .A4(new_n1132), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1128), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT119), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1121), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT120), .B1(new_n1142), .B2(new_n1119), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1110), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1060), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1064), .A2(KEYINPUT125), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1064), .A2(KEYINPUT125), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1094), .B(KEYINPUT53), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1146), .A2(G301), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1062), .ZN(new_n1151));
  AOI21_X1  g726(.A(G301), .B1(new_n1146), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1145), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1146), .A2(G301), .A3(new_n1151), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1060), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1155), .A2(new_n1156), .A3(new_n1149), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1154), .B(KEYINPUT54), .C1(new_n1157), .C2(G301), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1038), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1153), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1077), .B1(new_n1144), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(G290), .A2(G1986), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1162), .A2(KEYINPUT108), .A3(new_n955), .ZN(new_n1163));
  INV_X1    g738(.A(new_n938), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1163), .B(new_n1164), .C1(KEYINPUT108), .C2(new_n1162), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n954), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n963), .B1(new_n1161), .B2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g742(.A1(new_n917), .A2(new_n920), .ZN(new_n1169));
  INV_X1    g743(.A(new_n458), .ZN(new_n1170));
  NOR3_X1   g744(.A1(G401), .A2(new_n1170), .A3(G227), .ZN(new_n1171));
  NAND3_X1  g745(.A1(new_n850), .A2(new_n677), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n1169), .A2(new_n1172), .ZN(G308));
  AND2_X1   g747(.A1(new_n1171), .A2(new_n677), .ZN(new_n1174));
  OAI211_X1 g748(.A(new_n1174), .B(new_n850), .C1(new_n917), .C2(new_n920), .ZN(G225));
endmodule


