//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1297,
    new_n1298, new_n1299, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n214), .B1(new_n203), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n213), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT65), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  AND2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  INV_X1    g0026(.A(G50), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n206), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n211), .ZN(new_n230));
  AND2_X1   g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n213), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT0), .Z(new_n234));
  NOR4_X1   g0034(.A1(new_n225), .A2(new_n226), .A3(new_n231), .A4(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G226), .B(G232), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n227), .A2(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n203), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n249), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1698), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G222), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G223), .A3(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G77), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n261), .B(new_n263), .C1(new_n264), .C2(new_n262), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G1), .A3(G13), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(G274), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI22_X1  g0077(.A1(G226), .A2(new_n272), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n267), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT68), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n279), .A2(new_n280), .ZN(new_n283));
  OAI21_X1  g0083(.A(G190), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n283), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G200), .A3(new_n281), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n229), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT69), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n290), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT8), .B(G58), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n257), .A2(G20), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G150), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n211), .B1(new_n206), .B2(new_n227), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n289), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G13), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n302), .A2(new_n211), .A3(G1), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G50), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n289), .B1(new_n210), .B2(G20), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(G50), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n308), .A2(KEYINPUT9), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(KEYINPUT9), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n287), .B(new_n311), .C1(KEYINPUT71), .C2(KEYINPUT10), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n284), .B(new_n286), .C1(new_n309), .C2(new_n310), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT71), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G179), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n282), .B2(new_n283), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n285), .A2(new_n319), .A3(new_n281), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n320), .A3(new_n308), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n312), .A2(new_n316), .A3(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n323), .A2(G20), .B1(G159), .B2(new_n297), .ZN(new_n324));
  AND2_X1   g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT75), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT75), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n258), .A2(new_n328), .A3(new_n259), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n329), .A3(new_n211), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT7), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n262), .A2(G20), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n330), .A2(new_n331), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(KEYINPUT16), .B(new_n324), .C1(new_n335), .C2(new_n203), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT16), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n323), .A2(G20), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n297), .A2(G159), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n333), .B1(new_n262), .B2(G20), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n259), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n203), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n337), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n336), .A2(new_n289), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n306), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n293), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n303), .B2(new_n293), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  OR2_X1    g0149(.A1(G223), .A2(G1698), .ZN(new_n350));
  INV_X1    g0150(.A(G226), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G1698), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n350), .B(new_n352), .C1(new_n325), .C2(new_n326), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G87), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT77), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT77), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n353), .A2(new_n357), .A3(new_n354), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n356), .A2(new_n266), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n277), .A2(new_n269), .A3(G274), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n269), .A2(G232), .A3(new_n270), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n361), .A3(KEYINPUT78), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT78), .B1(new_n360), .B2(new_n361), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(G169), .B1(new_n359), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n356), .A2(new_n266), .A3(new_n358), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n360), .A2(new_n361), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT78), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n362), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n367), .A2(new_n371), .A3(G179), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n349), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT18), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n345), .A2(new_n348), .B1(new_n366), .B2(new_n372), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT18), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n367), .A2(new_n371), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(G190), .ZN(new_n380));
  AOI21_X1  g0180(.A(G200), .B1(new_n367), .B2(new_n371), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n345), .B(new_n348), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT17), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(G190), .B2(new_n379), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n387), .A2(KEYINPUT17), .A3(new_n345), .A4(new_n348), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n375), .A2(new_n378), .A3(new_n384), .A4(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n322), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT13), .ZN(new_n391));
  OAI211_X1 g0191(.A(G232), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT72), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n262), .A2(KEYINPUT72), .A3(G232), .A4(G1698), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G97), .ZN(new_n396));
  INV_X1    g0196(.A(G1698), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n262), .A2(G226), .A3(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n394), .A2(new_n395), .A3(new_n396), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n266), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n360), .B1(new_n215), .B2(new_n271), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n391), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  AOI211_X1 g0203(.A(KEYINPUT13), .B(new_n401), .C1(new_n399), .C2(new_n266), .ZN(new_n404));
  OAI21_X1  g0204(.A(G169), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n403), .A2(new_n404), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n405), .A2(KEYINPUT14), .B1(new_n406), .B2(G179), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT14), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n408), .B(G169), .C1(new_n403), .C2(new_n404), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT74), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n409), .A2(new_n410), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n407), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n306), .A2(G68), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT12), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n304), .B2(G68), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n303), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT73), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n294), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(new_n264), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n298), .A2(new_n227), .B1(new_n211), .B2(G68), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n289), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT11), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n414), .A2(new_n416), .A3(KEYINPUT73), .A4(new_n417), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n425), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n420), .A2(new_n426), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n413), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(G200), .B1(new_n403), .B2(new_n404), .ZN(new_n431));
  INV_X1    g0231(.A(new_n429), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n400), .A2(new_n402), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT13), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n400), .A2(new_n391), .A3(new_n402), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(G190), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n431), .B(new_n432), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n306), .A2(G77), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n303), .A2(new_n264), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n292), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n442), .A2(new_n297), .B1(G20), .B2(G77), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT15), .B(G87), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n443), .B1(new_n421), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n441), .B1(new_n445), .B2(new_n289), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n260), .A2(G232), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n262), .A2(G238), .A3(G1698), .ZN(new_n448));
  INV_X1    g0248(.A(G107), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n447), .B(new_n448), .C1(new_n449), .C2(new_n262), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n266), .ZN(new_n451));
  INV_X1    g0251(.A(G244), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n360), .B1(new_n452), .B2(new_n271), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT70), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n454), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n451), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n446), .B1(new_n457), .B2(new_n319), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n451), .A2(new_n455), .A3(new_n317), .A4(new_n456), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n457), .A2(G200), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n457), .A2(new_n437), .ZN(new_n463));
  INV_X1    g0263(.A(new_n446), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n461), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n430), .A2(new_n438), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n390), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n210), .A2(G45), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT5), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G41), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT79), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n473), .B1(new_n275), .B2(KEYINPUT5), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n275), .A2(KEYINPUT5), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n266), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(G257), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n479));
  OAI211_X1 g0279(.A(G250), .B(new_n397), .C1(new_n325), .C2(new_n326), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G294), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n478), .A2(G264), .B1(new_n482), .B2(new_n266), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n474), .A2(new_n477), .A3(G274), .A4(new_n269), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(KEYINPUT85), .A3(G179), .A4(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n319), .B1(new_n483), .B2(new_n484), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n482), .A2(new_n266), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT79), .B1(new_n471), .B2(G41), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(new_n472), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n276), .A2(G1), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n476), .B2(KEYINPUT79), .ZN(new_n491));
  OAI211_X1 g0291(.A(G264), .B(new_n269), .C1(new_n489), .C2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n487), .A2(G179), .A3(new_n492), .A4(new_n484), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT85), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n485), .B1(new_n486), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT86), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT86), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n498), .B(new_n485), .C1(new_n486), .C2(new_n495), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT84), .B1(new_n211), .B2(G107), .ZN(new_n500));
  OR2_X1    g0300(.A1(new_n500), .A2(KEYINPUT23), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(KEYINPUT23), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n501), .A2(new_n502), .B1(G116), .B2(new_n294), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT24), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n211), .B(G87), .C1(new_n325), .C2(new_n326), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT22), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT22), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n262), .A2(new_n507), .A3(new_n211), .A4(G87), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n503), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n504), .B1(new_n503), .B2(new_n509), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n289), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT25), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n304), .A2(new_n513), .A3(G107), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n304), .B2(G107), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n257), .A2(G1), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n303), .A2(new_n289), .A3(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n515), .A2(new_n516), .B1(G107), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n497), .A2(new_n499), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n483), .A2(new_n437), .A3(new_n484), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n487), .A2(new_n492), .A3(new_n484), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n385), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(new_n512), .A3(new_n519), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT19), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT80), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT80), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT19), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n396), .ZN(new_n532));
  AOI21_X1  g0332(.A(G20), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n216), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT81), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g0337(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n211), .B1(new_n538), .B2(new_n396), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT81), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(new_n535), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n294), .A2(G97), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n538), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n262), .A2(new_n211), .A3(G68), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n289), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n444), .A2(new_n303), .ZN(new_n548));
  OAI211_X1 g0348(.A(G238), .B(new_n397), .C1(new_n325), .C2(new_n326), .ZN(new_n549));
  OAI211_X1 g0349(.A(G244), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G116), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n266), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n470), .A2(G250), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n273), .A2(new_n470), .B1(new_n266), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n556), .A3(new_n437), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n555), .B1(new_n266), .B2(new_n552), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n557), .B1(new_n558), .B2(G200), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n518), .A2(G87), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n547), .A2(new_n548), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(G169), .B1(new_n553), .B2(new_n556), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n317), .B2(new_n558), .ZN(new_n563));
  INV_X1    g0363(.A(new_n444), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n518), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n546), .B1(new_n537), .B2(new_n541), .ZN(new_n566));
  INV_X1    g0366(.A(new_n289), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n548), .B(new_n565), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n526), .A2(new_n561), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n304), .A2(G97), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n518), .ZN(new_n573));
  INV_X1    g0373(.A(G97), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT6), .ZN(new_n576));
  AND2_X1   g0376(.A1(G97), .A2(G107), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(new_n534), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n449), .A2(KEYINPUT6), .A3(G97), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n580), .A2(G20), .B1(G77), .B2(new_n297), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n341), .A2(new_n342), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n582), .B2(new_n449), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n575), .B1(new_n583), .B2(new_n289), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n489), .A2(new_n491), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n478), .A2(G257), .B1(new_n585), .B2(new_n274), .ZN(new_n586));
  OAI211_X1 g0386(.A(G250), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G283), .ZN(new_n588));
  OAI211_X1 g0388(.A(G244), .B(new_n397), .C1(new_n325), .C2(new_n326), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n587), .B(new_n588), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT4), .B1(new_n260), .B2(G244), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n266), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n584), .B(new_n595), .C1(new_n437), .C2(new_n594), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n319), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n580), .A2(G20), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n297), .A2(G77), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n449), .B1(new_n341), .B2(new_n342), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n289), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n571), .B1(new_n518), .B2(G97), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n586), .A2(new_n593), .A3(new_n317), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n597), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n596), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n570), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(G270), .B(new_n269), .C1(new_n489), .C2(new_n491), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n484), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(G264), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n612));
  OAI211_X1 g0412(.A(G257), .B(new_n397), .C1(new_n325), .C2(new_n326), .ZN(new_n613));
  INV_X1    g0413(.A(G303), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n262), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n615), .A2(KEYINPUT82), .A3(new_n266), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT82), .B1(new_n615), .B2(new_n266), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n611), .B(G190), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n588), .B(new_n211), .C1(G33), .C2(new_n574), .ZN(new_n619));
  INV_X1    g0419(.A(G116), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G20), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n289), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT20), .ZN(new_n623));
  XNOR2_X1  g0423(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n303), .A2(KEYINPUT83), .A3(new_n620), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n210), .A2(new_n620), .A3(G13), .A4(G20), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT83), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n518), .A2(G116), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n615), .A2(new_n266), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT82), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n615), .A2(KEYINPUT82), .A3(new_n266), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n610), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n618), .B(new_n632), .C1(new_n637), .C2(new_n385), .ZN(new_n638));
  AOI211_X1 g0438(.A(new_n317), .B(new_n610), .C1(new_n624), .C2(new_n630), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n635), .A2(new_n636), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n611), .B1(new_n616), .B2(new_n617), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT21), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n319), .B1(new_n624), .B2(new_n630), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n642), .B2(new_n644), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n638), .B(new_n641), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n469), .A2(new_n521), .A3(new_n608), .A4(new_n649), .ZN(G372));
  XNOR2_X1  g0450(.A(new_n569), .B(KEYINPUT87), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n561), .A2(new_n569), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n652), .B1(new_n653), .B2(new_n606), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n548), .B(new_n560), .C1(new_n566), .C2(new_n567), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n656), .A2(new_n559), .B1(new_n568), .B2(new_n563), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n597), .A2(new_n604), .A3(new_n605), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(KEYINPUT26), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n651), .B1(new_n654), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n641), .B1(new_n646), .B2(new_n647), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n496), .B1(new_n512), .B2(new_n519), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n608), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n469), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n321), .ZN(new_n666));
  INV_X1    g0466(.A(new_n438), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n430), .B1(new_n667), .B2(new_n460), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n384), .A2(new_n388), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n349), .A2(new_n377), .A3(new_n373), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n377), .B1(new_n349), .B2(new_n373), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n312), .A2(new_n316), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n666), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n665), .A2(new_n676), .ZN(G369));
  NOR3_X1   g0477(.A1(new_n302), .A2(G1), .A3(G20), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT88), .ZN(new_n679));
  OR3_X1    g0479(.A1(new_n679), .A2(KEYINPUT89), .A3(KEYINPUT27), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT89), .B1(new_n679), .B2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(KEYINPUT90), .B(G343), .ZN(new_n683));
  INV_X1    g0483(.A(G213), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n684), .B1(new_n679), .B2(KEYINPUT27), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n521), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n526), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n520), .B2(new_n686), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n521), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n687), .A2(new_n632), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n661), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n648), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n647), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n700), .A2(new_n645), .B1(new_n640), .B2(new_n639), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n686), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n521), .A3(new_n690), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n662), .A2(new_n687), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n699), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT91), .ZN(G399));
  INV_X1    g0508(.A(new_n232), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n535), .A2(G116), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G1), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n228), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n711), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  NAND2_X1  g0516(.A1(new_n521), .A2(new_n701), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT93), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT93), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n521), .A2(new_n701), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n718), .A2(new_n608), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT87), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n569), .B(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT26), .B1(new_n657), .B2(new_n658), .ZN(new_n724));
  AND4_X1   g0524(.A1(KEYINPUT26), .A2(new_n658), .A3(new_n561), .A4(new_n569), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT92), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT92), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n660), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n721), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n687), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n686), .B1(new_n660), .B2(new_n663), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(KEYINPUT29), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G330), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n609), .A2(new_n484), .A3(G179), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n739), .A2(new_n483), .A3(new_n558), .ZN(new_n740));
  INV_X1    g0540(.A(new_n594), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(KEYINPUT30), .A3(new_n741), .A4(new_n640), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n558), .A2(G179), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n642), .A2(new_n743), .A3(new_n523), .A4(new_n594), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n593), .B(new_n586), .C1(new_n616), .C2(new_n617), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n739), .A2(new_n483), .A3(new_n558), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n742), .A2(new_n744), .A3(new_n748), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT31), .B1(new_n749), .B2(new_n686), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n608), .A2(new_n649), .A3(new_n521), .A4(new_n687), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n738), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n737), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n716), .B1(new_n756), .B2(new_n210), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT94), .ZN(G364));
  NOR2_X1   g0558(.A1(new_n302), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n210), .B1(new_n759), .B2(G45), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n710), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n229), .B1(G20), .B2(new_n319), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n254), .A2(new_n276), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n327), .A2(new_n329), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n709), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n276), .B2(new_n228), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n768), .B1(new_n772), .B2(KEYINPUT95), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(KEYINPUT95), .B2(new_n772), .ZN(new_n774));
  INV_X1    g0574(.A(new_n262), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n709), .A2(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n776), .A2(G355), .B1(new_n620), .B2(new_n709), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n766), .B(new_n767), .C1(new_n774), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(G20), .A2(G179), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n779), .A2(new_n385), .A3(G190), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(KEYINPUT33), .B(G317), .Z(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n779), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G311), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n775), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n211), .A2(G179), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n785), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n783), .B(new_n788), .C1(G329), .C2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n789), .A2(G190), .A3(G200), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT97), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G303), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n437), .A2(G179), .A3(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n211), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n784), .A2(G190), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G200), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n798), .A2(G294), .B1(new_n800), .B2(G322), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n789), .A2(new_n437), .A3(G200), .ZN(new_n802));
  INV_X1    g0602(.A(G283), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n799), .A2(new_n385), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(G326), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n792), .A2(new_n795), .A3(new_n801), .A4(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n802), .A2(new_n449), .ZN(new_n808));
  INV_X1    g0608(.A(new_n793), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n775), .B(new_n808), .C1(G87), .C2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT96), .Z(new_n811));
  NOR2_X1   g0611(.A1(new_n797), .A2(new_n574), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G50), .B2(new_n805), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n791), .A2(G159), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n814), .A2(KEYINPUT32), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n814), .A2(KEYINPUT32), .B1(G58), .B2(new_n800), .ZN(new_n816));
  INV_X1    g0616(.A(new_n786), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n817), .A2(G77), .B1(G68), .B2(new_n780), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n813), .A2(new_n815), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n807), .B1(new_n811), .B2(new_n819), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n763), .B(new_n778), .C1(new_n767), .C2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT98), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n766), .B(KEYINPUT99), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n696), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n697), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n762), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(G330), .B2(new_n696), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  INV_X1    g0629(.A(KEYINPUT101), .ZN(new_n830));
  AND3_X1   g0630(.A1(new_n458), .A2(new_n830), .A3(new_n459), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n830), .B1(new_n458), .B2(new_n459), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n465), .A2(new_n462), .B1(new_n686), .B2(new_n464), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT102), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n460), .B2(new_n687), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n686), .A2(new_n458), .A3(KEYINPUT102), .A4(new_n459), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n833), .A2(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n734), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n838), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n664), .A2(new_n687), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n754), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n711), .B2(new_n760), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n839), .A2(new_n754), .A3(new_n841), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n767), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n817), .A2(G159), .B1(G150), .B2(new_n780), .ZN(new_n847));
  INV_X1    g0647(.A(new_n800), .ZN(new_n848));
  INV_X1    g0648(.A(G143), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  INV_X1    g0650(.A(new_n805), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n847), .B1(new_n848), .B2(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT34), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n794), .A2(G50), .ZN(new_n856));
  INV_X1    g0656(.A(new_n769), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n797), .A2(new_n202), .B1(new_n802), .B2(new_n203), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n857), .B(new_n858), .C1(G132), .C2(new_n791), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n802), .A2(new_n216), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n851), .A2(new_n614), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n861), .B(new_n862), .C1(G294), .C2(new_n800), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n262), .B(new_n812), .C1(G311), .C2(new_n791), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n817), .A2(G116), .B1(G283), .B2(new_n780), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT100), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n794), .A2(G107), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n863), .A2(new_n864), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n846), .B1(new_n860), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n767), .A2(new_n764), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n763), .B(new_n869), .C1(new_n264), .C2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n840), .B2(new_n765), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n845), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(G384));
  OR2_X1    g0674(.A1(new_n580), .A2(KEYINPUT35), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n580), .A2(KEYINPUT35), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n875), .A2(G116), .A3(new_n230), .A4(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT36), .Z(new_n878));
  OAI211_X1 g0678(.A(new_n228), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n210), .B(G13), .C1(new_n879), .C2(new_n250), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n752), .A2(new_n753), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n840), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT103), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n434), .A2(G179), .A3(new_n435), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n319), .B1(new_n434), .B2(new_n435), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n885), .B1(new_n886), .B2(new_n408), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n409), .A2(new_n410), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(KEYINPUT74), .A3(new_n408), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n884), .B1(new_n890), .B2(new_n432), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n413), .A2(KEYINPUT103), .A3(new_n429), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n687), .A2(new_n432), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n667), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n407), .B(new_n438), .C1(new_n411), .C2(new_n412), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n893), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT104), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n896), .A2(KEYINPUT104), .A3(new_n893), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n883), .B1(new_n895), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n682), .A2(new_n685), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n349), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n669), .B2(new_n673), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n374), .A2(new_n905), .A3(new_n907), .A4(new_n382), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT105), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT37), .B1(new_n349), .B2(new_n904), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n911), .A2(KEYINPUT105), .A3(new_n374), .A4(new_n382), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n374), .A2(new_n905), .A3(new_n382), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n910), .A2(new_n912), .B1(KEYINPUT37), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n906), .B1(new_n914), .B2(KEYINPUT106), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(KEYINPUT37), .ZN(new_n916));
  INV_X1    g0716(.A(new_n349), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n376), .B1(new_n917), .B2(new_n387), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT105), .B1(new_n918), .B2(new_n911), .ZN(new_n919));
  INV_X1    g0719(.A(new_n912), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT106), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n915), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n330), .A2(new_n331), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n262), .A2(new_n333), .A3(G20), .ZN(new_n926));
  OAI21_X1  g0726(.A(G68), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT16), .B1(new_n927), .B2(new_n324), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n336), .A2(new_n289), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n348), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n373), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n904), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n932), .A3(new_n382), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT37), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n908), .ZN(new_n935));
  INV_X1    g0735(.A(new_n932), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n389), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n935), .A2(KEYINPUT38), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n902), .B(KEYINPUT40), .C1(new_n924), .C2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n901), .A2(new_n895), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT38), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n932), .B1(new_n669), .B2(new_n673), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n933), .A2(KEYINPUT37), .B1(new_n918), .B2(new_n911), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n938), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n838), .B1(new_n752), .B2(new_n753), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n941), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT40), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n940), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n468), .B1(new_n753), .B2(new_n752), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n953), .A2(new_n954), .A3(new_n738), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n833), .A2(new_n686), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n841), .A2(new_n957), .B1(new_n901), .B2(new_n895), .ZN(new_n958));
  INV_X1    g0758(.A(new_n673), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n958), .A2(new_n946), .B1(new_n959), .B2(new_n903), .ZN(new_n960));
  INV_X1    g0760(.A(new_n906), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n921), .B2(new_n922), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n914), .A2(KEYINPUT106), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n942), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT39), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n938), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n964), .A2(new_n967), .B1(KEYINPUT39), .B2(new_n946), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n891), .A2(new_n892), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n969), .A2(new_n686), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n960), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n676), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n737), .B2(new_n469), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n972), .B(new_n974), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n955), .A2(new_n975), .B1(new_n210), .B2(new_n759), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n955), .A2(new_n975), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n881), .B1(new_n976), .B2(new_n977), .ZN(G367));
  NOR2_X1   g0778(.A1(new_n766), .A2(new_n767), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n232), .B2(new_n444), .C1(new_n771), .C2(new_n245), .ZN(new_n980));
  INV_X1    g0780(.A(new_n794), .ZN(new_n981));
  OAI21_X1  g0781(.A(KEYINPUT46), .B1(new_n981), .B2(new_n620), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n620), .A2(KEYINPUT46), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n982), .B1(new_n793), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n802), .A2(new_n574), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G303), .B2(new_n800), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n449), .B2(new_n797), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G317), .A2(new_n791), .B1(new_n817), .B2(G283), .ZN(new_n988));
  INV_X1    g0788(.A(G294), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(new_n989), .B2(new_n781), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n857), .B1(new_n851), .B2(new_n787), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n987), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n984), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT111), .Z(new_n994));
  OAI22_X1  g0794(.A1(new_n851), .A2(new_n849), .B1(new_n793), .B2(new_n202), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G150), .B2(new_n800), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n790), .A2(new_n850), .B1(new_n786), .B2(new_n227), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n775), .B(new_n997), .C1(G159), .C2(new_n780), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n797), .A2(new_n203), .ZN(new_n999));
  INV_X1    g0799(.A(new_n802), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n999), .B1(G77), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n996), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n994), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT47), .Z(new_n1004));
  OAI211_X1 g0804(.A(new_n762), .B(new_n980), .C1(new_n1004), .C2(new_n846), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT112), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n651), .A2(new_n655), .A3(new_n686), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n657), .B1(new_n656), .B2(new_n687), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n823), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1007), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT110), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n607), .B1(new_n604), .B2(new_n686), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT108), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n687), .A2(new_n606), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT109), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n703), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT42), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n606), .B1(new_n1027), .B2(new_n521), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n687), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1010), .A2(KEYINPUT107), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1010), .A2(KEYINPUT107), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1030), .A2(new_n1031), .A3(KEYINPUT43), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1026), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT43), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1011), .A2(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1017), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n699), .A2(new_n1027), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1041));
  OAI211_X1 g0841(.A(KEYINPUT110), .B(new_n1033), .C1(new_n1041), .C2(new_n1037), .ZN(new_n1042));
  AND3_X1   g0842(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1040), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT45), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1027), .A2(new_n1046), .A3(new_n705), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT45), .B1(new_n1022), .B2(new_n706), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT44), .B1(new_n1027), .B2(new_n705), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT44), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1022), .A2(new_n706), .A3(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1047), .A2(new_n1048), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(new_n699), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n703), .B1(new_n692), .B2(new_n702), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(new_n825), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n755), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n756), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n710), .B(KEYINPUT41), .Z(new_n1059));
  OAI21_X1  g0859(.A(new_n760), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1016), .B1(new_n1045), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(G387));
  AOI22_X1  g0862(.A1(new_n798), .A2(new_n564), .B1(new_n800), .B2(G50), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT114), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n793), .A2(new_n264), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n985), .B(new_n1065), .C1(G159), .C2(new_n805), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n790), .A2(new_n296), .B1(new_n786), .B2(new_n203), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1067), .B(new_n857), .C1(new_n293), .C2(new_n780), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1064), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n769), .B1(G326), .B2(new_n791), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n797), .A2(new_n803), .B1(new_n793), .B2(new_n989), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n817), .A2(G303), .B1(G311), .B2(new_n780), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n800), .A2(G317), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(KEYINPUT115), .B(G322), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1072), .B(new_n1073), .C1(new_n851), .C2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT48), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1071), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n1076), .B2(new_n1075), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT49), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1070), .B1(new_n620), .B2(new_n802), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1069), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n767), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n712), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n776), .A2(new_n1084), .B1(new_n449), .B2(new_n709), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n241), .A2(new_n276), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n442), .A2(new_n227), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT50), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n712), .B(new_n276), .C1(new_n203), .C2(new_n264), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n770), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1085), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n763), .B1(new_n1091), .B2(new_n979), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT113), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1083), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n1093), .B2(new_n1092), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n693), .A2(new_n1012), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n761), .A2(new_n1055), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1056), .A2(new_n710), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n755), .A2(new_n1055), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(G393));
  NAND2_X1  g0900(.A1(new_n1027), .A2(new_n766), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G150), .A2(new_n805), .B1(new_n800), .B2(G159), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT51), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n781), .A2(new_n227), .B1(new_n790), .B2(new_n849), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n442), .B2(new_n817), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n857), .A2(new_n861), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n797), .A2(new_n264), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G68), .B2(new_n809), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(KEYINPUT116), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G311), .A2(new_n800), .B1(new_n805), .B2(G317), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT52), .Z(new_n1114));
  OAI22_X1  g0914(.A1(new_n790), .A2(new_n1074), .B1(new_n786), .B2(new_n989), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n262), .B(new_n1115), .C1(G303), .C2(new_n780), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n793), .A2(new_n803), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n808), .B(new_n1117), .C1(G116), .C2(new_n798), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1112), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1111), .A2(KEYINPUT116), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n767), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n979), .B1(new_n574), .B2(new_n232), .C1(new_n771), .C2(new_n249), .ZN(new_n1123));
  AND4_X1   g0923(.A1(new_n762), .A2(new_n1101), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1052), .B(new_n698), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1125), .B1(new_n1126), .B2(new_n760), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1056), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n711), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(G390));
  NAND3_X1  g0931(.A1(new_n730), .A2(new_n687), .A3(new_n840), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n957), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n941), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n970), .B1(new_n964), .B2(new_n938), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n841), .A2(new_n957), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n941), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n971), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n964), .A2(new_n967), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n946), .A2(KEYINPUT39), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n738), .B(new_n838), .C1(new_n752), .C2(new_n753), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n941), .A2(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1136), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n1136), .B2(new_n1142), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n968), .A2(new_n764), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n870), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n762), .B1(new_n293), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(G125), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n781), .A2(new_n850), .B1(new_n790), .B2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT54), .B(G143), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n775), .B(new_n1152), .C1(new_n817), .C2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n793), .A2(new_n296), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT53), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G128), .A2(new_n805), .B1(new_n1000), .B2(G50), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n798), .A2(G159), .B1(new_n800), .B2(G132), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT118), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n817), .A2(G97), .B1(G107), .B2(new_n780), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n803), .B2(new_n851), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT119), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n775), .B1(new_n790), .B2(new_n989), .C1(new_n203), .C2(new_n802), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1107), .B(new_n1166), .C1(G116), .C2(new_n800), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(new_n216), .C2(new_n981), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1162), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1150), .B1(new_n1170), .B2(new_n767), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1147), .A2(new_n761), .B1(new_n1148), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT117), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n956), .B1(new_n733), .B2(new_n840), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n895), .B(new_n901), .C1(new_n883), .C2(new_n738), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n1144), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1133), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1144), .A2(new_n1175), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n469), .A2(new_n754), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n735), .B1(new_n731), .B2(KEYINPUT29), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1180), .B(new_n676), .C1(new_n1181), .C2(new_n468), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1173), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1144), .A2(new_n1175), .A3(new_n957), .A4(new_n1132), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1178), .B2(new_n1174), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n974), .A2(new_n1185), .A3(KEYINPUT117), .A4(new_n1180), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1183), .B(new_n1186), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1136), .A2(new_n1142), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1144), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1136), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n710), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1172), .B1(new_n1188), .B2(new_n1195), .ZN(G378));
  AOI21_X1  g0996(.A(new_n1182), .B1(new_n1147), .B2(new_n1192), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n738), .B1(new_n948), .B2(new_n949), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n308), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1199), .A2(new_n903), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n322), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1200), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n312), .A2(new_n316), .A3(new_n321), .A4(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1201), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1198), .A2(new_n940), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1209), .B1(new_n1198), .B2(new_n940), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1211), .A2(new_n1212), .A3(new_n972), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n959), .A2(new_n903), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n946), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1214), .B1(new_n1138), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1141), .B1(new_n924), .B2(new_n966), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n970), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1198), .A2(new_n940), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1209), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1218), .B1(new_n1221), .B2(new_n1210), .ZN(new_n1222));
  OAI21_X1  g1022(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n710), .B1(new_n1197), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1182), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1194), .A2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n972), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1221), .A2(new_n1218), .A3(new_n1210), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT57), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1224), .A2(new_n1230), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n848), .A2(new_n449), .B1(new_n851), .B2(new_n620), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n791), .A2(G283), .B1(G97), .B2(new_n780), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n444), .B2(new_n786), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n802), .A2(new_n202), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1232), .A2(new_n1234), .A3(new_n999), .A4(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n857), .A2(new_n275), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(new_n1065), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(KEYINPUT120), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(KEYINPUT120), .B2(new_n1238), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT58), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1241), .A2(KEYINPUT58), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1237), .B(new_n227), .C1(G33), .C2(G41), .ZN(new_n1244));
  INV_X1    g1044(.A(G132), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n781), .A2(new_n1245), .B1(new_n786), .B2(new_n850), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n800), .A2(G128), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1247), .B1(new_n296), .B2(new_n797), .C1(new_n851), .C2(new_n1151), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1246), .B(new_n1248), .C1(new_n809), .C2(new_n1154), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT59), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1000), .A2(G159), .ZN(new_n1253));
  AOI211_X1 g1053(.A(G33), .B(G41), .C1(new_n791), .C2(G124), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  AND4_X1   g1055(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n1255), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n762), .B1(G50), .B2(new_n1149), .C1(new_n1256), .C2(new_n846), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1220), .B2(new_n764), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1229), .B2(new_n761), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1231), .A2(new_n1259), .ZN(G375));
  NAND2_X1  g1060(.A1(new_n1185), .A2(new_n761), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G128), .A2(new_n791), .B1(new_n817), .B2(G150), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n781), .B2(new_n1153), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1263), .A2(new_n857), .A3(new_n1235), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n794), .A2(G159), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n851), .A2(new_n1245), .B1(new_n227), .B2(new_n797), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(G137), .B2(new_n800), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1264), .A2(new_n1265), .A3(new_n1267), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n781), .A2(new_n620), .B1(new_n786), .B2(new_n449), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n262), .B(new_n1269), .C1(G303), .C2(new_n791), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n794), .A2(G97), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n798), .A2(new_n564), .B1(new_n1000), .B2(G77), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(G283), .A2(new_n800), .B1(new_n805), .B2(G294), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n846), .B1(new_n1268), .B2(new_n1274), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n763), .B(new_n1275), .C1(new_n203), .C2(new_n870), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(KEYINPUT121), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n941), .B2(new_n765), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT122), .B1(new_n1261), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1261), .A2(KEYINPUT122), .A3(new_n1278), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1059), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1183), .A2(new_n1186), .A3(new_n1283), .A4(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1282), .A2(new_n1285), .ZN(G381));
  OR2_X1    g1086(.A1(G393), .A2(G396), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n873), .A3(new_n1130), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(G387), .A2(new_n1289), .A3(G381), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1191), .A2(new_n1193), .A3(new_n761), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1148), .A2(new_n1171), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1195), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1293), .B1(new_n1294), .B2(new_n1187), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1290), .A2(new_n1295), .A3(new_n1231), .A4(new_n1259), .ZN(G407));
  NOR2_X1   g1096(.A1(new_n683), .A2(new_n684), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1231), .A2(new_n1295), .A3(new_n1259), .ZN(new_n1299));
  OAI211_X1 g1099(.A(G407), .B(G213), .C1(new_n1298), .C2(new_n1299), .ZN(G409));
  AND2_X1   g1100(.A1(G393), .A2(G396), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1288), .A2(new_n1130), .A3(new_n1301), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(G393), .B(new_n828), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(G390), .A2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(G387), .B1(new_n1302), .B2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1130), .B1(new_n1288), .B2(new_n1301), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G390), .A2(new_n1303), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(new_n1307), .A3(new_n1061), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1305), .A2(new_n1308), .ZN(new_n1309));
  OAI211_X1 g1109(.A(G378), .B(new_n1259), .C1(new_n1224), .C2(new_n1230), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1226), .A2(new_n1283), .A3(new_n1229), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1259), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1295), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1310), .A2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(KEYINPUT60), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1315));
  AND2_X1   g1115(.A1(new_n1315), .A2(new_n1284), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1179), .A2(KEYINPUT60), .A3(new_n1182), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n710), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1281), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1320), .A2(new_n1279), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n873), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1282), .B(G384), .C1(new_n1316), .C2(new_n1318), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1314), .A2(new_n1298), .A3(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(KEYINPUT123), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1297), .B1(new_n1310), .B2(new_n1313), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT123), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1327), .A2(new_n1328), .A3(new_n1324), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT62), .B1(new_n1326), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1314), .A2(new_n1298), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1297), .A2(G2897), .ZN(new_n1332));
  XOR2_X1   g1132(.A(new_n1332), .B(KEYINPUT125), .Z(new_n1333));
  AND3_X1   g1133(.A1(new_n1322), .A2(new_n1323), .A3(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1333), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT61), .B1(new_n1331), .B2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1325), .A2(KEYINPUT62), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1309), .B1(new_n1330), .B2(new_n1339), .ZN(new_n1340));
  XOR2_X1   g1140(.A(KEYINPUT124), .B(KEYINPUT63), .Z(new_n1341));
  NAND3_X1  g1141(.A1(new_n1326), .A2(new_n1329), .A3(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1327), .A2(KEYINPUT63), .A3(new_n1324), .ZN(new_n1343));
  AND2_X1   g1143(.A1(new_n1305), .A2(new_n1308), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1342), .A2(new_n1343), .A3(new_n1337), .A4(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1340), .A2(new_n1345), .ZN(G405));
  INV_X1    g1146(.A(KEYINPUT126), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1324), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(KEYINPUT127), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT127), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1324), .A2(new_n1347), .A3(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1349), .A2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1344), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1309), .A2(new_n1349), .A3(new_n1351), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(G375), .A2(G378), .ZN(new_n1356));
  OR2_X1    g1156(.A1(new_n1324), .A2(new_n1347), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1356), .A2(new_n1357), .A3(new_n1299), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1355), .A2(new_n1358), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1358), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1353), .A2(new_n1360), .A3(new_n1354), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1359), .A2(new_n1361), .ZN(G402));
endmodule


