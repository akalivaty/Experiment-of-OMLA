//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G128), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT72), .A3(G119), .ZN(new_n191));
  OAI211_X1 g005(.A(new_n189), .B(new_n191), .C1(G119), .C2(new_n190), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT24), .B(G110), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT73), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n188), .B2(G128), .ZN(new_n196));
  AOI22_X1  g010(.A1(new_n196), .A2(KEYINPUT23), .B1(new_n188), .B2(G128), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n197), .B1(KEYINPUT23), .B2(new_n196), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n194), .B1(new_n198), .B2(G110), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G140), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n203), .A3(KEYINPUT16), .ZN(new_n204));
  OR3_X1    g018(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G146), .ZN(new_n206));
  XNOR2_X1  g020(.A(G125), .B(G140), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n199), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n198), .A2(G110), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n204), .A2(new_n205), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n208), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n206), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n211), .B(new_n214), .C1(new_n193), .C2(new_n192), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G137), .ZN(new_n217));
  INV_X1    g031(.A(G953), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(G221), .A3(G234), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n217), .B(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n216), .A2(new_n221), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT71), .B(G217), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G902), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n227), .B1(G234), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G902), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n231), .A2(KEYINPUT76), .ZN(new_n232));
  INV_X1    g046(.A(new_n224), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT75), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n234), .B1(KEYINPUT74), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(new_n234), .B2(new_n235), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n233), .A2(new_n228), .A3(new_n222), .A4(new_n237), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n223), .A2(G902), .A3(new_n224), .ZN(new_n239));
  INV_X1    g053(.A(new_n236), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n238), .B(new_n229), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n231), .A2(KEYINPUT76), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n232), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n208), .A2(G143), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G146), .ZN(new_n246));
  AND2_X1   g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n244), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n249));
  XNOR2_X1  g063(.A(G143), .B(G146), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT0), .B(G128), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n244), .A2(new_n246), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n253), .A2(new_n255), .A3(KEYINPUT64), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n248), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT11), .ZN(new_n258));
  INV_X1    g072(.A(G134), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(G137), .ZN(new_n260));
  INV_X1    g074(.A(G137), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT11), .A3(G134), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(G137), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n265), .A3(G131), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(G131), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n260), .A2(new_n262), .A3(new_n263), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n257), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT2), .ZN(new_n271));
  INV_X1    g085(.A(G113), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(KEYINPUT68), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(KEYINPUT2), .B2(G113), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n273), .A2(new_n275), .B1(KEYINPUT2), .B2(G113), .ZN(new_n276));
  XNOR2_X1  g090(.A(G116), .B(G119), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n276), .A2(new_n277), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OR2_X1    g095(.A1(new_n264), .A2(G131), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n244), .A2(new_n246), .A3(new_n283), .A4(G128), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n245), .A2(KEYINPUT1), .A3(G146), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n284), .B(new_n285), .C1(G128), .C2(new_n250), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n261), .A2(G134), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n263), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G131), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n282), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n270), .A2(new_n281), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT28), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n270), .A2(new_n281), .A3(new_n293), .A4(new_n290), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n269), .B1(new_n257), .B2(KEYINPUT65), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT65), .ZN(new_n297));
  AOI211_X1 g111(.A(new_n297), .B(new_n248), .C1(new_n252), .C2(new_n256), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n290), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n276), .B(new_n277), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(G237), .A2(G953), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G210), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n304), .B(KEYINPUT27), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT26), .B(G101), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n270), .A2(new_n290), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n300), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n290), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n264), .B(new_n267), .ZN(new_n315));
  INV_X1    g129(.A(new_n248), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n250), .A2(new_n251), .A3(new_n249), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT64), .B1(new_n253), .B2(new_n255), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n315), .B1(new_n319), .B2(new_n297), .ZN(new_n320));
  INV_X1    g134(.A(new_n298), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n314), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT67), .B1(new_n322), .B2(KEYINPUT30), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT67), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n299), .A2(new_n324), .A3(new_n312), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n313), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n291), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(new_n308), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT31), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n310), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n313), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n299), .A2(new_n324), .A3(new_n312), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n324), .B1(new_n299), .B2(new_n312), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n328), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT69), .B1(new_n337), .B2(KEYINPUT31), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT69), .ZN(new_n339));
  AOI211_X1 g153(.A(new_n339), .B(new_n331), .C1(new_n336), .C2(new_n328), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n332), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(G472), .A2(G902), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT32), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n281), .B1(new_n270), .B2(new_n290), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n292), .B2(new_n294), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n307), .A2(KEYINPUT29), .ZN(new_n348));
  AOI21_X1  g162(.A(G902), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n349), .A2(KEYINPUT70), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(KEYINPUT70), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n327), .A2(new_n307), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n336), .A2(new_n352), .B1(new_n302), .B2(new_n307), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n350), .B(new_n351), .C1(new_n353), .C2(KEYINPUT29), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n341), .A2(new_n345), .B1(G472), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n336), .A2(new_n331), .A3(new_n328), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n309), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT31), .B1(new_n326), .B2(new_n329), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n339), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n337), .A2(KEYINPUT69), .A3(KEYINPUT31), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n344), .B1(new_n361), .B2(new_n343), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n243), .B1(new_n355), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT9), .B(G234), .ZN(new_n364));
  OAI21_X1  g178(.A(G221), .B1(new_n364), .B2(G902), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G469), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(new_n228), .ZN(new_n368));
  INV_X1    g182(.A(G104), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(G107), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT3), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT78), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n370), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n369), .A2(G107), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n373), .A2(KEYINPUT78), .ZN(new_n377));
  INV_X1    g191(.A(G107), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G104), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n376), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(G101), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n371), .A2(KEYINPUT3), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n379), .B1(new_n377), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G101), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n370), .A2(new_n372), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n383), .A2(new_n384), .A3(new_n385), .A4(new_n376), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n381), .A2(new_n386), .A3(KEYINPUT4), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n388), .B(G101), .C1(new_n375), .C2(new_n380), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n387), .A2(new_n257), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n379), .A2(new_n376), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G101), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n386), .A2(new_n286), .A3(KEYINPUT10), .A4(new_n392), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT80), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT10), .ZN(new_n396));
  AOI21_X1  g210(.A(G128), .B1(new_n244), .B2(new_n246), .ZN(new_n397));
  INV_X1    g211(.A(new_n285), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT79), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n285), .B(new_n400), .C1(new_n250), .C2(G128), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n399), .A2(new_n284), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n386), .A2(new_n392), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n396), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n394), .A2(new_n395), .A3(new_n315), .A4(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n404), .A2(new_n315), .A3(new_n390), .A4(new_n393), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT80), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n386), .A2(new_n392), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n399), .A2(new_n284), .A3(new_n401), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n286), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n403), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n315), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT12), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n408), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G110), .B(G140), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n218), .A2(G227), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n417), .B(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT77), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n419), .B1(new_n405), .B2(new_n407), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n394), .A2(new_n404), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n269), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n416), .A2(new_n421), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n368), .B1(new_n425), .B2(G469), .ZN(new_n426));
  INV_X1    g240(.A(new_n419), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n408), .A2(new_n415), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n427), .B1(new_n408), .B2(new_n424), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n367), .B(new_n228), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n366), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n387), .A2(new_n300), .A3(new_n389), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n277), .A2(KEYINPUT5), .ZN(new_n433));
  INV_X1    g247(.A(G116), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(G119), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT5), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n272), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n276), .A2(new_n277), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n409), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G122), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n432), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n412), .A2(new_n202), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n202), .B2(new_n257), .ZN(new_n443));
  INV_X1    g257(.A(G224), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT7), .B1(new_n444), .B2(G953), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n445), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n442), .B(new_n447), .C1(new_n202), .C2(new_n257), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n441), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n188), .A2(G116), .ZN(new_n450));
  OAI21_X1  g264(.A(G113), .B1(new_n450), .B2(KEYINPUT5), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n451), .A2(KEYINPUT82), .B1(new_n277), .B2(KEYINPUT5), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(KEYINPUT82), .B2(new_n451), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n278), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n409), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n440), .B(KEYINPUT8), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n403), .A2(new_n438), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n455), .A2(new_n456), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n457), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n403), .B1(new_n278), .B2(new_n453), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT83), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(G902), .B1(new_n449), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n432), .A2(new_n439), .ZN(new_n465));
  INV_X1    g279(.A(new_n440), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(KEYINPUT6), .A3(new_n441), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n444), .A2(G953), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT81), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n443), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n465), .A2(new_n472), .A3(new_n466), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n468), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n464), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(G210), .B1(G237), .B2(G902), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT84), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n464), .A2(new_n474), .A3(new_n476), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G214), .B1(G237), .B2(G902), .ZN(new_n482));
  INV_X1    g296(.A(new_n480), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT84), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT87), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n303), .A2(G143), .A3(G214), .ZN(new_n487));
  AOI21_X1  g301(.A(G143), .B1(new_n303), .B2(G214), .ZN(new_n488));
  OAI211_X1 g302(.A(KEYINPUT17), .B(G131), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n213), .A2(new_n489), .A3(new_n206), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT86), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n488), .ZN(new_n493));
  INV_X1    g307(.A(G131), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n303), .A2(G143), .A3(G214), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G131), .B1(new_n487), .B2(new_n488), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n213), .A2(new_n489), .A3(KEYINPUT86), .A4(new_n206), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n492), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n207), .B(new_n208), .ZN(new_n502));
  OAI211_X1 g316(.A(KEYINPUT18), .B(G131), .C1(new_n487), .C2(new_n488), .ZN(new_n503));
  NAND2_X1  g317(.A1(KEYINPUT18), .A2(G131), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n493), .A2(new_n495), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G113), .B(G122), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(G104), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n509), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT19), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n207), .B(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n206), .B1(new_n514), .B2(G146), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT85), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n496), .B2(new_n497), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n496), .A2(new_n497), .A3(new_n516), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n512), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n511), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(G475), .A2(G902), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n486), .B(KEYINPUT20), .C1(new_n522), .C2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n509), .B1(new_n501), .B2(new_n506), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n526), .A2(new_n520), .A3(new_n524), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT20), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT87), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n524), .A2(KEYINPUT88), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n524), .A2(KEYINPUT88), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT89), .B1(new_n522), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n526), .A2(new_n520), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT89), .ZN(new_n535));
  INV_X1    g349(.A(new_n532), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n525), .A2(new_n529), .A3(new_n533), .A4(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n507), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n509), .A2(KEYINPUT90), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(G902), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n539), .B2(new_n541), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G475), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT13), .B1(new_n190), .B2(G143), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(new_n259), .ZN(new_n546));
  XNOR2_X1  g360(.A(G128), .B(G143), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G122), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G116), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT91), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n434), .A2(G122), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n551), .A2(new_n378), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n378), .B1(new_n551), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n548), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT91), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n550), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n552), .B(KEYINPUT14), .ZN(new_n558));
  OAI21_X1  g372(.A(G107), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n551), .A2(new_n378), .A3(new_n552), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n547), .B(new_n259), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n227), .A2(G953), .A3(new_n364), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n555), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n563), .B1(new_n555), .B2(new_n562), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n228), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G478), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n566), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n564), .ZN(new_n572));
  INV_X1    g386(.A(new_n569), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n228), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n218), .A2(G952), .ZN(new_n576));
  NAND2_X1  g390(.A1(G234), .A2(G237), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(G902), .A3(G953), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT21), .B(G898), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n575), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n538), .A2(new_n544), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT92), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT92), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n538), .A2(new_n587), .A3(new_n584), .A4(new_n544), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n485), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n363), .A2(new_n431), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  OAI21_X1  g405(.A(G472), .B1(new_n361), .B2(G902), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n341), .A2(new_n342), .ZN(new_n593));
  INV_X1    g407(.A(new_n243), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n592), .A2(new_n431), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n538), .A2(new_n544), .ZN(new_n596));
  AND2_X1   g410(.A1(KEYINPUT93), .A2(KEYINPUT33), .ZN(new_n597));
  NOR2_X1   g411(.A1(KEYINPUT93), .A2(KEYINPUT33), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n572), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n568), .A2(G902), .ZN(new_n601));
  INV_X1    g415(.A(new_n572), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n600), .B(new_n601), .C1(new_n602), .C2(new_n597), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n567), .A2(new_n568), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n596), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n482), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n478), .B2(new_n480), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NOR4_X1   g423(.A1(new_n595), .A2(new_n583), .A3(new_n606), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT34), .B(G104), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  NAND2_X1  g426(.A1(new_n527), .A2(new_n528), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n525), .A2(new_n529), .A3(new_n613), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n543), .A2(G475), .B1(new_n570), .B2(new_n574), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n608), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n595), .A2(new_n583), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT35), .B(G107), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G9));
  OR3_X1    g433(.A1(new_n216), .A2(KEYINPUT36), .A3(new_n221), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n216), .B1(KEYINPUT36), .B2(new_n221), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(new_n230), .A3(new_n621), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n622), .A2(KEYINPUT94), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(KEYINPUT94), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n241), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n589), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n592), .A2(new_n593), .ZN(new_n627));
  INV_X1    g441(.A(new_n368), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n422), .A2(new_n424), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n408), .A2(new_n415), .ZN(new_n630));
  OAI211_X1 g444(.A(G469), .B(new_n629), .C1(new_n630), .C2(new_n420), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n430), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n365), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT37), .B(G110), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G12));
  NAND2_X1  g451(.A1(new_n355), .A2(new_n362), .ZN(new_n638));
  AND4_X1   g452(.A1(new_n365), .A2(new_n632), .A3(new_n608), .A4(new_n625), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n578), .B(KEYINPUT96), .Z(new_n641));
  INV_X1    g455(.A(G900), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT95), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n642), .A2(KEYINPUT95), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n581), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n615), .A2(new_n614), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT97), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n640), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n341), .A2(new_n345), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n308), .B1(new_n336), .B2(new_n291), .ZN(new_n653));
  INV_X1    g467(.A(new_n352), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n228), .B1(new_n654), .B2(new_n346), .ZN(new_n655));
  OAI21_X1  g469(.A(G472), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n362), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n481), .A2(new_n484), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT38), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n596), .A2(new_n575), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT38), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n481), .A2(new_n663), .A3(new_n484), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n625), .A2(new_n607), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n660), .A2(new_n662), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n651), .B1(new_n658), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n646), .B(KEYINPUT39), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n431), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT40), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n660), .A2(new_n664), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n661), .A2(new_n607), .A3(new_n625), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n672), .A2(KEYINPUT98), .A3(new_n657), .A4(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n667), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  NAND3_X1  g490(.A1(new_n596), .A2(new_n605), .A3(new_n646), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n640), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G146), .ZN(G48));
  NOR2_X1   g494(.A1(new_n606), .A2(new_n583), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n408), .A2(new_n424), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n682), .A2(new_n419), .B1(new_n422), .B2(new_n415), .ZN(new_n683));
  OAI21_X1  g497(.A(G469), .B1(new_n683), .B2(G902), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n608), .A2(new_n684), .A3(new_n365), .A4(new_n430), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n638), .A2(new_n594), .A3(new_n681), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  INV_X1    g503(.A(new_n583), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n684), .A2(new_n365), .A3(new_n430), .A4(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n616), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n363), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G116), .ZN(G18));
  INV_X1    g508(.A(KEYINPUT99), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT32), .B1(new_n341), .B2(new_n342), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n350), .A2(new_n351), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n336), .A2(new_n352), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n302), .A2(new_n307), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT29), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n345), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n701), .B1(new_n361), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n625), .B1(new_n696), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n586), .A2(new_n588), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n686), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n695), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n685), .B1(new_n588), .B2(new_n586), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(KEYINPUT99), .A3(new_n638), .A4(new_n625), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  OR2_X1    g525(.A1(new_n347), .A2(new_n307), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n358), .A2(new_n356), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n342), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT100), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n713), .A2(KEYINPUT100), .A3(new_n342), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(G472), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n341), .B2(new_n228), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n608), .A2(new_n596), .A3(new_n575), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n691), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(new_n594), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT101), .B(G122), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G24));
  NAND4_X1  g540(.A1(new_n721), .A2(new_n625), .A3(new_n678), .A4(new_n686), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  INV_X1    g542(.A(KEYINPUT102), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n594), .B1(new_n696), .B2(new_n703), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n607), .B1(new_n481), .B2(new_n484), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n678), .A2(new_n431), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n729), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n431), .A2(new_n731), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n677), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(KEYINPUT102), .A3(new_n363), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT42), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n733), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT103), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n361), .A2(new_n702), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n739), .B1(new_n696), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n362), .A2(new_n652), .A3(KEYINPUT103), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n701), .A3(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(KEYINPUT42), .A3(new_n594), .A4(new_n735), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G131), .ZN(G33));
  NAND3_X1  g560(.A1(new_n638), .A2(new_n594), .A3(new_n648), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n734), .ZN(new_n748));
  XOR2_X1   g562(.A(KEYINPUT104), .B(G134), .Z(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G36));
  OAI211_X1 g564(.A(KEYINPUT45), .B(new_n629), .C1(new_n630), .C2(new_n420), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n408), .A2(new_n424), .A3(new_n427), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n420), .B1(new_n408), .B2(new_n415), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n751), .A2(new_n755), .A3(G469), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n757), .A3(new_n430), .A4(new_n628), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n365), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n757), .B1(new_n756), .B2(new_n628), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n668), .A3(new_n731), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n538), .A2(KEYINPUT105), .A3(new_n544), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT105), .B1(new_n538), .B2(new_n544), .ZN(new_n764));
  INV_X1    g578(.A(new_n605), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n605), .A2(new_n767), .ZN(new_n768));
  OAI22_X1  g582(.A1(new_n766), .A2(new_n767), .B1(new_n596), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n361), .A2(new_n343), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n625), .B1(new_n720), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n627), .A2(KEYINPUT106), .A3(new_n625), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n769), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n762), .B1(new_n775), .B2(KEYINPUT44), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n775), .A2(new_n777), .A3(KEYINPUT44), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n768), .A2(new_n596), .ZN(new_n779));
  OR3_X1    g593(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n779), .B1(new_n780), .B2(KEYINPUT43), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT106), .B1(new_n627), .B2(new_n625), .ZN(new_n782));
  INV_X1    g596(.A(new_n625), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n772), .B(new_n783), .C1(new_n592), .C2(new_n593), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n781), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT107), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n776), .B1(new_n778), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  AND2_X1   g603(.A1(new_n758), .A2(new_n365), .ZN(new_n790));
  INV_X1    g604(.A(new_n760), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n790), .A2(KEYINPUT108), .A3(KEYINPUT47), .A4(new_n791), .ZN(new_n792));
  OR2_X1    g606(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n793));
  NAND2_X1  g607(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n793), .B(new_n794), .C1(new_n759), .C2(new_n760), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n731), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n638), .A2(new_n594), .A3(new_n797), .A4(new_n677), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  NAND3_X1  g614(.A1(new_n594), .A2(new_n365), .A3(new_n482), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT109), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n684), .A2(new_n430), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(KEYINPUT49), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(KEYINPUT49), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  OR4_X1    g620(.A1(new_n657), .A2(new_n806), .A3(new_n672), .A4(new_n780), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n769), .A2(new_n641), .ZN(new_n808));
  INV_X1    g622(.A(new_n803), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n365), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n797), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n721), .A2(new_n625), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n811), .A2(new_n658), .A3(new_n594), .A4(new_n579), .ZN(new_n814));
  INV_X1    g628(.A(new_n596), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n765), .ZN(new_n816));
  OAI22_X1  g630(.A1(new_n812), .A2(new_n813), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n672), .A2(new_n482), .A3(new_n810), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n718), .A2(new_n720), .A3(new_n243), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n808), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n817), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n808), .A2(new_n819), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n797), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n803), .A2(new_n365), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n826), .B1(new_n796), .B2(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n824), .A2(KEYINPUT51), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n830));
  OAI22_X1  g644(.A1(new_n796), .A2(new_n830), .B1(new_n365), .B2(new_n803), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT115), .B1(new_n792), .B2(new_n795), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n826), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT51), .B1(new_n824), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n743), .A2(new_n594), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n808), .A3(new_n811), .ZN(new_n836));
  XOR2_X1   g650(.A(new_n836), .B(KEYINPUT48), .Z(new_n837));
  OAI221_X1 g651(.A(new_n576), .B1(new_n606), .B2(new_n814), .C1(new_n825), .C2(new_n685), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n829), .A2(new_n834), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n589), .A2(new_n431), .ZN(new_n840));
  INV_X1    g654(.A(new_n485), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n681), .A2(new_n841), .ZN(new_n842));
  OAI22_X1  g656(.A1(new_n840), .A2(new_n730), .B1(new_n595), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT111), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n595), .A2(new_n583), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n815), .A2(new_n575), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n485), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n846), .A2(new_n848), .B1(new_n626), .B2(new_n634), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n590), .B(KEYINPUT111), .C1(new_n595), .C2(new_n842), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n845), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT110), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n707), .A2(new_n709), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n724), .A2(new_n693), .A3(new_n687), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n734), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n716), .A2(new_n717), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(new_n592), .A3(new_n625), .A4(new_n678), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n570), .A2(new_n574), .A3(new_n646), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(G475), .B2(new_n543), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n860), .A2(new_n614), .A3(KEYINPUT112), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT112), .B1(new_n860), .B2(new_n614), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n863), .B(new_n625), .C1(new_n696), .C2(new_n703), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n747), .A2(new_n858), .A3(new_n864), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n738), .A2(new_n744), .B1(new_n856), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n854), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(KEYINPUT110), .A3(new_n710), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n851), .A2(new_n855), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(KEYINPUT53), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n638), .B(new_n639), .C1(new_n648), .C2(new_n678), .ZN(new_n871));
  INV_X1    g685(.A(new_n722), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n625), .B1(new_n641), .B2(new_n645), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n657), .A2(new_n431), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n727), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n875), .A2(KEYINPUT113), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT52), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n875), .B(KEYINPUT52), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n877), .B1(new_n878), .B2(new_n876), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n870), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT53), .B1(new_n869), .B2(new_n878), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(KEYINPUT54), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n865), .B2(new_n856), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(new_n850), .A3(new_n845), .A4(new_n849), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n854), .B1(new_n707), .B2(new_n709), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n745), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n885), .B1(new_n887), .B2(KEYINPUT114), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT114), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n886), .A2(new_n745), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n879), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n883), .B1(new_n869), .B2(new_n878), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n839), .A2(new_n882), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(G952), .A2(G953), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT116), .Z(new_n897));
  OAI21_X1  g711(.A(new_n807), .B1(new_n895), .B2(new_n897), .ZN(G75));
  NOR2_X1   g712(.A1(new_n218), .A2(G952), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n228), .B1(new_n891), .B2(new_n892), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(G210), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT117), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n468), .A2(new_n473), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(new_n471), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT55), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT56), .B1(new_n901), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n907), .B1(new_n903), .B2(KEYINPUT56), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n899), .B1(new_n911), .B2(new_n912), .ZN(G51));
  NAND2_X1  g727(.A1(new_n891), .A2(new_n892), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT54), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n916), .A3(new_n894), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n914), .A2(KEYINPUT119), .A3(KEYINPUT54), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n368), .B(KEYINPUT57), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n683), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n756), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n900), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n899), .B1(new_n922), .B2(new_n924), .ZN(G54));
  NAND2_X1  g739(.A1(KEYINPUT58), .A2(G475), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT120), .Z(new_n927));
  AND3_X1   g741(.A1(new_n900), .A2(new_n534), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n534), .B1(new_n900), .B2(new_n927), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n899), .ZN(G60));
  INV_X1    g744(.A(new_n899), .ZN(new_n931));
  NAND2_X1  g745(.A1(G478), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT59), .Z(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n882), .B2(new_n894), .ZN(new_n934));
  MUX2_X1   g748(.A(new_n599), .B(new_n597), .S(new_n572), .Z(new_n935));
  OAI21_X1  g749(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n917), .A2(new_n918), .ZN(new_n937));
  INV_X1    g751(.A(new_n933), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n936), .B1(new_n937), .B2(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT60), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n891), .B2(new_n892), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(new_n620), .A3(new_n621), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n944), .B(new_n931), .C1(new_n225), .C2(new_n943), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G66));
  OAI21_X1  g761(.A(G953), .B1(new_n582), .B2(new_n444), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n851), .A2(new_n855), .A3(new_n868), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT121), .Z(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(KEYINPUT122), .B(new_n948), .C1(new_n951), .C2(G953), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT122), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n950), .A2(new_n953), .A3(new_n218), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n905), .B1(G898), .B2(new_n218), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n952), .A2(new_n956), .A3(new_n954), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(G69));
  AOI21_X1  g774(.A(new_n218), .B1(G227), .B2(G900), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT127), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n761), .A2(new_n668), .A3(new_n872), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n748), .B1(new_n835), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n727), .A2(new_n871), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT124), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n727), .A2(new_n871), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n964), .A2(new_n969), .A3(new_n745), .A4(new_n799), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n777), .B1(new_n775), .B2(KEYINPUT44), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n785), .A2(KEYINPUT107), .A3(new_n786), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n970), .B1(new_n973), .B2(new_n776), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n218), .ZN(new_n975));
  OAI22_X1  g789(.A1(new_n334), .A2(new_n335), .B1(new_n312), .B2(new_n311), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT123), .Z(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(new_n514), .Z(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(G900), .B2(G953), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n727), .A2(new_n871), .A3(new_n967), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n967), .B1(new_n727), .B2(new_n871), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n675), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g799(.A(KEYINPUT62), .B(new_n675), .C1(new_n981), .C2(new_n982), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI211_X1 g801(.A(new_n797), .B(new_n669), .C1(new_n606), .C2(new_n847), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n363), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n799), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(new_n973), .B2(new_n776), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n987), .A2(new_n991), .A3(KEYINPUT125), .ZN(new_n992));
  AOI21_X1  g806(.A(KEYINPUT125), .B1(new_n987), .B2(new_n991), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n218), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n978), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT126), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n980), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n994), .A2(KEYINPUT126), .A3(new_n978), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n962), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT125), .ZN(new_n1000));
  AOI21_X1  g814(.A(KEYINPUT62), .B1(new_n969), .B2(new_n675), .ZN(new_n1001));
  INV_X1    g815(.A(new_n986), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n990), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n788), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1000), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n987), .A2(new_n991), .A3(KEYINPUT125), .ZN(new_n1007));
  AOI21_X1  g821(.A(G953), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n978), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n996), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n980), .ZN(new_n1011));
  AND4_X1   g825(.A1(new_n962), .A2(new_n1010), .A3(new_n998), .A4(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n999), .A2(new_n1012), .ZN(G72));
  NAND2_X1  g827(.A1(new_n880), .A2(new_n881), .ZN(new_n1014));
  INV_X1    g828(.A(new_n653), .ZN(new_n1015));
  NAND2_X1  g829(.A1(G472), .A2(G902), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT63), .Z(new_n1017));
  NAND3_X1  g831(.A1(new_n1015), .A2(new_n698), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1017), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1019), .B1(new_n951), .B2(new_n974), .ZN(new_n1020));
  OAI221_X1 g834(.A(new_n931), .B1(new_n1014), .B2(new_n1018), .C1(new_n1020), .C2(new_n698), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n951), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1015), .B1(new_n1022), .B2(new_n1017), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1021), .A2(new_n1023), .ZN(G57));
endmodule


