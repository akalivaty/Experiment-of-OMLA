//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT85), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT85), .ZN(new_n195));
  NOR2_X1   g009(.A1(G237), .A2(G953), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(G214), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT86), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n199), .A2(KEYINPUT18), .A3(G131), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n193), .A2(new_n197), .A3(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n202), .A2(KEYINPUT86), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(G125), .A2(G140), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(G125), .A2(G140), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n208), .B(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n199), .A2(KEYINPUT18), .A3(G131), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n202), .A2(KEYINPUT86), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n204), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT16), .ZN(new_n215));
  INV_X1    g029(.A(G125), .ZN(new_n216));
  INV_X1    g030(.A(G140), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n215), .B1(new_n218), .B2(new_n205), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n216), .A2(KEYINPUT16), .A3(G140), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n214), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT76), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT16), .B1(new_n206), .B2(new_n207), .ZN(new_n223));
  INV_X1    g037(.A(new_n220), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(G146), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(KEYINPUT76), .B(new_n214), .C1(new_n219), .C2(new_n220), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n193), .A2(new_n197), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT66), .B(G131), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT17), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n234));
  INV_X1    g048(.A(new_n230), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n193), .A3(new_n197), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n231), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n228), .A2(new_n233), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G113), .B(G122), .ZN(new_n239));
  INV_X1    g053(.A(G104), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n239), .B(new_n240), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n213), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(new_n213), .B2(new_n238), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n187), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G475), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n231), .A2(new_n236), .ZN(new_n246));
  OR2_X1    g060(.A1(new_n208), .A2(KEYINPUT19), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n208), .A2(KEYINPUT19), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n246), .B(new_n225), .C1(new_n249), .C2(G146), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n241), .B1(new_n213), .B2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n245), .B(new_n187), .C1(new_n242), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT20), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n213), .A2(new_n250), .ZN(new_n254));
  INV_X1    g068(.A(new_n241), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n213), .A2(new_n238), .A3(new_n241), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n258), .A2(new_n259), .A3(new_n245), .A4(new_n187), .ZN(new_n260));
  AOI221_X4 g074(.A(KEYINPUT88), .B1(G475), .B2(new_n244), .C1(new_n253), .C2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT88), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n253), .A2(new_n260), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n244), .A2(G475), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n189), .A2(G952), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(G234), .B2(G237), .ZN(new_n268));
  XOR2_X1   g082(.A(KEYINPUT73), .B(G902), .Z(new_n269));
  AOI21_X1  g083(.A(new_n189), .B1(G234), .B2(G237), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  XOR2_X1   g086(.A(KEYINPUT21), .B(G898), .Z(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n268), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(G128), .B(G143), .ZN(new_n277));
  INV_X1    g091(.A(G134), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n279), .B(KEYINPUT89), .ZN(new_n280));
  XOR2_X1   g094(.A(G116), .B(G122), .Z(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(G107), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n278), .B1(new_n277), .B2(KEYINPUT13), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n194), .A2(G128), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n283), .B1(KEYINPUT13), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n280), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n277), .B(new_n278), .ZN(new_n287));
  INV_X1    g101(.A(G116), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(KEYINPUT14), .A3(G122), .ZN(new_n289));
  OAI211_X1 g103(.A(G107), .B(new_n289), .C1(new_n281), .C2(KEYINPUT14), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n287), .B(new_n290), .C1(G107), .C2(new_n281), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  XOR2_X1   g106(.A(KEYINPUT9), .B(G234), .Z(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(G217), .A3(new_n189), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n292), .B(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(new_n269), .ZN(new_n297));
  INV_X1    g111(.A(G478), .ZN(new_n298));
  NOR2_X1   g112(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n297), .B(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n266), .A2(new_n276), .A3(new_n305), .ZN(new_n306));
  XOR2_X1   g120(.A(G110), .B(G122), .Z(new_n307));
  INV_X1    g121(.A(G119), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT68), .B1(new_n308), .B2(G116), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT68), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(new_n288), .A3(G119), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n309), .A2(new_n311), .B1(G116), .B2(new_n308), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT2), .B(G113), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(new_n240), .B2(G107), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n316));
  INV_X1    g130(.A(G107), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(G104), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n240), .A2(G107), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n315), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G101), .ZN(new_n322));
  INV_X1    g136(.A(G101), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n315), .A2(new_n318), .A3(new_n323), .A4(new_n319), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT4), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT4), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n314), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT5), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(new_n308), .A3(G116), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n309), .A2(new_n311), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n308), .A2(G116), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g148(.A(G113), .B(new_n331), .C1(new_n334), .C2(new_n330), .ZN(new_n335));
  INV_X1    g149(.A(new_n319), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n240), .A2(G107), .ZN(new_n337));
  OAI21_X1  g151(.A(G101), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n338), .A2(new_n324), .ZN(new_n339));
  INV_X1    g153(.A(new_n313), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n312), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n335), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n307), .B1(new_n329), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n312), .A2(new_n340), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n341), .ZN(new_n347));
  INV_X1    g161(.A(new_n328), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n327), .B1(new_n322), .B2(new_n324), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n307), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n342), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n344), .A2(KEYINPUT6), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT80), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n344), .A2(new_n352), .A3(new_n355), .A4(KEYINPUT6), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n194), .A2(G146), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n214), .A2(G143), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT1), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n358), .A2(new_n359), .A3(new_n360), .A4(G128), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n214), .A2(G143), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(G128), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n194), .A2(G128), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n214), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n361), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n216), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n358), .A2(new_n359), .ZN(new_n369));
  NAND2_X1  g183(.A1(KEYINPUT0), .A2(G128), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n371));
  NOR2_X1   g185(.A1(KEYINPUT0), .A2(G128), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT64), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n369), .A2(new_n370), .A3(new_n371), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT65), .ZN(new_n376));
  XNOR2_X1  g190(.A(G143), .B(G146), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(KEYINPUT0), .A3(G128), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n358), .A2(new_n359), .B1(new_n372), .B2(new_n373), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT65), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n379), .A2(new_n380), .A3(new_n370), .A4(new_n371), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n376), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n368), .B1(new_n382), .B2(new_n216), .ZN(new_n383));
  INV_X1    g197(.A(G224), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(G953), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n385), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n350), .A2(new_n342), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n307), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n389), .A2(KEYINPUT82), .A3(new_n307), .A4(new_n390), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n357), .A2(new_n388), .A3(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n386), .B(new_n387), .C1(KEYINPUT7), .C2(new_n385), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT83), .B(KEYINPUT8), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n307), .B(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n339), .B1(new_n335), .B2(new_n341), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n399), .B1(new_n343), .B2(new_n400), .ZN(new_n401));
  OR3_X1    g215(.A1(new_n383), .A2(KEYINPUT7), .A3(new_n385), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n397), .A2(new_n352), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n396), .A2(new_n187), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(G210), .B1(G237), .B2(G902), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(KEYINPUT84), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n406), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n396), .A2(new_n187), .A3(new_n408), .A4(new_n403), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G214), .B1(G237), .B2(G902), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n306), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G469), .ZN(new_n414));
  INV_X1    g228(.A(new_n269), .ZN(new_n415));
  XNOR2_X1  g229(.A(G110), .B(G140), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n189), .A2(G227), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n416), .B(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n367), .B1(new_n324), .B2(new_n338), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n361), .A2(KEYINPUT78), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT78), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n377), .A2(new_n422), .A3(new_n360), .A4(G128), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n214), .A2(new_n365), .B1(new_n362), .B2(new_n363), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n420), .B1(new_n339), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT11), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n278), .B2(G137), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n278), .A2(G137), .ZN(new_n429));
  INV_X1    g243(.A(G137), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(KEYINPUT11), .A3(G134), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(new_n230), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n428), .A2(new_n431), .A3(new_n434), .A4(new_n429), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n435), .A2(G131), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(KEYINPUT67), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n433), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT12), .B1(new_n426), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n425), .A2(new_n339), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(new_n339), .B2(new_n367), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT12), .ZN(new_n442));
  INV_X1    g256(.A(new_n433), .ZN(new_n443));
  INV_X1    g257(.A(new_n437), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n435), .A2(G131), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n441), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n439), .A2(new_n447), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n376), .A2(new_n378), .A3(new_n381), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n349), .B2(new_n348), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT10), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n424), .B2(new_n361), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n440), .A2(new_n451), .B1(new_n339), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT79), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n450), .A2(new_n453), .A3(new_n454), .A4(new_n438), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n450), .A2(new_n453), .A3(new_n438), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT79), .ZN(new_n457));
  AOI211_X1 g271(.A(new_n419), .B(new_n448), .C1(new_n455), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n455), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n450), .A2(new_n453), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n446), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n418), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n414), .B(new_n415), .C1(new_n458), .C2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n414), .A2(new_n187), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n459), .A2(new_n461), .A3(new_n418), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n448), .B1(new_n455), .B2(new_n457), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n466), .B(G469), .C1(new_n418), .C2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n463), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n308), .A2(G128), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT74), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n308), .A2(G128), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT24), .B(G110), .Z(new_n474));
  INV_X1    g288(.A(KEYINPUT75), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT23), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT23), .ZN(new_n477));
  OAI211_X1 g291(.A(KEYINPUT75), .B(new_n477), .C1(new_n308), .C2(G128), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n470), .A3(new_n478), .ZN(new_n479));
  OAI22_X1  g293(.A1(new_n473), .A2(new_n474), .B1(G110), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n480), .B(new_n225), .C1(G146), .C2(new_n208), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n473), .A2(new_n474), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(G110), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n482), .A2(new_n227), .A3(new_n226), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT22), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(G137), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n481), .A2(new_n484), .A3(new_n488), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n415), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT25), .ZN(new_n493));
  INV_X1    g307(.A(G217), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n494), .B1(new_n415), .B2(G234), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT25), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n490), .A2(new_n496), .A3(new_n415), .A4(new_n491), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n490), .A2(new_n491), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n495), .A2(G902), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n293), .ZN(new_n503));
  OAI21_X1  g317(.A(G221), .B1(new_n503), .B2(G902), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n469), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT32), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n449), .A2(new_n446), .ZN(new_n508));
  INV_X1    g322(.A(new_n429), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n278), .A2(G137), .ZN(new_n510));
  OAI21_X1  g324(.A(G131), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n443), .A2(new_n367), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n507), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n507), .B(new_n512), .C1(new_n438), .C2(new_n382), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n347), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n512), .B1(new_n438), .B2(new_n382), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT69), .ZN(new_n518));
  INV_X1    g332(.A(new_n341), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n518), .B1(new_n519), .B2(new_n345), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n346), .A2(KEYINPUT69), .A3(new_n341), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n525));
  NAND2_X1  g339(.A1(new_n196), .A2(G210), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT26), .B(G101), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n516), .A2(new_n524), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT31), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n520), .A2(new_n521), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n367), .A2(new_n511), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n449), .A2(new_n446), .B1(new_n443), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT28), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT28), .B1(new_n517), .B2(new_n522), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n517), .A2(new_n347), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n529), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n517), .A2(KEYINPUT30), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n514), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n523), .B1(new_n544), .B2(new_n347), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT31), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n546), .A3(new_n530), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n532), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(G472), .A2(G902), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT71), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n548), .A2(KEYINPUT72), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT72), .B1(new_n548), .B2(new_n551), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n506), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n541), .A2(new_n530), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n545), .A2(new_n529), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT29), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n517), .A2(new_n522), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n539), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n530), .A2(KEYINPUT29), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n415), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G472), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n548), .A2(KEYINPUT32), .A3(new_n551), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n554), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n413), .A2(new_n505), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(G101), .ZN(G3));
  INV_X1    g381(.A(KEYINPUT72), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n546), .B1(new_n545), .B2(new_n530), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n314), .B1(new_n543), .B2(new_n514), .ZN(new_n570));
  NOR4_X1   g384(.A1(new_n570), .A2(KEYINPUT31), .A3(new_n523), .A4(new_n529), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n530), .B1(new_n539), .B2(new_n540), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n568), .B1(new_n573), .B2(new_n550), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n548), .A2(KEYINPUT72), .A3(new_n551), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT91), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n548), .A2(new_n415), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n577), .B1(new_n578), .B2(G472), .ZN(new_n579));
  INV_X1    g393(.A(G472), .ZN(new_n580));
  AOI211_X1 g394(.A(KEYINPUT91), .B(new_n580), .C1(new_n548), .C2(new_n415), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n576), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n469), .A2(new_n502), .A3(new_n504), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT92), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n578), .A2(G472), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT91), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n578), .A2(new_n577), .A3(G472), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n588), .A2(new_n505), .A3(new_n589), .A4(new_n576), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n591), .B(KEYINPUT93), .Z(new_n592));
  NOR2_X1   g406(.A1(new_n405), .A2(KEYINPUT94), .ZN(new_n593));
  INV_X1    g407(.A(new_n405), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT94), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n404), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n596), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n396), .A2(new_n187), .A3(new_n403), .A4(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n593), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n600), .A2(new_n412), .A3(new_n275), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n297), .A2(new_n298), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n294), .B2(KEYINPUT95), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n296), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n296), .A2(new_n605), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n415), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n603), .B1(new_n608), .B2(G478), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n261), .B2(new_n265), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT96), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n592), .A2(new_n601), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  NAND2_X1  g429(.A1(new_n263), .A2(KEYINPUT97), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n253), .A2(new_n260), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n616), .A2(new_n304), .A3(new_n264), .A4(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n592), .A2(new_n601), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT35), .B(G107), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  INV_X1    g437(.A(new_n582), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n489), .A2(KEYINPUT36), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n485), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n500), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n498), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n469), .A2(new_n504), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n413), .A2(new_n624), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n631), .B(KEYINPUT37), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G110), .ZN(G12));
  XNOR2_X1  g447(.A(new_n268), .B(KEYINPUT99), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT98), .B(G900), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n271), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT100), .B1(new_n619), .B2(new_n637), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n253), .A2(new_n260), .A3(new_n617), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n617), .B1(new_n253), .B2(new_n260), .ZN(new_n640));
  INV_X1    g454(.A(new_n264), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n643));
  INV_X1    g457(.A(new_n637), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n642), .A2(new_n643), .A3(new_n304), .A4(new_n644), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n629), .B1(new_n554), .B2(new_n564), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n597), .A2(new_n599), .ZN(new_n648));
  INV_X1    g462(.A(new_n593), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n412), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n646), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n653));
  INV_X1    g467(.A(new_n628), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n469), .A2(new_n504), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n637), .B(KEYINPUT101), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT39), .Z(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n655), .A2(KEYINPUT102), .A3(new_n657), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT40), .B1(new_n660), .B2(new_n661), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n654), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n410), .B(KEYINPUT38), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n266), .A2(new_n305), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n545), .A2(new_n529), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n558), .A2(new_n529), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n187), .B1(new_n671), .B2(new_n523), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n554), .A2(new_n563), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n668), .A2(new_n411), .A3(new_n669), .A4(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n653), .B1(new_n666), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n662), .B(new_n663), .ZN(new_n677));
  INV_X1    g491(.A(new_n675), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n677), .A2(new_n678), .A3(KEYINPUT103), .A4(new_n654), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n194), .ZN(G45));
  OAI211_X1 g495(.A(new_n609), .B(new_n644), .C1(new_n261), .C2(new_n265), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n647), .A2(new_n650), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  OAI21_X1  g499(.A(new_n415), .B1(new_n458), .B2(new_n462), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(KEYINPUT104), .A3(G469), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n459), .A2(new_n461), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n419), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n467), .A2(new_n418), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n269), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(KEYINPUT104), .A2(G469), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n687), .A2(new_n693), .A3(new_n504), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n687), .A2(new_n693), .A3(KEYINPUT105), .A4(new_n504), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n498), .A2(new_n501), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n554), .B2(new_n564), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n612), .A2(new_n601), .A3(new_n698), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND4_X1  g517(.A1(new_n601), .A2(new_n698), .A3(new_n620), .A4(new_n700), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  NOR3_X1   g519(.A1(new_n600), .A2(new_n694), .A3(new_n412), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n306), .A2(new_n654), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n565), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  AND3_X1   g523(.A1(new_n498), .A2(KEYINPUT107), .A3(new_n501), .ZN(new_n710));
  AOI21_X1  g524(.A(KEYINPUT107), .B1(new_n498), .B2(new_n501), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n559), .A2(new_n529), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n532), .A2(new_n713), .A3(new_n547), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n551), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT106), .B1(new_n578), .B2(G472), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n717), .B(new_n580), .C1(new_n548), .C2(new_n415), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n712), .B(new_n715), .C1(new_n716), .C2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n720), .A2(new_n601), .A3(new_n698), .A4(new_n669), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  OAI211_X1 g536(.A(new_n628), .B(new_n715), .C1(new_n716), .C2(new_n718), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n682), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n706), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n407), .A2(new_n411), .A3(new_n409), .ZN(new_n728));
  INV_X1    g542(.A(new_n504), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n464), .B1(new_n691), .B2(new_n414), .ZN(new_n730));
  INV_X1    g544(.A(new_n467), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(KEYINPUT108), .A3(new_n419), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n733), .B1(new_n467), .B2(new_n418), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n732), .A2(new_n734), .A3(G469), .A4(new_n466), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n729), .B1(new_n730), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n728), .A2(new_n683), .A3(new_n736), .A4(KEYINPUT42), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n506), .B1(new_n573), .B2(new_n550), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n564), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n712), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n727), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n735), .A2(new_n463), .A3(new_n465), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n504), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n407), .A2(new_n411), .A3(new_n409), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n682), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n710), .A2(new_n711), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(new_n564), .B2(new_n738), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n745), .A2(new_n747), .A3(KEYINPUT109), .A4(KEYINPUT42), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n743), .A2(new_n744), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n700), .A2(new_n749), .A3(new_n683), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n741), .A2(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT110), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  AOI21_X1  g568(.A(KEYINPUT32), .B1(new_n574), .B2(new_n575), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n562), .A2(new_n563), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n502), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n728), .A2(new_n736), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n760), .A3(new_n646), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n646), .A2(new_n700), .A3(new_n749), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT111), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NOR2_X1   g579(.A1(new_n624), .A2(new_n654), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n266), .A2(new_n767), .A3(new_n609), .ZN(new_n768));
  INV_X1    g582(.A(new_n609), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n266), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(KEYINPUT112), .B1(new_n261), .B2(new_n265), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n766), .B(new_n768), .C1(new_n767), .C2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n776));
  OR3_X1    g590(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n732), .A2(new_n734), .A3(KEYINPUT45), .A4(new_n466), .ZN(new_n778));
  INV_X1    g592(.A(new_n466), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n779), .B1(new_n419), .B2(new_n731), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n778), .B(G469), .C1(new_n780), .C2(KEYINPUT45), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n465), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT46), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n781), .A2(KEYINPUT46), .A3(new_n465), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n463), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n504), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n657), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n744), .B1(new_n774), .B2(new_n776), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n775), .B1(new_n774), .B2(new_n776), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n777), .A2(new_n790), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n787), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n786), .A2(KEYINPUT47), .A3(new_n504), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n744), .A2(new_n502), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n565), .A2(new_n682), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G140), .ZN(G42));
  INV_X1    g616(.A(new_n773), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n687), .A2(new_n693), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n804), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n808), .A2(new_n674), .A3(new_n729), .A4(new_n746), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n807), .A2(new_n809), .A3(new_n411), .A4(new_n667), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n811));
  INV_X1    g625(.A(new_n723), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n745), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n565), .A2(new_n642), .A3(new_n630), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n305), .A3(new_n644), .A4(new_n728), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n760), .B1(new_n759), .B2(new_n646), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n760), .A2(new_n646), .A3(new_n700), .A4(new_n749), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n813), .B(new_n815), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n263), .A2(new_n264), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT88), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n263), .A2(new_n262), .A3(new_n264), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n304), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n610), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n412), .B1(new_n407), .B2(new_n409), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n823), .A2(new_n824), .A3(new_n276), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n584), .A2(new_n825), .A3(new_n590), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n566), .A3(new_n631), .A4(new_n708), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n701), .A2(new_n721), .A3(new_n704), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n818), .A2(new_n752), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n650), .A2(new_n565), .A3(new_n630), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n830), .A2(new_n646), .B1(new_n706), .B2(new_n724), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n650), .A2(new_n669), .A3(new_n644), .A4(new_n736), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n674), .A2(new_n654), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n831), .A2(new_n834), .A3(KEYINPUT52), .A4(new_n684), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n725), .A2(new_n651), .A3(new_n684), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n832), .A2(new_n833), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT53), .B1(new_n829), .B2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n827), .A2(new_n752), .A3(new_n828), .ZN(new_n842));
  INV_X1    g656(.A(new_n818), .ZN(new_n843));
  AND4_X1   g657(.A1(KEYINPUT53), .A2(new_n842), .A3(new_n840), .A4(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n811), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(new_n840), .A3(new_n843), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n829), .A2(KEYINPUT53), .A3(new_n840), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n849), .A3(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n634), .B(new_n768), .C1(new_n773), .C2(new_n767), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n719), .ZN(new_n853));
  INV_X1    g667(.A(new_n694), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n410), .A2(KEYINPUT38), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n410), .A2(KEYINPUT38), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n412), .B(new_n854), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT114), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n667), .A2(new_n859), .A3(new_n412), .A4(new_n854), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n853), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT50), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n853), .A2(new_n858), .A3(KEYINPUT50), .A4(new_n860), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n805), .A2(new_n504), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n728), .B(new_n853), .C1(new_n798), .C2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n744), .A2(new_n694), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n268), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n869), .A2(new_n674), .A3(new_n699), .A4(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n266), .A3(new_n769), .ZN(new_n872));
  OR3_X1    g686(.A1(new_n852), .A2(new_n723), .A3(new_n869), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n865), .A2(new_n867), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n875), .A2(KEYINPUT51), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n874), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(KEYINPUT51), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n267), .B1(new_n853), .B2(new_n706), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n851), .A2(new_n877), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n871), .A2(new_n612), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n852), .A2(new_n740), .A3(new_n869), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT48), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(G952), .A2(G953), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n810), .B1(new_n884), .B2(new_n885), .ZN(G75));
  NOR2_X1   g700(.A1(new_n189), .A2(G952), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n415), .B1(new_n848), .B2(new_n849), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT56), .B1(new_n889), .B2(new_n594), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n357), .A2(new_n395), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(new_n388), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT116), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT55), .Z(new_n894));
  OAI21_X1  g708(.A(new_n888), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n848), .A2(new_n849), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT117), .B1(new_n896), .B2(new_n269), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n898));
  AOI211_X1 g712(.A(new_n898), .B(new_n415), .C1(new_n848), .C2(new_n849), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT56), .B1(new_n900), .B2(new_n594), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n895), .B1(new_n901), .B2(new_n894), .ZN(G51));
  INV_X1    g716(.A(new_n781), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n464), .B(KEYINPUT57), .Z(new_n905));
  OAI22_X1  g719(.A1(new_n851), .A2(new_n905), .B1(new_n462), .B2(new_n458), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n887), .B1(new_n904), .B2(new_n906), .ZN(G54));
  NAND2_X1  g721(.A1(new_n896), .A2(new_n269), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n898), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n889), .A2(KEYINPUT117), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n909), .A2(KEYINPUT58), .A3(G475), .A4(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n258), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n900), .A2(KEYINPUT58), .A3(G475), .A4(new_n258), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n888), .ZN(G60));
  NAND2_X1  g729(.A1(new_n606), .A2(new_n607), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT118), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT59), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n845), .A2(new_n850), .A3(new_n918), .A4(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n921), .A2(KEYINPUT119), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n921), .A2(KEYINPUT119), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n888), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n845), .A2(new_n850), .A3(new_n920), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n925), .A2(new_n926), .A3(new_n917), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n926), .B1(new_n925), .B2(new_n917), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n924), .A2(new_n929), .ZN(G63));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT61), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT123), .Z(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT60), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n896), .A2(new_n626), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n936), .B1(new_n848), .B2(new_n849), .ZN(new_n941));
  OAI221_X1 g755(.A(new_n888), .B1(new_n931), .B2(KEYINPUT61), .C1(new_n941), .C2(new_n499), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n934), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n938), .B(KEYINPUT121), .ZN(new_n944));
  INV_X1    g758(.A(new_n942), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n933), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n943), .A2(new_n946), .ZN(G66));
  OAI21_X1  g761(.A(G953), .B1(new_n274), .B2(new_n384), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n827), .A2(new_n828), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(G953), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n891), .B1(G898), .B2(new_n189), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G69));
  XOR2_X1   g766(.A(new_n544), .B(new_n249), .Z(new_n953));
  XOR2_X1   g767(.A(KEYINPUT125), .B(G900), .Z(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n956), .B(KEYINPUT124), .Z(new_n958));
  NAND3_X1  g772(.A1(new_n777), .A2(new_n791), .A3(new_n792), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n747), .A2(new_n650), .A3(new_n669), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n764), .B1(new_n961), .B2(new_n789), .ZN(new_n962));
  INV_X1    g776(.A(new_n801), .ZN(new_n963));
  OR3_X1    g777(.A1(new_n963), .A2(new_n752), .A3(new_n837), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n189), .B(new_n953), .C1(new_n962), .C2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT62), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n680), .B2(new_n837), .ZN(new_n967));
  INV_X1    g781(.A(new_n837), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n676), .A2(new_n679), .A3(KEYINPUT62), .A4(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n963), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n662), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n971), .A2(new_n700), .A3(new_n728), .A4(new_n823), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n793), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(G953), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n958), .B(new_n965), .C1(new_n974), .C2(new_n953), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n189), .A2(G900), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n957), .B1(new_n975), .B2(new_n976), .ZN(G72));
  XNOR2_X1  g791(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n580), .A2(new_n187), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n978), .B(new_n979), .Z(new_n980));
  INV_X1    g794(.A(new_n556), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n981), .A2(new_n670), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n896), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT127), .Z(new_n984));
  NAND2_X1  g798(.A1(new_n967), .A2(new_n969), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n985), .A2(new_n801), .A3(new_n949), .A4(new_n973), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n980), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n887), .B1(new_n987), .B2(new_n670), .ZN(new_n988));
  NOR4_X1   g802(.A1(new_n962), .A2(new_n827), .A3(new_n964), .A4(new_n828), .ZN(new_n989));
  INV_X1    g803(.A(new_n980), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n981), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n984), .A2(new_n988), .A3(new_n991), .ZN(G57));
endmodule


