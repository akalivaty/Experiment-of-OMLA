//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1193, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1256, new_n1257,
    new_n1258, new_n1259;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G107), .A2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n212), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n202), .C2(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(G58), .A2(G232), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n211), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n211), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n228), .A2(new_n209), .A3(new_n229), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n224), .A2(new_n227), .A3(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G264), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n218), .ZN(new_n241));
  INV_X1    g0041(.A(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT66), .B(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G351));
  NAND2_X1  g0048(.A1(G33), .A2(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n250), .B1(G232), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G226), .A2(G1698), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n229), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT68), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n229), .B1(KEYINPUT67), .B2(new_n256), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT67), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G33), .A3(G41), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n256), .A2(KEYINPUT67), .ZN(new_n268));
  AND4_X1   g0068(.A1(new_n263), .A2(new_n268), .A3(new_n266), .A4(new_n255), .ZN(new_n269));
  OAI211_X1 g0069(.A(G274), .B(new_n262), .C1(new_n267), .C2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n262), .ZN(new_n271));
  OAI211_X1 g0071(.A(G238), .B(new_n271), .C1(new_n267), .C2(new_n269), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n259), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT13), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT13), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n259), .A2(new_n270), .A3(new_n272), .A4(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(G179), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT70), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n274), .A2(new_n279), .A3(new_n276), .ZN(new_n280));
  OR3_X1    g0080(.A1(new_n273), .A2(new_n279), .A3(KEYINPUT13), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(new_n281), .A3(G169), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT14), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT14), .A4(G169), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n278), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n229), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(G1), .B2(new_n209), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G50), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n209), .A2(G33), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(new_n202), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n214), .A2(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n288), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT11), .ZN(new_n299));
  AOI22_X1  g0099(.A1(G68), .A2(new_n291), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n298), .A2(new_n299), .ZN(new_n301));
  INV_X1    g0101(.A(G13), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G1), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT71), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT12), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(new_n305), .B2(new_n306), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n300), .A2(new_n301), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n286), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n280), .A2(new_n281), .A3(G200), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n273), .B2(KEYINPUT13), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n310), .B1(new_n315), .B2(new_n276), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT72), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n313), .A2(KEYINPUT72), .A3(new_n316), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n268), .A2(new_n266), .A3(new_n255), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT68), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n264), .A2(new_n263), .A3(new_n266), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n262), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G244), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n251), .A2(G232), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n250), .B(new_n327), .C1(new_n215), .C2(new_n251), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n328), .B(new_n258), .C1(G107), .C2(new_n250), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n326), .A2(new_n270), .A3(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n330), .A2(G200), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n314), .ZN(new_n332));
  XOR2_X1   g0132(.A(KEYINPUT8), .B(G58), .Z(new_n333));
  AOI22_X1  g0133(.A1(new_n333), .A2(new_n292), .B1(G20), .B2(G77), .ZN(new_n334));
  XOR2_X1   g0134(.A(KEYINPUT15), .B(G87), .Z(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n334), .B1(new_n294), .B2(new_n336), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n337), .A2(new_n288), .B1(G77), .B2(new_n291), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(G77), .B2(new_n339), .ZN(new_n340));
  OR3_X1    g0140(.A1(new_n331), .A2(new_n332), .A3(new_n340), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n312), .A2(new_n321), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  NOR2_X1   g0143(.A1(KEYINPUT3), .A2(G33), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(G223), .B2(G1698), .ZN(new_n346));
  INV_X1    g0146(.A(G222), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(G1698), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n348), .B(new_n258), .C1(G77), .C2(new_n250), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n325), .A2(G226), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n270), .A3(new_n350), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n351), .A2(G179), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n209), .B1(new_n201), .B2(new_n203), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(G150), .B2(new_n292), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n333), .A2(KEYINPUT69), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT8), .B(G58), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT69), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n354), .B1(new_n359), .B2(new_n294), .ZN(new_n360));
  INV_X1    g0160(.A(new_n339), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n360), .A2(new_n288), .B1(new_n218), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n218), .B2(new_n290), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n351), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n352), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n351), .A2(G200), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n363), .A2(KEYINPUT9), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n363), .A2(KEYINPUT9), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n368), .B1(new_n314), .B2(new_n351), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n371), .A2(KEYINPUT10), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(KEYINPUT10), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT17), .ZN(new_n375));
  OAI211_X1 g0175(.A(G232), .B(new_n271), .C1(new_n267), .C2(new_n269), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n219), .A2(G1698), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n377), .B1(G223), .B2(G1698), .C1(new_n343), .C2(new_n344), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G33), .ZN(new_n380));
  INV_X1    g0180(.A(G87), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n258), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n270), .A2(new_n376), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT74), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT74), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n270), .A2(new_n376), .A3(new_n383), .A4(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(G200), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n384), .A2(G190), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n345), .B2(new_n209), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NOR4_X1   g0192(.A1(new_n343), .A2(new_n344), .A3(new_n392), .A4(G20), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n292), .A2(G159), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n242), .A2(new_n214), .ZN(new_n396));
  OAI21_X1  g0196(.A(G20), .B1(new_n396), .B2(new_n203), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n394), .A2(KEYINPUT16), .A3(new_n395), .A4(new_n397), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n288), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n355), .A2(new_n358), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n291), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n404), .B(KEYINPUT73), .C1(new_n339), .C2(new_n403), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT73), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n403), .A2(new_n339), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n290), .B1(new_n358), .B2(new_n355), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n402), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n375), .B1(new_n390), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n411), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n413), .B(KEYINPUT17), .C1(new_n388), .C2(new_n389), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n385), .A2(new_n387), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n364), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n384), .A2(G179), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n417), .A2(KEYINPUT18), .A3(new_n411), .A4(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT75), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n417), .A2(new_n411), .A3(new_n419), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n423), .A2(new_n421), .A3(new_n424), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n415), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n330), .A2(new_n364), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n340), .B(new_n429), .C1(G179), .C2(new_n330), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n342), .A2(new_n374), .A3(new_n428), .A4(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT83), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n208), .A2(G45), .ZN(new_n434));
  OR2_X1    g0234(.A1(KEYINPUT5), .A2(G41), .ZN(new_n435));
  NAND2_X1  g0235(.A1(KEYINPUT5), .A2(G41), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(G274), .B(new_n437), .C1(new_n267), .C2(new_n269), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT76), .ZN(new_n439));
  INV_X1    g0239(.A(G274), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(new_n323), .B2(new_n324), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT76), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(new_n437), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n437), .B1(new_n323), .B2(new_n324), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n250), .B1(G257), .B2(new_n251), .ZN(new_n446));
  NOR2_X1   g0246(.A1(G250), .A2(G1698), .ZN(new_n447));
  INV_X1    g0247(.A(G294), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n446), .A2(new_n447), .B1(new_n380), .B2(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(G264), .A2(new_n445), .B1(new_n449), .B2(new_n258), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n444), .A2(G179), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n364), .B1(new_n444), .B2(new_n450), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n433), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n444), .A2(new_n450), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G169), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(KEYINPUT83), .A3(new_n451), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n250), .A2(new_n209), .A3(G87), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT22), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT22), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n250), .A2(new_n461), .A3(new_n209), .A4(G87), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT24), .ZN(new_n464));
  INV_X1    g0264(.A(G107), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT81), .B1(new_n465), .B2(G20), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT23), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G116), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n294), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n466), .A2(KEYINPUT23), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n463), .A2(new_n464), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n464), .B1(new_n463), .B2(new_n472), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n288), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n208), .A2(G33), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n339), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(new_n288), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(new_n465), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n303), .A2(G20), .A3(new_n465), .ZN(new_n482));
  XOR2_X1   g0282(.A(new_n482), .B(KEYINPUT25), .Z(new_n483));
  NAND3_X1  g0283(.A1(new_n475), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT82), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT82), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n475), .A2(new_n486), .A3(new_n481), .A4(new_n483), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n455), .A2(G200), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n444), .A2(G190), .A3(new_n450), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n484), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n458), .A2(new_n488), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n250), .A2(KEYINPUT4), .A3(G244), .A4(new_n251), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G283), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n345), .A2(new_n220), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n494), .B(new_n495), .C1(new_n496), .C2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n250), .A2(G250), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n251), .B1(new_n498), .B2(KEYINPUT4), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n258), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n445), .A2(G257), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n444), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G200), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n465), .A2(KEYINPUT6), .A3(G97), .ZN(new_n504));
  XOR2_X1   g0304(.A(G97), .B(G107), .Z(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(KEYINPUT6), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(G20), .B1(G77), .B2(new_n292), .ZN(new_n507));
  OAI21_X1  g0307(.A(G107), .B1(new_n391), .B2(new_n393), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n289), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G97), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n479), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n339), .A2(G97), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n503), .B(new_n513), .C1(new_n314), .C2(new_n502), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n502), .A2(new_n364), .ZN(new_n515));
  INV_X1    g0315(.A(new_n513), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n439), .A2(new_n443), .B1(G257), .B2(new_n445), .ZN(new_n517));
  INV_X1    g0317(.A(G179), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(new_n500), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n251), .A2(G257), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G264), .A2(G1698), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n250), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g0324(.A(KEYINPUT79), .B(G303), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n524), .B(new_n258), .C1(new_n250), .C2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(G270), .B2(new_n445), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n444), .A2(new_n528), .A3(G190), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n361), .A2(new_n469), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n289), .A2(G116), .A3(new_n339), .A4(new_n476), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n287), .A2(new_n229), .B1(G20), .B2(new_n469), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n495), .B(new_n209), .C1(G33), .C2(new_n510), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n532), .A2(KEYINPUT20), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT20), .B1(new_n532), .B2(new_n533), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n530), .B(new_n531), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n536), .A2(KEYINPUT80), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n536), .A2(KEYINPUT80), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n445), .A2(G270), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n526), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(new_n443), .B2(new_n439), .ZN(new_n542));
  INV_X1    g0342(.A(G200), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n529), .B(new_n539), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT21), .ZN(new_n545));
  OAI21_X1  g0345(.A(G169), .B1(new_n537), .B2(new_n538), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(new_n542), .ZN(new_n547));
  XNOR2_X1  g0347(.A(new_n536), .B(KEYINPUT80), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n542), .A2(G179), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n444), .A2(new_n528), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n550), .A2(new_n548), .A3(KEYINPUT21), .A4(G169), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n544), .A2(new_n547), .A3(new_n549), .A4(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n381), .A2(new_n510), .A3(new_n465), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n249), .A2(new_n209), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT19), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n209), .B(G68), .C1(new_n343), .C2(new_n344), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n249), .A2(G20), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n555), .B(new_n556), .C1(KEYINPUT19), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n288), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n336), .A2(new_n361), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n478), .A2(G87), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(G250), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n440), .B1(new_n563), .B2(KEYINPUT77), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(new_n208), .A3(G45), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n434), .A2(KEYINPUT77), .A3(G250), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n323), .A2(new_n324), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n220), .A2(G1698), .ZN(new_n568));
  OAI221_X1 g0368(.A(new_n568), .B1(G238), .B2(G1698), .C1(new_n343), .C2(new_n344), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G116), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n257), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(G200), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n562), .A2(KEYINPUT78), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT78), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n565), .A2(new_n566), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n267), .B2(new_n269), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n569), .A2(new_n570), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n258), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n543), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n574), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n567), .A2(new_n571), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G190), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n573), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n582), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n364), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n582), .A2(new_n518), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n559), .B(new_n560), .C1(new_n336), .C2(new_n479), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n552), .A2(new_n590), .ZN(new_n591));
  AND4_X1   g0391(.A1(new_n432), .A2(new_n493), .A3(new_n521), .A4(new_n591), .ZN(G372));
  NAND2_X1  g0392(.A1(new_n520), .A2(KEYINPUT84), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT26), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n579), .A2(new_n580), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n583), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT84), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n515), .A2(new_n516), .A3(new_n597), .A4(new_n519), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n593), .A2(new_n594), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n484), .B1(new_n452), .B2(new_n453), .ZN(new_n600));
  AND4_X1   g0400(.A1(new_n549), .A2(new_n600), .A3(new_n547), .A4(new_n551), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n475), .A2(new_n481), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n602), .A2(new_n489), .A3(new_n483), .A4(new_n490), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n603), .A2(new_n514), .A3(new_n520), .A4(new_n596), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n599), .B(new_n589), .C1(new_n601), .C2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n520), .A2(new_n590), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(new_n594), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n432), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n412), .A2(new_n414), .ZN(new_n610));
  INV_X1    g0410(.A(new_n312), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n430), .B1(new_n319), .B2(new_n320), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n425), .A2(new_n420), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n372), .A2(new_n373), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n367), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n609), .A2(new_n617), .ZN(G369));
  NAND3_X1  g0418(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n303), .A2(new_n209), .ZN(new_n621));
  OR3_X1    g0421(.A1(new_n621), .A2(KEYINPUT85), .A3(KEYINPUT27), .ZN(new_n622));
  INV_X1    g0422(.A(G213), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n621), .B2(KEYINPUT27), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT85), .B1(new_n621), .B2(KEYINPUT27), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(G343), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n539), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n620), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g0431(.A(new_n552), .B(KEYINPUT86), .Z(new_n632));
  OAI21_X1  g0432(.A(new_n631), .B1(new_n632), .B2(new_n630), .ZN(new_n633));
  XOR2_X1   g0433(.A(new_n633), .B(KEYINPUT87), .Z(new_n634));
  INV_X1    g0434(.A(new_n488), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n493), .B1(new_n635), .B2(new_n629), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n458), .A2(new_n488), .A3(new_n628), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n634), .A2(G330), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n600), .A2(new_n628), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n620), .A2(new_n628), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n640), .B1(new_n641), .B2(new_n493), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT88), .ZN(G399));
  INV_X1    g0444(.A(new_n225), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(G41), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n553), .A2(G116), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G1), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n228), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT28), .ZN(new_n651));
  INV_X1    g0451(.A(new_n589), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n606), .B2(new_n594), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n619), .B1(new_n458), .B2(new_n488), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(new_n604), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n520), .A2(KEYINPUT84), .B1(new_n595), .B2(new_n583), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n594), .B1(new_n656), .B2(new_n598), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n629), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT89), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(KEYINPUT89), .B(new_n629), .C1(new_n655), .C2(new_n657), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(KEYINPUT29), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT29), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n608), .A2(new_n663), .A3(new_n629), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n493), .A2(new_n591), .A3(new_n521), .A4(new_n629), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n517), .A2(new_n450), .A3(new_n500), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n444), .A2(new_n528), .A3(G179), .A4(new_n582), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT30), .ZN(new_n669));
  OR3_X1    g0469(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(G179), .B1(new_n517), .B2(new_n500), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n671), .A2(new_n455), .A3(new_n585), .A4(new_n550), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n669), .B1(new_n667), .B2(new_n668), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT31), .B1(new_n674), .B2(new_n628), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(KEYINPUT31), .A3(new_n628), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n666), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n665), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n651), .B1(new_n681), .B2(G1), .ZN(G364));
  NOR2_X1   g0482(.A1(new_n302), .A2(G20), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G45), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n647), .A2(G1), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n634), .B2(G330), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(G330), .B2(new_n634), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n229), .B1(G20), .B2(new_n364), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n209), .A2(new_n314), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n691), .A2(new_n518), .A3(G200), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(G179), .A2(G200), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n209), .B1(new_n694), .B2(G190), .ZN(new_n695));
  OAI22_X1  g0495(.A1(new_n693), .A2(new_n242), .B1(new_n695), .B2(new_n510), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n518), .B2(G200), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n543), .A2(KEYINPUT92), .A3(G179), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n209), .A2(G190), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G107), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n700), .A2(new_n691), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n705), .B(new_n250), .C1(new_n381), .C2(new_n707), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT93), .Z(new_n709));
  NAND3_X1  g0509(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G190), .ZN(new_n711));
  AOI211_X1 g0511(.A(new_n696), .B(new_n709), .C1(G68), .C2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n702), .A2(new_n694), .ZN(new_n713));
  INV_X1    g0513(.A(G159), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT32), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n710), .A2(new_n314), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n712), .B(new_n716), .C1(new_n218), .C2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n702), .A2(G179), .A3(new_n543), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT91), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(KEYINPUT91), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n719), .B1(G77), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n720), .ZN(new_n725));
  INV_X1    g0525(.A(new_n713), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n725), .A2(G311), .B1(new_n726), .B2(G329), .ZN(new_n727));
  INV_X1    g0527(.A(G303), .ZN(new_n728));
  OAI221_X1 g0528(.A(new_n727), .B1(new_n448), .B2(new_n695), .C1(new_n707), .C2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n711), .ZN(new_n730));
  INV_X1    g0530(.A(G317), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n730), .B1(KEYINPUT33), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(KEYINPUT33), .B2(new_n731), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n250), .B1(new_n717), .B2(G326), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G322), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n693), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G283), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n703), .A2(new_n738), .ZN(new_n739));
  NOR4_X1   g0539(.A1(new_n729), .A2(new_n735), .A3(new_n737), .A4(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n689), .B1(new_n724), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(G355), .A2(new_n225), .A3(new_n250), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n243), .A2(G45), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n645), .A2(new_n250), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G45), .B2(new_n228), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n742), .B1(G116), .B2(new_n225), .C1(new_n743), .C2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT90), .Z(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n689), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n685), .B1(new_n633), .B2(new_n750), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n741), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n688), .A2(new_n754), .ZN(G396));
  NAND2_X1  g0555(.A1(new_n340), .A2(new_n628), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n341), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n430), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n430), .A2(new_n628), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n749), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n689), .A2(new_n747), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT94), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n202), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n703), .A2(new_n381), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n693), .A2(new_n448), .B1(new_n695), .B2(new_n510), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n250), .B1(new_n768), .B2(KEYINPUT95), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n769), .B1(KEYINPUT95), .B2(new_n768), .C1(new_n738), .C2(new_n730), .ZN(new_n770));
  INV_X1    g0570(.A(new_n723), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n469), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n718), .A2(new_n728), .ZN(new_n773));
  INV_X1    g0573(.A(G311), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n707), .A2(new_n465), .B1(new_n774), .B2(new_n713), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n770), .A2(new_n772), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G132), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n707), .A2(new_n218), .B1(new_n777), .B2(new_n713), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n703), .A2(new_n214), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n695), .A2(new_n242), .ZN(new_n780));
  NOR4_X1   g0580(.A1(new_n778), .A2(new_n779), .A3(new_n345), .A4(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT97), .Z(new_n782));
  AOI22_X1  g0582(.A1(new_n723), .A2(G159), .B1(G143), .B2(new_n692), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n717), .A2(G137), .ZN(new_n784));
  INV_X1    g0584(.A(G150), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n783), .B(new_n784), .C1(new_n785), .C2(new_n730), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT96), .B(KEYINPUT34), .Z(new_n787));
  XNOR2_X1  g0587(.A(new_n786), .B(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n767), .A2(new_n776), .B1(new_n782), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n689), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n765), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n686), .B1(new_n762), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n761), .B1(new_n608), .B2(new_n629), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n629), .B(new_n761), .C1(new_n605), .C2(new_n607), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(new_n679), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n792), .B1(new_n797), .B2(new_n686), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT98), .Z(G384));
  INV_X1    g0599(.A(KEYINPUT100), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n311), .A2(new_n629), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n800), .B(new_n802), .C1(new_n321), .C2(new_n286), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n284), .A2(new_n285), .ZN(new_n804));
  AND3_X1   g0604(.A1(new_n313), .A2(KEYINPUT72), .A3(new_n316), .ZN(new_n805));
  AOI21_X1  g0605(.A(KEYINPUT72), .B1(new_n313), .B2(new_n316), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n804), .B(new_n277), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(KEYINPUT100), .B1(new_n807), .B2(new_n801), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n312), .A2(new_n321), .A3(new_n802), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n809), .A2(new_n810), .B1(new_n794), .B2(new_n759), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n413), .B1(new_n388), .B2(new_n389), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT37), .ZN(new_n813));
  INV_X1    g0613(.A(new_n626), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n411), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n812), .A2(new_n423), .A3(new_n813), .A4(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n418), .B1(new_n416), .B2(new_n364), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n402), .B(new_n404), .C1(new_n339), .C2(new_n403), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n814), .ZN(new_n820));
  AND3_X1   g0620(.A1(new_n812), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n816), .B1(new_n821), .B2(new_n813), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n428), .B2(new_n820), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT38), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(KEYINPUT38), .B(new_n822), .C1(new_n428), .C2(new_n820), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n811), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n425), .A2(new_n420), .A3(new_n626), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT101), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n825), .A2(KEYINPUT39), .A3(new_n826), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n812), .A2(new_n423), .A3(new_n815), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(new_n813), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n815), .B1(new_n610), .B2(new_n614), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n824), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT39), .B1(new_n836), .B2(new_n826), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n611), .A2(new_n629), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT101), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n828), .A2(new_n842), .A3(new_n829), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n831), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT102), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n665), .B2(new_n432), .ZN(new_n846));
  AOI211_X1 g0646(.A(KEYINPUT102), .B(new_n431), .C1(new_n662), .C2(new_n664), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n617), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n844), .B(new_n848), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n674), .A2(KEYINPUT31), .A3(new_n628), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(new_n675), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n760), .B1(new_n851), .B2(new_n666), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n807), .A2(new_n801), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n800), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n807), .A2(KEYINPUT100), .A3(new_n801), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(new_n810), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n827), .A2(new_n852), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT40), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n856), .A2(new_n852), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n858), .B1(new_n836), .B2(new_n826), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n857), .A2(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n432), .A2(new_n678), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n861), .B(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n863), .A2(G330), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n849), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n208), .B2(new_n683), .ZN(new_n866));
  OAI211_X1 g0666(.A(G20), .B(new_n255), .C1(new_n506), .C2(KEYINPUT35), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n469), .B(new_n867), .C1(KEYINPUT35), .C2(new_n506), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT36), .Z(new_n869));
  NAND2_X1  g0669(.A1(new_n201), .A2(G68), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT99), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n396), .A2(new_n228), .A3(new_n202), .ZN(new_n872));
  OAI211_X1 g0672(.A(G1), .B(new_n302), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n866), .A2(new_n869), .A3(new_n873), .ZN(G367));
  NOR2_X1   g0674(.A1(new_n703), .A2(new_n202), .ZN(new_n875));
  XNOR2_X1  g0675(.A(KEYINPUT105), .B(G137), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n726), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n707), .B2(new_n242), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n875), .B(new_n878), .C1(G143), .C2(new_n717), .ZN(new_n879));
  INV_X1    g0679(.A(new_n201), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n723), .A2(new_n880), .B1(G159), .B2(new_n711), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n695), .A2(new_n214), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n692), .B2(G150), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT104), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n879), .A2(new_n250), .A3(new_n881), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n704), .A2(G97), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n886), .B1(new_n465), .B2(new_n695), .C1(new_n448), .C2(new_n730), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n250), .B(new_n887), .C1(G283), .C2(new_n723), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n692), .A2(new_n525), .B1(G311), .B2(new_n717), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n888), .B(new_n889), .C1(new_n731), .C2(new_n713), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n706), .A2(G116), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT46), .Z(new_n892));
  OAI21_X1  g0692(.A(new_n885), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT106), .Z(new_n894));
  AOI21_X1  g0694(.A(new_n790), .B1(new_n894), .B2(KEYINPUT47), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(KEYINPUT47), .B2(new_n894), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n628), .A2(new_n580), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n589), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n589), .A2(new_n596), .A3(new_n897), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n234), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n744), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n689), .B(new_n750), .C1(new_n645), .C2(new_n335), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n901), .A2(new_n750), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n896), .A2(new_n686), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n641), .A2(new_n493), .A3(new_n521), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT42), .Z(new_n908));
  OAI21_X1  g0708(.A(new_n521), .B1(new_n513), .B2(new_n629), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n458), .A2(new_n488), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n520), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n629), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT103), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT43), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(new_n900), .A3(new_n913), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n900), .B2(new_n915), .ZN(new_n917));
  INV_X1    g0717(.A(new_n639), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n520), .A2(new_n629), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n909), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n917), .A2(new_n921), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n684), .A2(G1), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n920), .A2(new_n642), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT45), .Z(new_n927));
  NOR2_X1   g0727(.A1(new_n920), .A2(new_n642), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT44), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n918), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n639), .A2(new_n927), .A3(new_n929), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n634), .A2(G330), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n641), .A2(new_n493), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n638), .B2(new_n641), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n934), .B(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n681), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n646), .B(KEYINPUT41), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n925), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n906), .B1(new_n924), .B2(new_n940), .ZN(G387));
  INV_X1    g0741(.A(new_n925), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n681), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n937), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT110), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n937), .A2(new_n944), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n647), .B1(new_n945), .B2(new_n946), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n943), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n723), .A2(new_n525), .B1(G317), .B2(new_n692), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n952), .B1(new_n774), .B2(new_n730), .C1(new_n736), .C2(new_n718), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT48), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n954), .B1(new_n738), .B2(new_n695), .C1(new_n448), .C2(new_n707), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT107), .Z(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT49), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n345), .B1(new_n703), .B2(new_n469), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(G326), .B2(new_n726), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT108), .Z(new_n960));
  NOR2_X1   g0760(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n693), .A2(new_n218), .B1(new_n214), .B2(new_n720), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n707), .A2(new_n202), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n962), .B(new_n963), .C1(new_n403), .C2(new_n711), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n785), .B2(new_n713), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n336), .A2(new_n695), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n886), .B1(new_n714), .B2(new_n718), .ZN(new_n967));
  NOR4_X1   g0767(.A1(new_n965), .A2(new_n345), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n689), .B1(new_n961), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n636), .A2(new_n637), .A3(new_n750), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n356), .A2(G50), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT50), .ZN(new_n972));
  NAND2_X1  g0772(.A1(G68), .A2(G77), .ZN(new_n973));
  AND4_X1   g0773(.A1(new_n261), .A2(new_n972), .A3(new_n973), .A4(new_n648), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n744), .B1(new_n238), .B2(new_n261), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n225), .B(new_n250), .C1(G116), .C2(new_n553), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n225), .A2(G107), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n751), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n969), .A2(new_n686), .A3(new_n970), .A4(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT109), .Z(new_n981));
  NAND2_X1  g0781(.A1(new_n951), .A2(new_n981), .ZN(G393));
  INV_X1    g0782(.A(KEYINPUT111), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n931), .A2(new_n983), .A3(new_n932), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n918), .A2(KEYINPUT111), .A3(new_n930), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT113), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n986), .A2(new_n948), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n987), .B1(new_n986), .B2(new_n948), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n948), .A2(new_n931), .A3(new_n932), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n988), .A2(new_n989), .A3(new_n646), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n986), .A2(new_n925), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n692), .A2(G311), .B1(new_n717), .B2(G317), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT52), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n250), .B1(new_n711), .B2(new_n525), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n705), .B(new_n995), .C1(new_n448), .C2(new_n720), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n994), .B(new_n996), .C1(G322), .C2(new_n726), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n469), .B2(new_n695), .C1(new_n738), .C2(new_n707), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n692), .A2(G159), .B1(new_n717), .B2(G150), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT51), .Z(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n202), .B2(new_n695), .C1(new_n356), .C2(new_n771), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n726), .A2(G143), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n880), .A2(new_n711), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n345), .B(new_n766), .C1(G68), .C2(new_n706), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n790), .B1(new_n998), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n751), .B1(new_n510), .B2(new_n225), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n247), .B2(new_n744), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT112), .Z(new_n1010));
  NOR3_X1   g0810(.A1(new_n1007), .A2(new_n685), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n750), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1011), .B1(new_n920), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n991), .A2(new_n992), .A3(new_n1013), .ZN(G390));
  NAND3_X1  g0814(.A1(new_n856), .A2(new_n680), .A3(new_n761), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n856), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n678), .A2(G330), .A3(new_n761), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n794), .A2(new_n759), .ZN(new_n1020));
  AND3_X1   g0820(.A1(new_n1019), .A2(KEYINPUT114), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(KEYINPUT114), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n660), .A2(new_n661), .A3(new_n759), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1023), .A2(new_n758), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n680), .B(new_n761), .C1(new_n856), .C2(KEYINPUT115), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n761), .A2(KEYINPUT115), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1016), .A2(new_n1017), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n1021), .A2(new_n1022), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n432), .A2(G330), .A3(new_n678), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n617), .B(new_n1030), .C1(new_n846), .C2(new_n847), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1023), .A2(new_n758), .A3(new_n856), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n840), .B1(new_n836), .B2(new_n826), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n832), .A2(new_n837), .B1(new_n811), .B2(new_n840), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1015), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1036), .A2(new_n1015), .A3(new_n1037), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1033), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g0843(.A1(new_n1036), .A2(new_n1015), .A3(new_n1037), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1015), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1046), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1043), .A2(new_n646), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n925), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n693), .A2(new_n777), .ZN(new_n1050));
  XOR2_X1   g0850(.A(KEYINPUT54), .B(G143), .Z(new_n1051));
  AOI22_X1  g0851(.A1(new_n723), .A2(new_n1051), .B1(G128), .B2(new_n717), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n345), .B1(new_n711), .B2(new_n876), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(new_n201), .C2(new_n703), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1050), .B(new_n1054), .C1(G125), .C2(new_n726), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n706), .A2(G150), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT53), .Z(new_n1057));
  OAI211_X1 g0857(.A(new_n1055), .B(new_n1057), .C1(new_n714), .C2(new_n695), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n707), .A2(new_n381), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n779), .B(new_n1059), .C1(G97), .C2(new_n723), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n717), .A2(G283), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n730), .A2(new_n465), .B1(new_n695), .B2(new_n202), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n250), .B(new_n1062), .C1(G294), .C2(new_n726), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n692), .A2(G116), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1060), .A2(new_n1061), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1058), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n686), .B1(new_n1066), .B2(new_n790), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n359), .B2(new_n764), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT116), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n838), .B2(new_n749), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1049), .A2(new_n1070), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1071), .A2(KEYINPUT117), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1071), .A2(KEYINPUT117), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1048), .B1(new_n1072), .B2(new_n1073), .ZN(G378));
  AOI21_X1  g0874(.A(KEYINPUT18), .B1(new_n817), .B2(new_n411), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n421), .B2(new_n420), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n427), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n610), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n820), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT38), .B1(new_n1080), .B2(new_n822), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n826), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n856), .A2(new_n852), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n858), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n859), .A2(new_n860), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(G330), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT120), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT120), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1085), .A2(new_n1086), .A3(new_n1089), .A4(G330), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n374), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n374), .A2(new_n1092), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n363), .A2(new_n814), .ZN(new_n1095));
  OR3_X1    g0895(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1095), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1088), .A2(new_n1090), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1098), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1100), .A2(KEYINPUT120), .A3(new_n1087), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1099), .A2(new_n844), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n844), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n925), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1100), .A2(new_n749), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n963), .B1(G116), .B2(new_n717), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1106), .B1(new_n242), .B2(new_n703), .C1(new_n465), .C2(new_n693), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n343), .A2(G41), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1108), .B1(new_n713), .B2(new_n738), .C1(new_n730), .C2(new_n510), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n1107), .A2(new_n344), .A3(new_n882), .A4(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n336), .B2(new_n720), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT58), .ZN(new_n1112));
  AOI21_X1  g0912(.A(G33), .B1(new_n726), .B2(G124), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n260), .B(new_n1113), .C1(new_n703), .C2(new_n714), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT118), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n717), .A2(G125), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n730), .B2(new_n777), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n725), .A2(G137), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(new_n706), .C2(new_n1051), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n692), .A2(G128), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1119), .B(new_n1120), .C1(new_n785), .C2(new_n695), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT59), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1112), .B1(G50), .B2(new_n1108), .C1(new_n1115), .C2(new_n1122), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT119), .Z(new_n1124));
  NOR2_X1   g0924(.A1(new_n1124), .A2(new_n790), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n763), .A2(new_n201), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NOR4_X1   g0927(.A1(new_n1105), .A2(new_n1125), .A3(new_n685), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1104), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1028), .A2(new_n1024), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT114), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1019), .A2(KEYINPUT114), .A3(new_n1020), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1131), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1032), .B1(new_n1136), .B2(new_n1042), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT57), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n647), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1031), .B1(new_n1046), .B2(new_n1029), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1141), .A2(new_n1139), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n844), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1090), .A2(new_n1098), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1089), .B1(new_n861), .B2(G330), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1100), .A2(KEYINPUT120), .A3(new_n1087), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1143), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT121), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1099), .A2(new_n844), .A3(new_n1101), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1103), .A2(KEYINPUT121), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1142), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1130), .B1(new_n1140), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(G375));
  INV_X1    g0955(.A(KEYINPUT122), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1136), .B2(new_n942), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1016), .A2(new_n747), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n764), .A2(new_n214), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n713), .A2(new_n728), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1160), .B(new_n875), .C1(G283), .C2(new_n692), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1161), .B1(new_n465), .B2(new_n771), .C1(new_n469), .C2(new_n730), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n707), .A2(new_n510), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n345), .B1(new_n718), .B2(new_n448), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1162), .A2(new_n966), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n692), .A2(new_n876), .B1(new_n711), .B2(new_n1051), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n777), .B2(new_n718), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT123), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1167), .A2(new_n1168), .B1(G58), .B2(new_n704), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n720), .A2(new_n785), .B1(new_n695), .B2(new_n218), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n706), .B2(G159), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n250), .A3(new_n1172), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1169), .B(new_n1173), .C1(G128), .C2(new_n726), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n689), .B1(new_n1165), .B2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1158), .A2(new_n686), .A3(new_n1159), .A4(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1029), .A2(KEYINPUT122), .A3(new_n925), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1157), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1136), .A2(new_n1031), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n1033), .A3(new_n939), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1180), .ZN(G381));
  AND2_X1   g0981(.A1(G375), .A2(KEYINPUT124), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(G375), .A2(KEYINPUT124), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1071), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1048), .A2(new_n1184), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(G381), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(G390), .A2(G384), .ZN(new_n1188));
  INV_X1    g0988(.A(G396), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n951), .A2(new_n1189), .A3(new_n981), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1190), .A2(G387), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .A4(new_n1191), .ZN(G407));
  AOI21_X1  g0992(.A(new_n623), .B1(new_n1186), .B2(new_n627), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(G407), .ZN(G409));
  AOI21_X1  g0994(.A(new_n1141), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1128), .B1(new_n1195), .B2(new_n939), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1151), .A2(new_n925), .A3(new_n1152), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1185), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1140), .A2(new_n1153), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1130), .ZN(new_n1201));
  AND4_X1   g1001(.A1(KEYINPUT125), .A2(new_n1200), .A3(G378), .A4(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT125), .B1(new_n1154), .B2(G378), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1199), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n623), .A2(G343), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT60), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1179), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1136), .A2(KEYINPUT60), .A3(new_n1031), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1208), .A2(new_n646), .A3(new_n1033), .A4(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(G384), .B1(new_n1210), .B2(new_n1178), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1178), .A3(G384), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1204), .A2(new_n1206), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT62), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT61), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1205), .A2(G2897), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1214), .B(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n646), .B1(new_n1195), .B2(KEYINPUT57), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1142), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1222));
  OAI211_X1 g1022(.A(G378), .B(new_n1201), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT125), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1154), .A2(KEYINPUT125), .A3(G378), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1198), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1220), .B1(new_n1227), .B2(new_n1205), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT62), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1204), .A2(new_n1229), .A3(new_n1206), .A4(new_n1215), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1217), .A2(new_n1218), .A3(new_n1228), .A4(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(G387), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(G390), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(G387), .A2(new_n991), .A3(new_n992), .A4(new_n1013), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1190), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1189), .B1(new_n951), .B2(new_n981), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT127), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n1232), .B2(G390), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1235), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1237), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1190), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1243), .A2(new_n1239), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1231), .A2(new_n1246), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1228), .A2(new_n1245), .A3(new_n1218), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1227), .A2(new_n1205), .A3(new_n1214), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT126), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT63), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1216), .A2(KEYINPUT126), .A3(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1248), .A2(new_n1251), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1247), .A2(new_n1254), .ZN(G405));
  NAND2_X1  g1055(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1154), .A2(new_n1185), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(new_n1215), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(new_n1246), .ZN(G402));
endmodule


