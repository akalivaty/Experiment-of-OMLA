//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XOR2_X1   g0005(.A(KEYINPUT66), .B(G77), .Z(new_n206));
  INV_X1    g0006(.A(G244), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G87), .A2(G250), .ZN(new_n212));
  NAND4_X1  g0012(.A1(new_n209), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n205), .B1(new_n208), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT1), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n216), .A2(G50), .A3(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OR3_X1    g0024(.A1(new_n205), .A2(KEYINPUT64), .A3(G13), .ZN(new_n225));
  OAI21_X1  g0025(.A(KEYINPUT64), .B1(new_n205), .B2(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  INV_X1    g0029(.A(G264), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n224), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n223), .B1(new_n231), .B2(KEYINPUT0), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n215), .B(new_n232), .C1(KEYINPUT0), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT69), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(new_n239), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  XOR2_X1   g0046(.A(KEYINPUT70), .B(G50), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G97), .B(G107), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n254));
  INV_X1    g0054(.A(G274), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n258), .A2(new_n254), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n256), .B1(new_n259), .B2(G232), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT78), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  AOI21_X1  g0064(.A(KEYINPUT78), .B1(new_n264), .B2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(G33), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G223), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(G226), .B2(new_n269), .ZN(new_n271));
  INV_X1    g0071(.A(G87), .ZN(new_n272));
  OAI22_X1  g0072(.A1(new_n267), .A2(new_n271), .B1(new_n262), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n257), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n260), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G169), .ZN(new_n276));
  INV_X1    g0076(.A(G179), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n276), .B1(new_n277), .B2(new_n275), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n220), .ZN(new_n281));
  INV_X1    g0081(.A(G58), .ZN(new_n282));
  INV_X1    g0082(.A(G68), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(G20), .B1(new_n284), .B2(new_n201), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G159), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT7), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n264), .A2(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n288), .B1(new_n296), .B2(G68), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n281), .B1(new_n297), .B2(KEYINPUT16), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT79), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n267), .A2(new_n221), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n283), .B1(new_n301), .B2(KEYINPUT7), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n267), .A2(new_n289), .A3(new_n221), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n288), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n300), .B1(new_n304), .B2(KEYINPUT16), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n264), .A2(KEYINPUT78), .A3(G33), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n261), .B1(new_n262), .B2(KEYINPUT3), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n306), .B1(new_n292), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT7), .B1(new_n308), .B2(G20), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(G68), .A3(new_n303), .ZN(new_n310));
  INV_X1    g0110(.A(new_n288), .ZN(new_n311));
  AND4_X1   g0111(.A1(new_n300), .A2(new_n310), .A3(KEYINPUT16), .A4(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n299), .B1(new_n305), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n221), .A2(G1), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G13), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT8), .B(G58), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n281), .B(KEYINPUT71), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n314), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n317), .B1(new_n319), .B2(new_n316), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n313), .A2(KEYINPUT80), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT80), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n307), .A2(new_n292), .ZN(new_n323));
  AOI21_X1  g0123(.A(G20), .B1(new_n323), .B2(new_n263), .ZN(new_n324));
  OAI21_X1  g0124(.A(G68), .B1(new_n324), .B2(new_n289), .ZN(new_n325));
  INV_X1    g0125(.A(new_n303), .ZN(new_n326));
  OAI211_X1 g0126(.A(KEYINPUT16), .B(new_n311), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT79), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n310), .A2(new_n300), .A3(KEYINPUT16), .A4(new_n311), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n298), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n320), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n322), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n279), .B1(new_n321), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT18), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT17), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n330), .A2(new_n331), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n275), .A2(G200), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n338), .A2(KEYINPUT81), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(KEYINPUT81), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n337), .B1(new_n275), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n335), .B1(new_n336), .B2(new_n343), .ZN(new_n344));
  NOR4_X1   g0144(.A1(new_n330), .A2(new_n342), .A3(KEYINPUT17), .A4(new_n331), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n333), .A2(new_n334), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI211_X1 g0146(.A(KEYINPUT18), .B(new_n279), .C1(new_n321), .C2(new_n332), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XOR2_X1   g0148(.A(KEYINPUT15), .B(G87), .Z(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(new_n221), .A3(G33), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT73), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n350), .B(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT72), .ZN(new_n353));
  INV_X1    g0153(.A(new_n286), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n316), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n353), .B2(new_n354), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n352), .B(new_n356), .C1(new_n221), .C2(new_n206), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n281), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n281), .A2(new_n314), .ZN(new_n359));
  INV_X1    g0159(.A(G77), .ZN(new_n360));
  INV_X1    g0160(.A(new_n206), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n359), .A2(new_n360), .B1(new_n361), .B2(new_n315), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT74), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT74), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n358), .A2(new_n366), .A3(new_n363), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n290), .A2(G232), .A3(new_n269), .ZN(new_n368));
  INV_X1    g0168(.A(G107), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n290), .A2(G1698), .ZN(new_n370));
  INV_X1    g0170(.A(G238), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n368), .B1(new_n369), .B2(new_n290), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n257), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n256), .B1(new_n259), .B2(G244), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(G190), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n374), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G200), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n365), .A2(new_n367), .A3(new_n375), .A4(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n376), .A2(G179), .ZN(new_n379));
  INV_X1    g0179(.A(G169), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(new_n376), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n366), .B1(new_n358), .B2(new_n363), .ZN(new_n382));
  AOI211_X1 g0182(.A(KEYINPUT74), .B(new_n362), .C1(new_n357), .C2(new_n281), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n385));
  INV_X1    g0185(.A(G150), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n221), .A2(G33), .ZN(new_n387));
  OAI221_X1 g0187(.A(new_n385), .B1(new_n386), .B2(new_n354), .C1(new_n316), .C2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G50), .ZN(new_n389));
  INV_X1    g0189(.A(new_n315), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n388), .A2(new_n318), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n319), .A2(G50), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n290), .A2(G222), .A3(new_n269), .ZN(new_n394));
  OAI221_X1 g0194(.A(new_n394), .B1(new_n206), .B2(new_n290), .C1(new_n370), .C2(new_n268), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n257), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n256), .B1(new_n259), .B2(G226), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n393), .B1(new_n399), .B2(G169), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n398), .A2(G179), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n378), .A2(new_n384), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n393), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(KEYINPUT9), .B1(new_n399), .B2(G190), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT9), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n393), .A2(new_n407), .B1(new_n398), .B2(G200), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT10), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT10), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n406), .A2(new_n411), .A3(new_n408), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n404), .A2(new_n413), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n387), .A2(new_n360), .B1(new_n221), .B2(G68), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n415), .A2(KEYINPUT75), .B1(G50), .B2(new_n286), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(KEYINPUT75), .B2(new_n415), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n318), .ZN(new_n418));
  XOR2_X1   g0218(.A(new_n418), .B(KEYINPUT11), .Z(new_n419));
  NAND2_X1  g0219(.A1(new_n390), .A2(new_n283), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT76), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT12), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(KEYINPUT12), .B2(new_n420), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n421), .B1(new_n420), .B2(KEYINPUT12), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n423), .A2(new_n424), .B1(new_n283), .B2(new_n359), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT77), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n256), .B1(new_n259), .B2(G238), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n290), .A2(G232), .A3(G1698), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n290), .A2(G226), .A3(new_n269), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G97), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n257), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n435), .A2(KEYINPUT13), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(KEYINPUT13), .ZN(new_n437));
  OAI21_X1  g0237(.A(G169), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n436), .A2(new_n437), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n438), .A2(KEYINPUT14), .B1(new_n439), .B2(G179), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT14), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(G169), .C1(new_n436), .C2(new_n437), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n428), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n438), .A2(KEYINPUT14), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n439), .A2(G179), .ZN(new_n445));
  AND4_X1   g0245(.A1(new_n428), .A2(new_n444), .A3(new_n442), .A4(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n427), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n427), .B1(G190), .B2(new_n439), .ZN(new_n448));
  INV_X1    g0248(.A(G200), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n448), .B1(new_n449), .B2(new_n439), .ZN(new_n450));
  AND4_X1   g0250(.A1(new_n348), .A2(new_n414), .A3(new_n447), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G283), .ZN(new_n452));
  INV_X1    g0252(.A(G97), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n452), .B(new_n221), .C1(G33), .C2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n454), .B(new_n281), .C1(new_n221), .C2(G116), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT20), .ZN(new_n456));
  OR3_X1    g0256(.A1(new_n455), .A2(KEYINPUT86), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n456), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT86), .B1(new_n455), .B2(new_n456), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n315), .B1(G1), .B2(new_n262), .ZN(new_n461));
  INV_X1    g0261(.A(G116), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n461), .A2(new_n462), .A3(new_n281), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n462), .B2(new_n390), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n230), .A2(G1698), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(G257), .B2(G1698), .ZN(new_n467));
  INV_X1    g0267(.A(G303), .ZN(new_n468));
  OAI22_X1  g0268(.A1(new_n267), .A2(new_n467), .B1(new_n468), .B2(new_n290), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n257), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n257), .A2(new_n255), .ZN(new_n471));
  INV_X1    g0271(.A(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G1), .ZN(new_n473));
  INV_X1    g0273(.A(G41), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n473), .B(KEYINPUT83), .C1(KEYINPUT5), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(KEYINPUT5), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n253), .B(G45), .C1(new_n474), .C2(KEYINPUT5), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT83), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n471), .A2(new_n475), .A3(new_n476), .A4(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n470), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n475), .A2(new_n479), .A3(new_n476), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n258), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G270), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n465), .B1(G200), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n341), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n481), .A2(new_n488), .A3(new_n485), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n486), .A2(new_n465), .A3(G169), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT21), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n486), .A2(new_n465), .A3(KEYINPUT21), .A4(G169), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n465), .A2(G179), .A3(new_n485), .A4(new_n481), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n490), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT87), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n494), .A2(new_n495), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT87), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(new_n493), .A4(new_n490), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n229), .A2(G1698), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(G250), .B2(G1698), .ZN(new_n503));
  INV_X1    g0303(.A(G294), .ZN(new_n504));
  OAI22_X1  g0304(.A1(new_n267), .A2(new_n503), .B1(new_n262), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n257), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n482), .A2(G264), .A3(new_n258), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(G179), .A3(new_n480), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT88), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n506), .A2(new_n507), .A3(new_n480), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G169), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n308), .A2(KEYINPUT22), .A3(new_n221), .A4(G87), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT22), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n221), .A2(G87), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n294), .B2(new_n516), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n262), .A2(new_n462), .A3(G20), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT23), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n221), .B2(G107), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n369), .A2(KEYINPUT23), .A3(G20), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n514), .A2(new_n517), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT24), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n514), .A2(KEYINPUT24), .A3(new_n517), .A4(new_n522), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n281), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n318), .A2(new_n461), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT25), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n315), .B2(G107), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n390), .A2(KEYINPUT25), .A3(new_n369), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n528), .A2(G107), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n510), .B1(new_n509), .B2(new_n512), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n513), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n511), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G190), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n511), .A2(G200), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n538), .A2(new_n527), .A3(new_n532), .A4(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n528), .A2(G97), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n390), .A2(new_n453), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g0345(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(G97), .A3(new_n369), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n249), .B2(new_n546), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(G20), .B1(G77), .B2(new_n286), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n296), .A2(G107), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n545), .B1(new_n551), .B2(new_n281), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n290), .A2(KEYINPUT4), .A3(G244), .A4(new_n269), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n290), .A2(G250), .A3(G1698), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n553), .A2(new_n452), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT4), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n269), .A2(G244), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(new_n267), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n258), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n480), .B1(new_n483), .B2(new_n229), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G190), .ZN(new_n562));
  OAI21_X1  g0362(.A(G200), .B1(new_n559), .B2(new_n560), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n552), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n551), .A2(new_n281), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n543), .A2(new_n544), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n561), .A2(new_n277), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n380), .B1(new_n559), .B2(new_n560), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n272), .A2(new_n453), .A3(new_n369), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n572), .B(KEYINPUT85), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT19), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n221), .B1(new_n432), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n308), .A2(new_n221), .A3(G68), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n574), .B1(new_n387), .B2(new_n453), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n349), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n579), .A2(new_n281), .B1(new_n390), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n207), .A2(G1698), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(G238), .B2(G1698), .ZN(new_n583));
  OAI22_X1  g0383(.A1(new_n267), .A2(new_n583), .B1(new_n262), .B2(new_n462), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n257), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n257), .A2(new_n224), .A3(new_n473), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(G274), .B2(new_n473), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G200), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n528), .A2(G87), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n581), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n588), .A2(new_n338), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n588), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G179), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n380), .B1(new_n585), .B2(new_n587), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(KEYINPUT84), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT84), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n588), .A2(new_n277), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n600), .B2(new_n596), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n528), .A2(new_n349), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n581), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n598), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n571), .A2(new_n593), .A3(new_n604), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n451), .A2(new_n501), .A3(new_n542), .A4(new_n605), .ZN(G372));
  NAND3_X1  g0406(.A1(new_n410), .A2(KEYINPUT90), .A3(new_n412), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT90), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n413), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n345), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n313), .A2(new_n343), .A3(new_n320), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT17), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n384), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n450), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n614), .B1(new_n616), .B2(new_n447), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n278), .B1(new_n330), .B2(new_n331), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n334), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n278), .B(KEYINPUT18), .C1(new_n330), .C2(new_n331), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n607), .B(new_n609), .C1(new_n617), .C2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n623), .A2(new_n403), .ZN(new_n624));
  INV_X1    g0424(.A(new_n570), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n593), .A3(new_n604), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT26), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n595), .A2(new_n597), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n603), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n581), .A2(new_n590), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(KEYINPUT89), .A3(new_n589), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT89), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n592), .B1(new_n591), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n625), .A3(new_n629), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n627), .B(new_n629), .C1(new_n635), .C2(KEYINPUT26), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n509), .A2(new_n512), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n533), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n498), .A2(new_n493), .A3(new_n638), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n631), .A2(new_n633), .B1(new_n628), .B2(new_n603), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n564), .A2(new_n570), .A3(new_n540), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n451), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n624), .A2(new_n644), .ZN(G369));
  INV_X1    g0445(.A(G13), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(G20), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n253), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G213), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n465), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n501), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n498), .A2(new_n493), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(new_n654), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n653), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n542), .B1(new_n534), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n536), .A2(new_n653), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n638), .A2(new_n653), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n658), .A2(new_n653), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(new_n542), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(G399));
  NOR2_X1   g0472(.A1(new_n573), .A2(G116), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n228), .A2(G41), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n674), .A2(new_n675), .A3(new_n253), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n219), .B2(new_n675), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT91), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT28), .Z(new_n679));
  NOR2_X1   g0479(.A1(new_n486), .A2(new_n277), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n680), .A2(new_n508), .A3(new_n561), .A4(new_n594), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT30), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n486), .A2(new_n277), .A3(new_n588), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT92), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n561), .A2(new_n537), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n681), .A2(new_n682), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n683), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n691), .A2(new_n692), .A3(new_n653), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n501), .A2(new_n605), .A3(new_n542), .A4(new_n664), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n692), .B1(new_n691), .B2(new_n653), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n643), .A2(new_n664), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT29), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT26), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n625), .A2(new_n593), .A3(new_n604), .A4(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n703), .A2(new_n629), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n641), .B(new_n640), .C1(new_n657), .C2(new_n536), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n635), .A2(KEYINPUT26), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n707), .A2(KEYINPUT29), .A3(new_n664), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n698), .B1(new_n701), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n679), .B1(new_n709), .B2(G1), .ZN(G364));
  AOI21_X1  g0510(.A(new_n253), .B1(new_n647), .B2(G45), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n675), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n661), .A2(G330), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n713), .B1(new_n715), .B2(new_n662), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n380), .A2(KEYINPUT93), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n221), .B1(KEYINPUT93), .B2(new_n380), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n220), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G13), .A2(G33), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT94), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n228), .A2(new_n308), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n248), .A2(new_n472), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n728), .B(new_n729), .C1(new_n472), .C2(new_n219), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n227), .A2(new_n290), .ZN(new_n731));
  INV_X1    g0531(.A(G355), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n731), .A2(new_n732), .B1(G116), .B2(new_n227), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n726), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n221), .A2(new_n277), .A3(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n488), .A2(new_n735), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n221), .A2(new_n277), .A3(new_n449), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n338), .ZN(new_n738));
  OAI22_X1  g0538(.A1(new_n736), .A2(new_n282), .B1(new_n738), .B2(new_n283), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n488), .A2(new_n737), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n735), .A2(new_n338), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n741), .A2(G50), .B1(new_n361), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G179), .A2(G200), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n746), .A2(new_n221), .A3(G190), .ZN(new_n747));
  XNOR2_X1  g0547(.A(KEYINPUT95), .B(G159), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n744), .B(new_n290), .C1(KEYINPUT32), .C2(new_n749), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n739), .B(new_n750), .C1(KEYINPUT32), .C2(new_n749), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n221), .A2(G179), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(new_n338), .A3(G200), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT97), .Z(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n369), .ZN(new_n755));
  OAI21_X1  g0555(.A(G20), .B1(new_n746), .B2(new_n338), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT98), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n453), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n752), .A2(G190), .A3(G200), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n762), .A2(KEYINPUT96), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(KEYINPUT96), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n755), .B(new_n761), .C1(G87), .C2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n290), .B1(new_n747), .B2(G329), .ZN(new_n768));
  INV_X1    g0568(.A(G311), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n769), .B2(new_n742), .ZN(new_n770));
  INV_X1    g0570(.A(new_n738), .ZN(new_n771));
  NOR2_X1   g0571(.A1(KEYINPUT33), .A2(G317), .ZN(new_n772));
  AND2_X1   g0572(.A1(KEYINPUT33), .A2(G317), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n774), .B1(new_n775), .B2(new_n736), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT99), .B(G326), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n770), .B(new_n776), .C1(new_n741), .C2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n760), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n779), .A2(G294), .B1(new_n766), .B2(G303), .ZN(new_n780));
  INV_X1    g0580(.A(G283), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n781), .B2(new_n754), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n751), .A2(new_n767), .B1(new_n778), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n720), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n734), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(new_n660), .B2(new_n723), .ZN(new_n787));
  INV_X1    g0587(.A(new_n713), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n716), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT100), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n790), .B(new_n791), .ZN(G396));
  NOR2_X1   g0592(.A1(new_n720), .A2(new_n721), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n788), .B1(new_n360), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n267), .B1(new_n747), .B2(G132), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n741), .A2(G137), .B1(new_n743), .B2(new_n748), .ZN(new_n796));
  INV_X1    g0596(.A(G143), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n796), .B1(new_n797), .B2(new_n736), .C1(new_n386), .C2(new_n738), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT34), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n795), .B1(new_n282), .B2(new_n760), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n799), .B2(new_n798), .ZN(new_n801));
  INV_X1    g0601(.A(new_n754), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G68), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n389), .B2(new_n765), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT101), .Z(new_n805));
  INV_X1    g0605(.A(new_n747), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n294), .B1(new_n806), .B2(new_n769), .C1(new_n736), .C2(new_n504), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n740), .A2(new_n468), .B1(new_n738), .B2(new_n781), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n807), .B(new_n808), .C1(G116), .C2(new_n743), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n754), .A2(new_n272), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n810), .B(new_n761), .C1(G107), .C2(new_n766), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n801), .A2(new_n805), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n384), .A2(new_n653), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n653), .B1(new_n382), .B2(new_n383), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n378), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n813), .B1(new_n815), .B2(new_n384), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n794), .B1(new_n812), .B2(new_n785), .C1(new_n816), .C2(new_n722), .ZN(new_n817));
  INV_X1    g0617(.A(new_n816), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n699), .A2(new_n818), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n816), .B(new_n664), .C1(new_n636), .C2(new_n642), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n820), .A2(KEYINPUT102), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n819), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n698), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT103), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n822), .A2(new_n697), .A3(new_n823), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n827), .A2(new_n788), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n825), .A2(new_n826), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n817), .B1(new_n829), .B2(new_n830), .ZN(G384));
  NAND3_X1  g0631(.A1(new_n701), .A2(new_n451), .A3(new_n708), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n624), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT106), .ZN(new_n834));
  INV_X1    g0634(.A(new_n651), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n318), .B1(new_n304), .B2(KEYINPUT16), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n329), .B2(new_n328), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n835), .B1(new_n837), .B2(new_n331), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n346), .B2(new_n347), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT80), .B1(new_n313), .B2(new_n320), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n330), .A2(new_n322), .A3(new_n331), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n278), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n835), .B1(new_n841), .B2(new_n842), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT37), .B1(new_n336), .B2(new_n343), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n278), .B1(new_n837), .B2(new_n331), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n838), .A2(new_n847), .A3(new_n611), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(KEYINPUT37), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n840), .A2(KEYINPUT38), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT38), .B1(new_n840), .B2(new_n850), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT39), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT104), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT104), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n855), .B(KEYINPUT39), .C1(new_n851), .C2(new_n852), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT105), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n651), .B1(new_n321), .B2(new_n332), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n611), .A2(new_n859), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n333), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n611), .A2(new_n618), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n859), .B1(new_n844), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n857), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n611), .A2(new_n618), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT37), .B1(new_n858), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n846), .A2(new_n866), .A3(KEYINPUT105), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n844), .B1(new_n613), .B2(new_n621), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n864), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT39), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n840), .A2(KEYINPUT38), .A3(new_n850), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n854), .A2(new_n856), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n447), .A2(new_n653), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n813), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n820), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n427), .A2(new_n653), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n447), .A2(new_n450), .A3(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n427), .B(new_n653), .C1(new_n443), .C2(new_n446), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n840), .A2(new_n850), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n871), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n885), .B1(new_n887), .B2(new_n874), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n621), .A2(new_n835), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n878), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n834), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n846), .A2(new_n866), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n868), .B1(new_n893), .B2(new_n857), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n894), .B2(new_n867), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT107), .B1(new_n895), .B2(new_n851), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT107), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n872), .A2(new_n897), .A3(new_n874), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n696), .A2(new_n884), .A3(KEYINPUT40), .A4(new_n816), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n696), .A2(new_n884), .A3(new_n816), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n887), .A2(new_n874), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT40), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n902), .A2(G330), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n698), .A2(new_n451), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n905), .B1(new_n899), .B2(new_n901), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n451), .A2(new_n696), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n907), .A2(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n892), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n913), .A2(KEYINPUT108), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(KEYINPUT108), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n647), .A2(new_n253), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n892), .B2(new_n911), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n548), .A2(KEYINPUT35), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(G116), .A3(new_n222), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(KEYINPUT35), .B2(new_n548), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT36), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n921), .A2(KEYINPUT36), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n206), .A2(new_n284), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n218), .A2(new_n924), .B1(G50), .B2(new_n283), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(G1), .A3(new_n646), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n918), .A2(new_n922), .A3(new_n923), .A4(new_n926), .ZN(G367));
  OAI21_X1  g0727(.A(new_n571), .B1(new_n552), .B2(new_n664), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n570), .B2(new_n664), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n542), .A3(new_n670), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT42), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(KEYINPUT109), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n536), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n570), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n931), .B1(new_n935), .B2(new_n664), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n640), .B1(new_n630), .B2(new_n664), .ZN(new_n937));
  OR3_X1    g0737(.A1(new_n629), .A2(new_n630), .A3(new_n664), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT43), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n936), .A2(KEYINPUT110), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT110), .B1(new_n936), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n668), .B2(new_n932), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n668), .A2(new_n932), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n947), .B(new_n941), .C1(new_n943), .C2(new_n944), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n675), .B(KEYINPUT41), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n709), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n670), .A2(new_n542), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n667), .B2(new_n670), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n662), .B(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n671), .A2(new_n929), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT45), .Z(new_n957));
  NOR2_X1   g0757(.A1(new_n671), .A2(new_n929), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT44), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(new_n663), .A3(new_n667), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n668), .A2(new_n957), .A3(new_n959), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n955), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n950), .B1(new_n963), .B2(new_n709), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n946), .B(new_n948), .C1(new_n964), .C2(new_n712), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n726), .B1(new_n227), .B2(new_n580), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n238), .A2(new_n728), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n713), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(G137), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n290), .B1(new_n806), .B2(new_n969), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n740), .A2(new_n797), .B1(new_n206), .B2(new_n753), .ZN(new_n971));
  INV_X1    g0771(.A(new_n736), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n970), .B(new_n971), .C1(G150), .C2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n779), .A2(G68), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(new_n282), .C2(new_n765), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n771), .A2(new_n748), .B1(new_n743), .B2(G50), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT112), .Z(new_n977));
  NAND3_X1  g0777(.A1(new_n766), .A2(KEYINPUT46), .A3(G116), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT46), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n765), .B2(new_n462), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n308), .B1(G317), .B2(new_n747), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n738), .A2(new_n504), .B1(new_n453), .B2(new_n753), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G283), .B2(new_n743), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n978), .A2(new_n980), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n468), .A2(new_n736), .B1(new_n740), .B2(new_n769), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT111), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G107), .A2(new_n779), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n986), .B2(new_n985), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n975), .A2(new_n977), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT47), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n785), .B1(new_n989), .B2(new_n990), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n968), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n723), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n939), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n965), .A2(new_n995), .ZN(G387));
  INV_X1    g0796(.A(new_n954), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n709), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n951), .A2(new_n954), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n998), .A2(new_n675), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n997), .A2(new_n712), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n316), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT50), .B1(new_n316), .B2(G50), .ZN(new_n1003));
  AOI21_X1  g0803(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n727), .B1(new_n674), .B2(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n243), .A2(G45), .B1(new_n1006), .B2(KEYINPUT113), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(KEYINPUT113), .B2(new_n1006), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(G107), .B2(new_n227), .C1(new_n673), .C2(new_n731), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n726), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n713), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n741), .A2(G159), .B1(G68), .B2(new_n743), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n389), .B2(new_n736), .C1(new_n316), .C2(new_n738), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n267), .B(new_n1013), .C1(G150), .C2(new_n747), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n766), .A2(new_n361), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n779), .A2(new_n349), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n802), .A2(G97), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n308), .B1(new_n747), .B2(new_n777), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G317), .A2(new_n972), .B1(new_n741), .B2(G322), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n468), .B2(new_n742), .C1(new_n769), .C2(new_n738), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT48), .Z(new_n1022));
  OAI22_X1  g0822(.A1(new_n760), .A2(new_n781), .B1(new_n765), .B2(new_n504), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1019), .B1(new_n462), .B2(new_n753), .C1(new_n1024), .C2(KEYINPUT49), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1024), .A2(KEYINPUT49), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1018), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1011), .B1(new_n1027), .B2(new_n720), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n667), .B2(new_n994), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1000), .A2(new_n1001), .A3(new_n1029), .ZN(G393));
  AOI22_X1  g0830(.A1(G311), .A2(new_n972), .B1(new_n741), .B2(G317), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1031), .A2(KEYINPUT52), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G116), .B2(new_n779), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n294), .B1(new_n504), .B2(new_n742), .C1(new_n806), .C2(new_n775), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1034), .B(new_n755), .C1(G303), .C2(new_n771), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1031), .A2(KEYINPUT52), .B1(G283), .B2(new_n766), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(G159), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n386), .A2(new_n740), .B1(new_n736), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT51), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n738), .A2(new_n389), .B1(new_n742), .B2(new_n316), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n308), .B1(new_n806), .B2(new_n797), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n810), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n766), .A2(G68), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n779), .A2(G77), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1040), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n785), .B1(new_n1037), .B2(new_n1046), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n728), .A2(new_n251), .B1(new_n453), .B2(new_n227), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n713), .B1(new_n1048), .B2(new_n725), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT114), .Z(new_n1050));
  AOI211_X1 g0850(.A(new_n1047), .B(new_n1050), .C1(new_n932), .C2(new_n723), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n961), .A2(new_n962), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1051), .B1(new_n1053), .B2(new_n712), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n675), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1053), .B2(new_n955), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n998), .A2(new_n1052), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1056), .A2(KEYINPUT115), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT115), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1054), .B1(new_n1059), .B2(new_n1060), .ZN(G390));
  NAND4_X1  g0861(.A1(new_n696), .A2(new_n884), .A3(G330), .A4(new_n816), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n877), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n885), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n854), .A2(new_n856), .A3(new_n875), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n815), .A2(new_n384), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n707), .A2(new_n664), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n879), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n884), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n1064), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n896), .B2(new_n898), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT116), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1066), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI211_X1 g0874(.A(KEYINPUT116), .B(new_n1071), .C1(new_n896), .C2(new_n898), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1063), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n877), .B1(new_n1069), .B2(new_n884), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n895), .A2(KEYINPUT107), .A3(new_n851), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n897), .B1(new_n872), .B2(new_n874), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(KEYINPUT116), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1062), .B(KEYINPUT117), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .A4(new_n1066), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1076), .A2(new_n712), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT119), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n741), .A2(G283), .B1(G97), .B2(new_n743), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n369), .B2(new_n738), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT118), .Z(new_n1089));
  NAND2_X1  g0889(.A1(new_n766), .A2(G87), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n294), .B1(new_n806), .B2(new_n504), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G116), .B2(new_n972), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1045), .A2(new_n803), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n766), .A2(G150), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT53), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n779), .A2(G159), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n738), .A2(new_n969), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n294), .B(new_n1097), .C1(G125), .C2(new_n747), .ZN(new_n1098));
  XOR2_X1   g0898(.A(KEYINPUT54), .B(G143), .Z(new_n1099));
  AOI22_X1  g0899(.A1(new_n741), .A2(G128), .B1(new_n743), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n753), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n972), .A2(G132), .B1(G50), .B2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .A4(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1089), .A2(new_n1093), .B1(new_n1095), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n720), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n788), .B1(new_n316), .B2(new_n793), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(new_n876), .C2(new_n722), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1085), .A2(new_n1086), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1086), .B1(new_n1085), .B2(new_n1107), .ZN(new_n1109));
  OAI21_X1  g0909(.A(KEYINPUT120), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1085), .A2(new_n1107), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(KEYINPUT119), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT120), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1085), .A2(new_n1086), .A3(new_n1107), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1076), .A2(new_n1084), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n624), .A2(new_n832), .A3(new_n908), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n884), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n696), .A2(new_n816), .ZN(new_n1120));
  INV_X1    g0920(.A(G330), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1069), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1083), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1062), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n880), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1118), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1117), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1076), .A2(new_n1127), .A3(new_n1084), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n675), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1116), .A2(new_n1131), .ZN(G378));
  NAND3_X1  g0932(.A1(new_n609), .A2(new_n403), .A3(new_n607), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n405), .A2(new_n651), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1134), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n609), .A2(new_n403), .A3(new_n607), .A4(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1135), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n721), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n974), .A2(new_n1015), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G97), .A2(new_n771), .B1(new_n743), .B2(new_n349), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1101), .A2(G58), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(new_n369), .C2(new_n736), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n308), .A2(G41), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n806), .B2(new_n781), .C1(new_n740), .C2(new_n462), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1143), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT58), .Z(new_n1150));
  NAND2_X1  g0950(.A1(new_n779), .A2(G150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n972), .A2(G128), .B1(G137), .B2(new_n743), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n741), .A2(G125), .B1(new_n771), .B2(G132), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n766), .A2(new_n1099), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1101), .A2(new_n748), .ZN(new_n1158));
  AOI211_X1 g0958(.A(G33), .B(G41), .C1(new_n747), .C2(G124), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n389), .B1(G33), .B2(G41), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1150), .B1(new_n1156), .B2(new_n1160), .C1(new_n1147), .C2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT121), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n785), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n1163), .B2(new_n1162), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n793), .A2(new_n389), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1142), .A2(new_n713), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n907), .A2(new_n1141), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n878), .A2(new_n890), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1141), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n909), .A2(G330), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1171), .B1(new_n909), .B2(G330), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n900), .B1(new_n896), .B2(new_n898), .ZN(new_n1175));
  NOR4_X1   g0975(.A1(new_n1175), .A2(new_n905), .A3(new_n1121), .A4(new_n1141), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n891), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1173), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1168), .B1(new_n1178), .B2(new_n712), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1118), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1130), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(KEYINPUT57), .A3(new_n1178), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n675), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT57), .B1(new_n1181), .B2(new_n1178), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1179), .B1(new_n1183), .B2(new_n1184), .ZN(G375));
  NAND3_X1  g0985(.A1(new_n1124), .A2(new_n1118), .A3(new_n1126), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1128), .A2(new_n949), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n788), .B1(new_n283), .B2(new_n793), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT122), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n741), .A2(G132), .B1(new_n771), .B2(new_n1099), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n386), .B2(new_n742), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n267), .B1(new_n747), .B2(G128), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n1145), .C1(new_n736), .C2(new_n969), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n760), .A2(new_n389), .B1(new_n765), .B2(new_n1038), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1016), .B1(new_n781), .B2(new_n736), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT123), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n754), .A2(new_n360), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n765), .A2(new_n453), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n294), .B1(new_n738), .B2(new_n462), .C1(new_n806), .C2(new_n468), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n740), .A2(new_n504), .B1(new_n369), .B2(new_n742), .ZN(new_n1201));
  NOR4_X1   g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1195), .B1(new_n1197), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1189), .B1(new_n1203), .B2(new_n785), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1119), .B2(new_n721), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1205), .B1(new_n1206), .B2(new_n712), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1187), .A2(new_n1207), .ZN(G381));
  INV_X1    g1008(.A(new_n1060), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1058), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1210), .A2(new_n995), .A3(new_n965), .A4(new_n1054), .ZN(new_n1211));
  OR2_X1    g1011(.A1(G393), .A2(G396), .ZN(new_n1212));
  OR3_X1    g1012(.A1(new_n1211), .A2(G384), .A3(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1131), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1214));
  OR2_X1    g1014(.A1(G375), .A2(new_n1214), .ZN(new_n1215));
  OR3_X1    g1015(.A1(new_n1213), .A2(new_n1215), .A3(G381), .ZN(G407));
  OAI211_X1 g1016(.A(G407), .B(G213), .C1(G343), .C2(new_n1215), .ZN(G409));
  NAND3_X1  g1017(.A1(new_n1181), .A2(new_n949), .A3(new_n1178), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n1179), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1219), .A2(new_n1131), .A3(new_n1114), .A4(new_n1112), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1131), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1220), .B1(new_n1222), .B2(G375), .ZN(new_n1223));
  INV_X1    g1023(.A(G213), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(G343), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT60), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1186), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1186), .A2(new_n1227), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1228), .A2(new_n675), .A3(new_n1128), .A4(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1230), .A2(new_n1207), .B1(KEYINPUT124), .B2(G384), .ZN(new_n1231));
  INV_X1    g1031(.A(G384), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT124), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1230), .A2(new_n1232), .A3(new_n1233), .A4(new_n1207), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1223), .A2(new_n1226), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(KEYINPUT62), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT61), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT62), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1223), .A2(new_n1241), .A3(new_n1226), .A4(new_n1237), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1225), .A2(G2897), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1235), .A2(new_n1236), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1218), .A2(new_n1179), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(new_n1214), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1179), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1180), .A2(new_n1130), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1055), .B1(new_n1250), .B2(KEYINPUT57), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1184), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1249), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1248), .B1(G378), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1246), .B1(new_n1254), .B2(new_n1225), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1239), .A2(new_n1240), .A3(new_n1242), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G393), .A2(G396), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1212), .A2(new_n1257), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1258), .A2(KEYINPUT125), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(KEYINPUT125), .ZN(new_n1260));
  AND2_X1   g1060(.A1(G390), .A2(G387), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(G390), .A2(G387), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1259), .B(new_n1260), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G390), .A2(G387), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1211), .A2(new_n1264), .A3(KEYINPUT125), .A4(new_n1258), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT127), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1266), .B(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1256), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT63), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1266), .B1(KEYINPUT126), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1238), .B1(KEYINPUT126), .B2(new_n1270), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT61), .B1(new_n1273), .B2(new_n1246), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1270), .A2(KEYINPUT126), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1223), .A2(new_n1226), .A3(new_n1237), .A4(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1271), .A2(new_n1272), .A3(new_n1274), .A4(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1269), .A2(new_n1277), .ZN(G405));
  NOR2_X1   g1078(.A1(new_n1222), .A2(G375), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1253), .A2(new_n1214), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1266), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1263), .B(new_n1265), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1237), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1284), .B(new_n1285), .ZN(G402));
endmodule


