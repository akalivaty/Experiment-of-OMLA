//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR3_X1   g0001(.A1(new_n201), .A2(G58), .A3(G68), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  NOR2_X1   g0010(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n211), .B1(new_n216), .B2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n217), .B(new_n218), .Z(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n210), .B(new_n219), .C1(new_n222), .C2(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT2), .B(G226), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G250), .B(G257), .Z(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n229), .B(new_n232), .Z(G358));
  XNOR2_X1  g0033(.A(G68), .B(G77), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G58), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT66), .B(G50), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G97), .B(G107), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G351));
  INV_X1    g0041(.A(G33), .ZN(new_n242));
  OAI21_X1  g0042(.A(KEYINPUT70), .B1(new_n242), .B2(G20), .ZN(new_n243));
  INV_X1    g0043(.A(KEYINPUT70), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n244), .A2(new_n221), .A3(G33), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n243), .A2(new_n245), .A3(G97), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT19), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G97), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n221), .B1(new_n248), .B2(new_n247), .ZN(new_n249));
  INV_X1    g0049(.A(G87), .ZN(new_n250));
  INV_X1    g0050(.A(G97), .ZN(new_n251));
  INV_X1    g0051(.A(G107), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n246), .A2(new_n247), .B1(new_n249), .B2(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT76), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT76), .A2(G33), .ZN(new_n256));
  OAI211_X1 g0056(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G68), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT76), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n242), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT76), .A2(G33), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT77), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n265), .B1(new_n260), .B2(G33), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n257), .B(new_n259), .C1(new_n264), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n254), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT68), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(new_n207), .B2(new_n242), .ZN(new_n270));
  NAND4_X1  g0070(.A1(KEYINPUT68), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(new_n220), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT69), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n270), .A2(KEYINPUT69), .A3(new_n220), .A4(new_n271), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n268), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G13), .A3(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n242), .A2(G1), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n274), .A2(G87), .A3(new_n275), .A4(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT15), .B(G87), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n280), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n277), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G1), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G1), .A3(G13), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(G250), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n288), .A2(G274), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT3), .B1(new_n255), .B2(new_n256), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n260), .A2(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT77), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G1698), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n298), .A2(G238), .A3(new_n299), .A4(new_n257), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n298), .A2(G244), .A3(G1698), .A4(new_n257), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n255), .A2(new_n256), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G116), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n291), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n294), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n286), .B1(G190), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n305), .ZN(new_n308));
  INV_X1    g0108(.A(new_n294), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G200), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n276), .ZN(new_n313));
  INV_X1    g0113(.A(new_n284), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(new_n282), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(new_n285), .A3(new_n277), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n308), .A2(G179), .A3(new_n309), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(new_n306), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT81), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n317), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n318), .B(KEYINPUT81), .C1(new_n319), .C2(new_n306), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n312), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(G20), .A2(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G150), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n243), .A2(new_n245), .ZN(new_n327));
  XOR2_X1   g0127(.A(KEYINPUT8), .B(G58), .Z(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OAI221_X1 g0129(.A(new_n326), .B1(new_n327), .B2(new_n329), .C1(new_n202), .C2(new_n221), .ZN(new_n330));
  INV_X1    g0130(.A(G50), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n330), .A2(new_n276), .B1(new_n331), .B2(new_n280), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n276), .B1(new_n278), .B2(G20), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G50), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT9), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT9), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n278), .B1(G41), .B2(G45), .ZN(new_n340));
  INV_X1    g0140(.A(G274), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n291), .A2(new_n340), .ZN(new_n344));
  INV_X1    g0144(.A(G226), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n242), .A2(KEYINPUT3), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n296), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT67), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n349), .A2(G223), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(G223), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n299), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(G222), .A2(G1698), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n296), .A2(new_n347), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n291), .B1(new_n355), .B2(new_n203), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n346), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G200), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(G190), .B2(new_n357), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n337), .A2(new_n339), .A3(new_n360), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n361), .B(KEYINPUT10), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n357), .A2(G169), .ZN(new_n363));
  INV_X1    g0163(.A(G179), .ZN(new_n364));
  AOI211_X1 g0164(.A(new_n363), .B(new_n336), .C1(new_n364), .C2(new_n357), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n333), .A2(G68), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n325), .A2(G50), .B1(G20), .B2(new_n258), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n327), .B2(new_n203), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n276), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT11), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n280), .A2(new_n258), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT12), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n276), .A2(KEYINPUT11), .A3(new_n370), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n368), .A2(new_n373), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n344), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n342), .B1(new_n378), .B2(G238), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT72), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n345), .A2(new_n299), .ZN(new_n381));
  INV_X1    g0181(.A(G232), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G1698), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n296), .A2(new_n381), .A3(new_n347), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n248), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n380), .B1(new_n385), .B2(new_n305), .ZN(new_n386));
  AOI211_X1 g0186(.A(KEYINPUT72), .B(new_n291), .C1(new_n384), .C2(new_n248), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n379), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT73), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT13), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT13), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n379), .B1(KEYINPUT73), .B2(new_n391), .C1(new_n386), .C2(new_n387), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(G179), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n388), .A2(KEYINPUT13), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n391), .B(new_n379), .C1(new_n386), .C2(new_n387), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n319), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  XOR2_X1   g0196(.A(KEYINPUT74), .B(KEYINPUT14), .Z(new_n397));
  OAI21_X1  g0197(.A(new_n393), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n394), .A2(new_n395), .ZN(new_n399));
  NAND2_X1  g0199(.A1(KEYINPUT74), .A2(KEYINPUT14), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n399), .A2(G169), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n377), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n377), .B1(new_n399), .B2(G200), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n390), .A2(G190), .A3(new_n392), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT75), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(new_n405), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT75), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n382), .A2(new_n299), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(G238), .B2(new_n299), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n291), .B1(new_n348), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n355), .A2(new_n252), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G244), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n343), .B1(new_n344), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G190), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n358), .B2(new_n417), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n279), .A2(G77), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT71), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n328), .A2(new_n325), .B1(G20), .B2(G77), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n284), .B2(new_n327), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n421), .B1(new_n423), .B2(new_n276), .ZN(new_n424));
  INV_X1    g0224(.A(new_n333), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(new_n203), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n417), .A2(new_n364), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n426), .B(new_n428), .C1(G169), .C2(new_n417), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NOR4_X1   g0230(.A1(new_n367), .A2(new_n406), .A3(new_n409), .A4(new_n430), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n298), .A2(new_n257), .ZN(new_n432));
  NOR2_X1   g0232(.A1(G223), .A2(G1698), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n345), .B2(G1698), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G87), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n305), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n342), .B1(new_n378), .B2(G232), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n358), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n291), .B1(new_n435), .B2(new_n436), .ZN(new_n441));
  INV_X1    g0241(.A(G190), .ZN(new_n442));
  INV_X1    g0242(.A(new_n439), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n425), .A2(new_n328), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n329), .A2(new_n279), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT16), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G58), .A2(G68), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n450), .B(KEYINPUT79), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(G58), .B2(G68), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n452), .A2(G20), .B1(G159), .B2(new_n325), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n298), .A2(new_n257), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT78), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT7), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n432), .B2(G20), .ZN(new_n459));
  AOI21_X1  g0259(.A(G20), .B1(new_n298), .B2(new_n257), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT78), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT7), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n457), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  AOI211_X1 g0263(.A(new_n449), .B(new_n454), .C1(new_n463), .C2(G68), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT3), .ZN(new_n465));
  INV_X1    g0265(.A(new_n347), .ZN(new_n466));
  OAI211_X1 g0266(.A(KEYINPUT7), .B(new_n221), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n458), .B1(new_n348), .B2(G20), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n453), .B1(new_n469), .B2(new_n258), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n313), .B1(new_n470), .B2(new_n449), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n445), .B(new_n448), .C1(new_n464), .C2(new_n472), .ZN(new_n473));
  OR2_X1    g0273(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n463), .A2(G68), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(KEYINPUT16), .A3(new_n453), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(new_n471), .B1(new_n446), .B2(new_n447), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n479), .A2(KEYINPUT80), .A3(KEYINPUT17), .A4(new_n445), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n441), .A2(new_n443), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(new_n319), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n441), .A2(new_n364), .A3(new_n443), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT18), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n479), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n448), .B1(new_n464), .B2(new_n472), .ZN(new_n487));
  INV_X1    g0287(.A(new_n483), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n319), .B2(new_n481), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT18), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n476), .B(new_n480), .C1(new_n486), .C2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n431), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT21), .ZN(new_n495));
  INV_X1    g0295(.A(G116), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n280), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(G20), .B1(G33), .B2(G283), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n242), .A2(G97), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n498), .A2(new_n499), .B1(G20), .B2(new_n496), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n272), .A2(KEYINPUT20), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT20), .B1(new_n272), .B2(new_n500), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n274), .A2(G116), .A3(new_n275), .A4(new_n282), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  MUX2_X1   g0306(.A(G257), .B(G264), .S(G1698), .Z(new_n507));
  OAI211_X1 g0307(.A(new_n257), .B(new_n507), .C1(new_n264), .C2(new_n266), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n355), .A2(G303), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n291), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g0310(.A(KEYINPUT5), .B(G41), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(G274), .A3(new_n288), .ZN(new_n512));
  INV_X1    g0312(.A(new_n511), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n291), .B1(new_n513), .B2(new_n289), .ZN(new_n514));
  INV_X1    g0314(.A(G270), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(G169), .B1(new_n510), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n495), .B1(new_n506), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n508), .A2(new_n509), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n305), .ZN(new_n520));
  INV_X1    g0320(.A(new_n512), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n305), .B1(new_n288), .B2(new_n511), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n521), .B1(new_n522), .B2(G270), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n504), .B(new_n497), .C1(new_n502), .C2(new_n501), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT21), .A4(G169), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n510), .A2(new_n516), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n527), .A3(G179), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n518), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(G257), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(new_n299), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n257), .B(new_n531), .C1(new_n264), .C2(new_n266), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT84), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n302), .A2(G294), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n298), .A2(G250), .A3(new_n299), .A4(new_n257), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT84), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n298), .A2(new_n536), .A3(new_n257), .A4(new_n531), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n533), .A2(new_n534), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n305), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n522), .A2(G264), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n539), .A2(new_n512), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT82), .B1(new_n252), .B2(G20), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT23), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT22), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n221), .A2(G87), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n355), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n545), .A2(new_n250), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n257), .B(new_n549), .C1(new_n264), .C2(new_n266), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n303), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n548), .B1(new_n551), .B2(new_n221), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT24), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT24), .ZN(new_n554));
  AOI21_X1  g0354(.A(G20), .B1(new_n550), .B2(new_n303), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n554), .B1(new_n555), .B2(new_n548), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n276), .A3(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n274), .A2(G107), .A3(new_n275), .A4(new_n282), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n279), .A2(G107), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n559), .B(KEYINPUT25), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT83), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT83), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n558), .A2(new_n563), .A3(new_n560), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n541), .A2(new_n364), .B1(new_n557), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n539), .A2(new_n512), .A3(new_n540), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n319), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n529), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n539), .A2(G190), .A3(new_n512), .A4(new_n540), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n570), .A2(new_n565), .A3(new_n557), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n538), .A2(new_n305), .B1(G264), .B2(new_n522), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n358), .B1(new_n572), .B2(new_n512), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n521), .B1(new_n522), .B2(G257), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n296), .A2(new_n347), .A3(G250), .A4(G1698), .ZN(new_n576));
  NAND2_X1  g0376(.A1(G33), .A2(G283), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT4), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n578), .A2(new_n415), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n299), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n576), .B(new_n577), .C1(new_n580), .C2(new_n355), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n298), .A2(G244), .A3(new_n299), .A4(new_n257), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(new_n582), .B2(new_n578), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n575), .B1(new_n583), .B2(new_n291), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G200), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n252), .B1(new_n467), .B2(new_n468), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT6), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n587), .A2(new_n251), .A3(G107), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n587), .B2(new_n239), .ZN(new_n589));
  INV_X1    g0389(.A(new_n325), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n589), .A2(new_n221), .B1(new_n203), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n276), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n274), .A2(G97), .A3(new_n275), .A4(new_n282), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n280), .A2(new_n251), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(G190), .B(new_n575), .C1(new_n583), .C2(new_n291), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n585), .A2(new_n592), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n592), .A2(new_n595), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n364), .B(new_n575), .C1(new_n583), .C2(new_n291), .ZN(new_n599));
  INV_X1    g0399(.A(new_n575), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n257), .B(G244), .C1(new_n264), .C2(new_n266), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n578), .B1(new_n601), .B2(G1698), .ZN(new_n602));
  INV_X1    g0402(.A(new_n581), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n600), .B1(new_n604), .B2(new_n305), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n598), .B(new_n599), .C1(new_n605), .C2(G169), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n527), .A2(G190), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n607), .B(new_n506), .C1(new_n358), .C2(new_n527), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n597), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n574), .A2(new_n609), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n324), .A2(new_n494), .A3(new_n569), .A4(new_n610), .ZN(G372));
  INV_X1    g0411(.A(KEYINPUT85), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n598), .B1(G200), .B2(new_n584), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n584), .A2(new_n319), .B1(new_n592), .B2(new_n595), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n613), .A2(new_n596), .B1(new_n614), .B2(new_n599), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n320), .A2(new_n316), .B1(new_n307), .B2(new_n311), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n567), .A2(G200), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(new_n565), .A3(new_n557), .A4(new_n570), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n612), .B1(new_n619), .B2(new_n569), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  INV_X1    g0421(.A(new_n606), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n616), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n320), .A2(new_n316), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n319), .B1(new_n308), .B2(new_n309), .ZN(new_n627));
  AOI211_X1 g0427(.A(new_n364), .B(new_n294), .C1(new_n304), .C2(new_n305), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n321), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(new_n323), .A3(new_n316), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n307), .A2(new_n311), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n631), .A3(new_n622), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT26), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n556), .A2(new_n276), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n555), .A2(new_n554), .A3(new_n548), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n565), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n572), .A2(new_n364), .A3(new_n512), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n568), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n518), .A2(new_n526), .A3(new_n528), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n640), .A2(new_n618), .A3(new_n615), .A4(new_n616), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n633), .B1(new_n641), .B2(new_n612), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n626), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n494), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n486), .A2(new_n490), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n476), .A2(new_n480), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n402), .A2(new_n429), .B1(new_n404), .B2(new_n403), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n362), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n366), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n644), .A2(new_n652), .ZN(G369));
  AND2_X1   g0453(.A1(new_n221), .A2(G13), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n278), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n557), .B2(new_n565), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n638), .B1(new_n574), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n638), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n661), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n639), .A2(new_n660), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(new_n665), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n525), .A2(new_n660), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n529), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n529), .A2(new_n670), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(new_n608), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G330), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n666), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n669), .A2(new_n676), .ZN(G399));
  AND2_X1   g0477(.A1(new_n643), .A2(new_n661), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n624), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n616), .A2(new_n622), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(KEYINPUT26), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n683), .B(new_n641), .C1(KEYINPUT26), .C2(new_n632), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n661), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT29), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n610), .A2(new_n324), .A3(new_n569), .A4(new_n661), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT31), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT86), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n520), .A2(new_n523), .A3(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n628), .A2(new_n572), .A3(new_n605), .A4(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n690), .A2(KEYINPUT86), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n527), .A2(new_n691), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(new_n584), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n628), .A3(new_n572), .A4(new_n694), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n527), .A2(G179), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n567), .A2(new_n310), .A3(new_n584), .A4(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n696), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n689), .B1(new_n702), .B2(new_n660), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n688), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n702), .A2(new_n660), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n674), .B1(new_n705), .B2(new_n689), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT87), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n704), .A2(new_n706), .A3(KEYINPUT87), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n687), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n278), .ZN(new_n713));
  INV_X1    g0513(.A(new_n208), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n253), .A2(G116), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G1), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n223), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n713), .A2(new_n720), .ZN(G364));
  NOR2_X1   g0521(.A1(new_n221), .A2(new_n442), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n364), .A2(G200), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n221), .A2(G190), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n723), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(G322), .A2(new_n725), .B1(new_n728), .B2(G311), .ZN(new_n729));
  INV_X1    g0529(.A(G303), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n358), .A2(G179), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n722), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n729), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n726), .A2(new_n731), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n348), .B(new_n733), .C1(G283), .C2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n364), .A2(new_n358), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n722), .ZN(new_n738));
  XNOR2_X1  g0538(.A(KEYINPUT91), .B(G326), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G179), .A2(G200), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n221), .B1(new_n740), .B2(G190), .ZN(new_n741));
  INV_X1    g0541(.A(G294), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n738), .A2(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT92), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT90), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n737), .A2(new_n745), .A3(new_n726), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n745), .B1(new_n737), .B2(new_n726), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(KEYINPUT33), .B(G317), .Z(new_n749));
  OAI211_X1 g0549(.A(new_n736), .B(new_n744), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n726), .A2(new_n740), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT89), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(KEYINPUT89), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT93), .Z(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n756), .A2(G329), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n738), .A2(new_n331), .B1(new_n734), .B2(new_n252), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n348), .B1(new_n741), .B2(new_n251), .C1(new_n203), .C2(new_n727), .ZN(new_n759));
  INV_X1    g0559(.A(new_n732), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n758), .B(new_n759), .C1(G87), .C2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G58), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n724), .B(KEYINPUT88), .Z(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n761), .B1(new_n762), .B2(new_n764), .C1(new_n258), .C2(new_n748), .ZN(new_n765));
  INV_X1    g0565(.A(new_n754), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G159), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT32), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n750), .A2(new_n757), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n220), .B1(G20), .B2(new_n319), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n278), .B1(new_n654), .B2(G45), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n715), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n348), .A2(G355), .A3(new_n208), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n237), .A2(new_n287), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n432), .A2(new_n714), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G45), .B2(new_n223), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n776), .B1(G116), .B2(new_n208), .C1(new_n777), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G13), .A2(G33), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n770), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n775), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n771), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(new_n673), .B2(new_n783), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n675), .A2(new_n774), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n673), .A2(new_n674), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(G396));
  NAND2_X1  g0591(.A1(new_n426), .A2(new_n660), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT94), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n427), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n792), .A2(new_n793), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n429), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n429), .A2(new_n660), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n711), .B(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n678), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n774), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n802), .B2(new_n801), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n355), .B1(new_n741), .B2(new_n251), .C1(new_n738), .C2(new_n730), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G107), .A2(new_n760), .B1(new_n725), .B2(G294), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n735), .A2(G87), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(new_n496), .C2(new_n727), .ZN(new_n808));
  INV_X1    g0608(.A(new_n748), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n805), .B(new_n808), .C1(G283), .C2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G311), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n811), .B2(new_n755), .ZN(new_n812));
  INV_X1    g0612(.A(new_n738), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n813), .A2(G137), .B1(new_n728), .B2(G159), .ZN(new_n814));
  INV_X1    g0614(.A(G150), .ZN(new_n815));
  INV_X1    g0615(.A(G143), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n814), .B1(new_n815), .B2(new_n748), .C1(new_n764), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n735), .A2(G68), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n331), .B2(new_n732), .ZN(new_n821));
  INV_X1    g0621(.A(new_n741), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n455), .B(new_n821), .C1(G58), .C2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G132), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n819), .B(new_n823), .C1(new_n824), .C2(new_n755), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n817), .A2(new_n818), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n812), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n770), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n770), .A2(new_n781), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n775), .B1(new_n203), .B2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n828), .B(new_n830), .C1(new_n800), .C2(new_n782), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n804), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G384));
  NAND2_X1  g0633(.A1(new_n377), .A2(new_n660), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n402), .A2(new_n405), .A3(new_n834), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n377), .B(new_n660), .C1(new_n398), .C2(new_n401), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n835), .A2(KEYINPUT96), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT96), .B1(new_n835), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n661), .B(new_n797), .C1(new_n626), .C2(new_n642), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n798), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT95), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT95), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n840), .A2(new_n843), .A3(new_n798), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n839), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n487), .A2(new_n489), .ZN(new_n846));
  INV_X1    g0646(.A(new_n658), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n487), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n846), .A2(new_n848), .A3(new_n849), .A4(new_n473), .ZN(new_n850));
  INV_X1    g0650(.A(new_n473), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n454), .B1(new_n463), .B2(G68), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n276), .B1(new_n852), .B2(KEYINPUT16), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT97), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(KEYINPUT97), .B(new_n276), .C1(new_n852), .C2(KEYINPUT16), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n478), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n448), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n484), .A2(new_n658), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n851), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n850), .B1(new_n860), .B2(new_n849), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT98), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n658), .B1(new_n857), .B2(new_n448), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n491), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n862), .B1(new_n491), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n861), .B(KEYINPUT38), .C1(new_n864), .C2(new_n865), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n845), .A2(new_n870), .B1(new_n645), .B2(new_n658), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n848), .A2(new_n846), .A3(new_n473), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n850), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n492), .B2(new_n848), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n867), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT39), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n869), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(KEYINPUT39), .B2(new_n870), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n402), .A2(new_n660), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n871), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n493), .B1(new_n680), .B2(new_n686), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n652), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n882), .B(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT40), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n869), .A2(new_n876), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n702), .A2(new_n660), .ZN(new_n889));
  NOR2_X1   g0689(.A1(KEYINPUT99), .A2(KEYINPUT31), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n890), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n702), .A2(new_n660), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n688), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n894), .B(new_n800), .C1(new_n837), .C2(new_n838), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n887), .B1(new_n888), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n887), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n868), .B2(new_n869), .ZN(new_n899));
  OAI21_X1  g0699(.A(G330), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n431), .A2(G330), .A3(new_n492), .A4(new_n894), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n494), .B(new_n894), .C1(new_n897), .C2(new_n899), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n886), .A2(new_n904), .B1(new_n278), .B2(new_n654), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n904), .B2(new_n886), .ZN(new_n906));
  INV_X1    g0706(.A(new_n589), .ZN(new_n907));
  OAI211_X1 g0707(.A(G116), .B(new_n222), .C1(new_n907), .C2(KEYINPUT35), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(KEYINPUT35), .B2(new_n907), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT36), .ZN(new_n910));
  INV_X1    g0710(.A(new_n201), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(G68), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n451), .A2(G77), .A3(new_n224), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n278), .B(G13), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  OR3_X1    g0714(.A1(new_n906), .A2(new_n910), .A3(new_n914), .ZN(G367));
  NAND2_X1  g0715(.A1(new_n286), .A2(new_n660), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT100), .B1(new_n616), .B2(new_n916), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n624), .A2(new_n916), .ZN(new_n918));
  MUX2_X1   g0718(.A(KEYINPUT100), .B(new_n917), .S(new_n918), .Z(new_n919));
  XNOR2_X1  g0719(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n622), .A2(new_n660), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n922), .A2(KEYINPUT103), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n598), .A2(new_n660), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n615), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n922), .A2(KEYINPUT103), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n666), .A2(new_n927), .A3(new_n675), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT102), .Z(new_n929));
  AND2_X1   g0729(.A1(new_n927), .A2(new_n664), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n661), .B1(new_n930), .B2(new_n622), .ZN(new_n931));
  INV_X1    g0731(.A(new_n668), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n927), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT42), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT104), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n936), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n934), .A2(new_n935), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT105), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n938), .A2(KEYINPUT105), .A3(new_n939), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT43), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n919), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n929), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n929), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n946), .B(new_n949), .C1(new_n942), .C2(new_n943), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n921), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n943), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT105), .B1(new_n938), .B2(new_n939), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n947), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n949), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n944), .A2(new_n947), .A3(new_n929), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n955), .A2(new_n956), .A3(new_n919), .A4(new_n920), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n669), .A2(new_n927), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT45), .Z(new_n959));
  NOR2_X1   g0759(.A1(new_n669), .A2(new_n927), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT44), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(new_n676), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n666), .A2(new_n667), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(KEYINPUT106), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(new_n675), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(new_n668), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n712), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n712), .B1(new_n963), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n715), .B(KEYINPUT41), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n772), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n951), .A2(new_n957), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n919), .A2(new_n783), .ZN(new_n974));
  INV_X1    g0774(.A(new_n770), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n809), .A2(G159), .B1(new_n201), .B2(new_n728), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT109), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(KEYINPUT109), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n766), .A2(G137), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n738), .A2(new_n816), .B1(new_n724), .B2(new_n815), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n348), .B1(new_n741), .B2(new_n258), .C1(new_n203), .C2(new_n734), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n980), .B(new_n981), .C1(G58), .C2(new_n760), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n977), .A2(new_n978), .A3(new_n979), .A4(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(KEYINPUT107), .B(G317), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n766), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n735), .A2(G97), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n985), .A2(new_n455), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT108), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(G283), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n738), .A2(new_n811), .B1(new_n727), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n732), .A2(new_n496), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT46), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n991), .B(new_n993), .C1(G107), .C2(new_n822), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n763), .A2(G303), .B1(new_n809), .B2(G294), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n989), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n987), .A2(new_n988), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n983), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT47), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n975), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n999), .B2(new_n998), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n778), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n784), .B1(new_n208), .B2(new_n284), .C1(new_n1002), .C2(new_n232), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n974), .A2(new_n774), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n973), .A2(new_n1004), .ZN(G387));
  AND2_X1   g0805(.A1(new_n712), .A2(new_n967), .ZN(new_n1006));
  OR3_X1    g0806(.A1(new_n1006), .A2(new_n968), .A3(new_n716), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n783), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n666), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n784), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n229), .A2(G45), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n348), .A2(new_n208), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1011), .A2(new_n1002), .B1(new_n717), .B2(new_n1012), .ZN(new_n1013));
  OR3_X1    g0813(.A1(new_n329), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1014));
  OAI21_X1  g0814(.A(KEYINPUT50), .B1(new_n329), .B2(G50), .ZN(new_n1015));
  AOI21_X1  g0815(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1014), .A2(new_n717), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n1013), .A2(new_n1017), .B1(new_n252), .B2(new_n714), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n432), .B1(new_n329), .B2(new_n748), .C1(new_n754), .C2(new_n815), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n813), .A2(G159), .B1(new_n728), .B2(G68), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n203), .B2(new_n732), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n986), .B1(new_n331), .B2(new_n724), .C1(new_n284), .C2(new_n741), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n813), .A2(G322), .B1(new_n728), .B2(G303), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n811), .B2(new_n748), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n763), .B2(new_n984), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT48), .Z(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n990), .B2(new_n741), .C1(new_n742), .C2(new_n732), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT49), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n455), .B1(new_n496), .B2(new_n734), .C1(new_n754), .C2(new_n739), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1023), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n774), .B1(new_n1010), .B2(new_n1018), .C1(new_n1033), .C2(new_n975), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT110), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1007), .B1(new_n772), .B2(new_n967), .C1(new_n1009), .C2(new_n1035), .ZN(G393));
  AOI21_X1  g0836(.A(new_n716), .B1(new_n963), .B2(new_n968), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n963), .B2(new_n968), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n927), .A2(new_n1008), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(KEYINPUT111), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(KEYINPUT111), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n778), .A2(new_n240), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n784), .B1(new_n251), .B2(new_n208), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n348), .B1(new_n735), .B2(G107), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n990), .B2(new_n732), .C1(new_n742), .C2(new_n727), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT52), .ZN(new_n1046));
  INV_X1    g0846(.A(G317), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n738), .A2(new_n1047), .B1(new_n724), .B2(new_n811), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n766), .A2(G322), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n1046), .B2(new_n1048), .C1(new_n730), .C2(new_n748), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1045), .B(new_n1050), .C1(G116), .C2(new_n822), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n754), .A2(new_n816), .B1(new_n258), .B2(new_n732), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT112), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1054), .A2(new_n432), .A3(new_n807), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT113), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(G159), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n738), .A2(new_n815), .B1(new_n724), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT51), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n728), .A2(new_n328), .B1(new_n822), .B2(G77), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n911), .C2(new_n748), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1051), .B1(new_n1058), .B2(new_n1064), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n774), .B1(new_n1042), .B2(new_n1043), .C1(new_n1065), .C2(new_n975), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1041), .A2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n963), .A2(new_n773), .B1(new_n1040), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1038), .A2(new_n1068), .ZN(G390));
  AOI21_X1  g0869(.A(new_n799), .B1(new_n709), .B2(new_n710), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n838), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n835), .A2(KEYINPUT96), .A3(new_n836), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n797), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n798), .B1(new_n685), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n880), .B1(new_n1076), .B2(new_n1073), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n888), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n491), .A2(new_n863), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(KEYINPUT98), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n491), .A2(new_n862), .A3(new_n863), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(KEYINPUT38), .B1(new_n1082), .B2(new_n861), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n869), .ZN(new_n1084));
  OAI21_X1  g0884(.A(KEYINPUT39), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n869), .A2(new_n876), .A3(new_n877), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n845), .A2(new_n880), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1074), .B(new_n1078), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1078), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n844), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n843), .B1(new_n840), .B2(new_n798), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1073), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n881), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1090), .B1(new_n879), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(KEYINPUT114), .B1(new_n895), .B2(new_n674), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n893), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n892), .B1(new_n702), .B2(new_n660), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n799), .B1(new_n1099), .B2(new_n688), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT114), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1100), .A2(new_n1073), .A3(new_n1101), .A4(G330), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1096), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1089), .B1(new_n1095), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(KEYINPUT119), .B1(new_n1105), .B2(new_n772), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1085), .B(new_n1086), .C1(new_n880), .C2(new_n845), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1104), .B1(new_n1107), .B2(new_n1078), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT119), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1109), .A2(new_n1110), .A3(new_n773), .A4(new_n1089), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n829), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1113), .A2(new_n328), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n756), .A2(G125), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n732), .A2(new_n815), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT53), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n355), .B(new_n1118), .C1(G132), .C2(new_n725), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n809), .A2(G137), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1116), .A2(new_n1117), .B1(G159), .B2(new_n822), .ZN(new_n1121));
  INV_X1    g0921(.A(G128), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n911), .A2(new_n734), .B1(new_n1122), .B2(new_n738), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT54), .B(G143), .Z(new_n1124));
  AOI21_X1  g0924(.A(new_n1123), .B1(new_n728), .B2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1125), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n820), .B1(new_n251), .B2(new_n727), .C1(new_n990), .C2(new_n738), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n348), .B(new_n1127), .C1(G87), .C2(new_n760), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n724), .A2(new_n496), .B1(new_n741), .B2(new_n203), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT120), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1128), .B(new_n1130), .C1(new_n252), .C2(new_n748), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n755), .A2(new_n742), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1115), .A2(new_n1126), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n775), .B(new_n1114), .C1(new_n1133), .C2(new_n770), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n1087), .B2(new_n782), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1112), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1100), .A2(G330), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1076), .B1(new_n1137), .B2(new_n839), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1074), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n842), .A2(new_n844), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1073), .B1(new_n711), .B2(new_n800), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(new_n1142), .B2(new_n1103), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT116), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1102), .B(new_n1096), .C1(new_n1070), .C2(new_n1073), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT116), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n1146), .A3(new_n1141), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1140), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n901), .A2(KEYINPUT115), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n901), .A2(KEYINPUT115), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n884), .A2(new_n652), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(KEYINPUT117), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1145), .A2(new_n1146), .A3(new_n1141), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1146), .B1(new_n1145), .B2(new_n1141), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1139), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1150), .A2(new_n1149), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1156), .A2(new_n883), .A3(new_n651), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT117), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1152), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT118), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1152), .A2(KEYINPUT118), .A3(new_n1159), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n1105), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1105), .B1(new_n1152), .B2(new_n1159), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1165), .A2(new_n716), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1136), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(G378));
  OAI21_X1  g0968(.A(new_n774), .B1(new_n1113), .B2(new_n201), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT123), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n336), .A2(new_n658), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n367), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n367), .A2(new_n1173), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1172), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1174), .A2(new_n1175), .A3(new_n1172), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1170), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1178), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(KEYINPUT123), .A3(new_n1176), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1182), .A2(new_n782), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n735), .A2(G58), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT121), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G97), .B2(new_n809), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n432), .A2(G41), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n724), .A2(new_n252), .B1(new_n727), .B2(new_n284), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n738), .A2(new_n496), .B1(new_n732), .B2(new_n203), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(G68), .C2(new_n822), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1186), .A2(new_n1187), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G283), .B2(new_n756), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT122), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1193), .A2(KEYINPUT58), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(KEYINPUT58), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(G33), .A2(G41), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1187), .A2(G50), .A3(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G125), .A2(new_n813), .B1(new_n725), .B2(G128), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n760), .A2(new_n1124), .B1(new_n728), .B2(G137), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n824), .B2(new_n748), .C1(new_n815), .C2(new_n741), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1202));
  INV_X1    g1002(.A(G124), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1196), .B1(new_n1059), .B2(new_n734), .C1(new_n754), .C2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1201), .B2(KEYINPUT59), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1197), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1194), .A2(new_n1195), .A3(new_n1206), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1169), .B(new_n1183), .C1(new_n770), .C2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n900), .A2(new_n1180), .A3(new_n1176), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1182), .B(G330), .C1(new_n897), .C2(new_n899), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1209), .A2(new_n882), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n882), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1208), .B1(new_n1213), .B2(new_n773), .ZN(new_n1214));
  OAI211_X1 g1014(.A(KEYINPUT57), .B(new_n1213), .C1(new_n1165), .C2(new_n1151), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n715), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1074), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1217), .B(new_n1090), .C1(new_n879), .C2(new_n1094), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1218), .A2(new_n1108), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1148), .A2(KEYINPUT117), .A3(new_n1151), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1158), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1219), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1157), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT57), .B1(new_n1223), .B2(new_n1213), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1214), .B1(new_n1216), .B2(new_n1224), .ZN(G375));
  NAND2_X1  g1025(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1162), .A2(new_n970), .A3(new_n1163), .A4(new_n1226), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT124), .Z(new_n1228));
  AOI21_X1  g1028(.A(new_n775), .B1(new_n258), .B2(new_n829), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n809), .A2(new_n1124), .ZN(new_n1230));
  INV_X1    g1030(.A(G137), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1230), .B1(new_n764), .B2(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G132), .A2(new_n813), .B1(new_n760), .B2(G159), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n331), .B2(new_n741), .C1(new_n815), .C2(new_n727), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(new_n1232), .A2(new_n1234), .A3(new_n455), .A4(new_n1185), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n756), .A2(G128), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n756), .A2(G303), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n748), .A2(new_n496), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n355), .B1(new_n741), .B2(new_n284), .C1(new_n203), .C2(new_n734), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n738), .A2(new_n742), .B1(new_n724), .B2(new_n990), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n732), .A2(new_n251), .B1(new_n727), .B2(new_n252), .ZN(new_n1241));
  NOR4_X1   g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1235), .A2(new_n1236), .B1(new_n1237), .B2(new_n1242), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1229), .B1(new_n975), .B2(new_n1243), .C1(new_n1073), .C2(new_n782), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1148), .B2(new_n772), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1228), .A2(new_n1246), .ZN(G381));
  INV_X1    g1047(.A(G375), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1167), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1038), .A2(new_n832), .A3(new_n1068), .ZN(new_n1251));
  NOR4_X1   g1051(.A1(G387), .A2(G396), .A3(G393), .A4(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1250), .A2(new_n1228), .A3(new_n1246), .A4(new_n1252), .ZN(G407));
  OAI211_X1 g1053(.A(G407), .B(G213), .C1(G343), .C2(new_n1249), .ZN(G409));
  AND3_X1   g1054(.A1(new_n973), .A2(new_n1004), .A3(G390), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G390), .B1(new_n973), .B2(new_n1004), .ZN(new_n1256));
  OAI21_X1  g1056(.A(KEYINPUT126), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(G393), .B(new_n790), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1257), .B(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(KEYINPUT61), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1213), .B1(new_n1165), .B2(new_n1151), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT57), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n715), .A3(new_n1215), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1167), .B1(new_n1264), .B2(new_n1214), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1136), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1223), .A2(new_n970), .A3(new_n1213), .ZN(new_n1268));
  AND4_X1   g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1214), .A4(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n659), .A2(G213), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1265), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT60), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1226), .B1(new_n1160), .B2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1226), .A2(new_n1273), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1275), .A2(new_n716), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1277), .B2(new_n1246), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n832), .B(new_n1245), .C1(new_n1274), .C2(new_n1276), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1272), .A2(KEYINPUT63), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT125), .B1(new_n1265), .B2(new_n1269), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G375), .A2(G378), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT125), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1167), .A2(new_n1214), .A3(new_n1268), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1284), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1283), .A2(new_n1287), .A3(new_n1270), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1271), .A2(G2897), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1280), .B(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1282), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1280), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1288), .A2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1260), .B(new_n1281), .C1(new_n1291), .C2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1284), .A2(new_n1286), .A3(new_n1270), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1290), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1272), .A2(KEYINPUT127), .A3(KEYINPUT62), .A4(new_n1280), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT127), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1284), .A2(new_n1280), .A3(new_n1286), .A4(new_n1270), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1300), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1299), .A2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1302), .B1(new_n1288), .B2(new_n1292), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1298), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1258), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1257), .B(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1294), .B1(new_n1306), .B2(new_n1308), .ZN(G405));
  OAI21_X1  g1109(.A(new_n1308), .B1(new_n1250), .B2(new_n1265), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1259), .A2(new_n1249), .A3(new_n1284), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1310), .A2(new_n1311), .A3(new_n1280), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1280), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(G402));
endmodule


