//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993, new_n994, new_n995;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g002(.A1(G127gat), .A2(G134gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(KEYINPUT68), .B(G127gat), .Z(new_n206));
  INV_X1    g005(.A(G134gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G113gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(G113gat), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT1), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(KEYINPUT69), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT69), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G120gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n218), .A3(G113gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT70), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n219), .A2(new_n220), .A3(new_n211), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n220), .B1(new_n219), .B2(new_n211), .ZN(new_n222));
  NAND2_X1  g021(.A1(G127gat), .A2(G134gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(KEYINPUT71), .A2(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g024(.A1(KEYINPUT71), .A2(KEYINPUT1), .ZN(new_n226));
  OAI22_X1  g025(.A1(new_n224), .A2(new_n204), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NOR4_X1   g026(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT72), .A4(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT72), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n219), .A2(new_n211), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n227), .B1(new_n230), .B2(KEYINPUT70), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT69), .B(G120gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n210), .B1(new_n232), .B2(G113gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n220), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n229), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n215), .B1(new_n228), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n237));
  XOR2_X1   g036(.A(G141gat), .B(G148gat), .Z(new_n238));
  INV_X1    g037(.A(G155gat), .ZN(new_n239));
  INV_X1    g038(.A(G162gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G155gat), .A2(G162gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(KEYINPUT2), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n238), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G141gat), .B(G148gat), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n242), .B(new_n241), .C1(new_n246), .C2(KEYINPUT2), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n237), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n247), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT79), .B1(new_n249), .B2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT79), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n245), .A2(new_n247), .A3(new_n251), .A4(new_n237), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n248), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n203), .B1(new_n236), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n249), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n255), .B(new_n215), .C1(new_n228), .C2(new_n235), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n227), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n233), .B2(new_n220), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT72), .B1(new_n260), .B2(new_n221), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n231), .A2(new_n229), .A3(new_n234), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n263), .A2(KEYINPUT4), .A3(new_n255), .A4(new_n215), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n254), .A2(new_n258), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT80), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT80), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n254), .A2(new_n258), .A3(new_n264), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n255), .B1(new_n263), .B2(new_n215), .ZN(new_n270));
  AOI211_X1 g069(.A(new_n249), .B(new_n214), .C1(new_n261), .C2(new_n262), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n203), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n265), .A2(KEYINPUT5), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G1gat), .B(G29gat), .Z(new_n278));
  XNOR2_X1  g077(.A(G57gat), .B(G85gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n280), .B(new_n281), .Z(new_n282));
  NAND3_X1  g081(.A1(new_n275), .A2(new_n277), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n284));
  INV_X1    g083(.A(new_n282), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n273), .B1(new_n266), .B2(new_n268), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n285), .B1(new_n286), .B2(new_n276), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n283), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(KEYINPUT6), .B(new_n285), .C1(new_n286), .C2(new_n276), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G226gat), .A2(G233gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT24), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(G183gat), .A3(G190gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G183gat), .B(G190gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n295), .B1(new_n296), .B2(new_n294), .ZN(new_n297));
  NOR2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT23), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT23), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(G169gat), .B2(G176gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n299), .A2(KEYINPUT25), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G183gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G183gat), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n294), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n295), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT66), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT66), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n312), .B(new_n295), .C1(new_n296), .C2(new_n294), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n299), .A2(new_n302), .A3(new_n301), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT65), .B(KEYINPUT25), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n304), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT26), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(new_n298), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n298), .A2(KEYINPUT26), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(new_n305), .B2(new_n307), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT27), .B(G183gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n307), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT28), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(KEYINPUT67), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(KEYINPUT67), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n324), .A2(new_n307), .A3(new_n328), .ZN(new_n329));
  AOI211_X1 g128(.A(new_n321), .B(new_n323), .C1(new_n327), .C2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n293), .B1(new_n318), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n329), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n323), .A2(new_n321), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n317), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n314), .B1(new_n297), .B2(KEYINPUT66), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(new_n313), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n334), .B(new_n291), .C1(new_n337), .C2(new_n304), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n331), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G197gat), .B(G204gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT22), .ZN(new_n341));
  INV_X1    g140(.A(G211gat), .ZN(new_n342));
  INV_X1    g141(.A(G218gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G211gat), .B(G218gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n340), .A3(new_n344), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n339), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT91), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT91), .A3(new_n351), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n331), .A2(new_n338), .A3(new_n350), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT90), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT90), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n331), .A2(new_n338), .A3(new_n358), .A4(new_n350), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n354), .A2(new_n355), .A3(new_n357), .A4(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT38), .B1(new_n360), .B2(KEYINPUT37), .ZN(new_n361));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n352), .A2(new_n365), .A3(new_n356), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n331), .A2(new_n338), .A3(KEYINPUT76), .A4(new_n350), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT37), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n364), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT92), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n361), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(new_n361), .B2(new_n370), .ZN(new_n373));
  INV_X1    g172(.A(new_n364), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n374), .B1(new_n366), .B2(new_n367), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n290), .A2(new_n376), .A3(KEYINPUT93), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT93), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n370), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT92), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n370), .A3(new_n371), .ZN(new_n381));
  INV_X1    g180(.A(new_n375), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n288), .A2(new_n289), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n378), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n370), .B1(new_n369), .B2(new_n368), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT38), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n377), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n250), .A2(new_n252), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n350), .B1(new_n389), .B2(new_n292), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT29), .B1(new_n348), .B2(new_n349), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(KEYINPUT3), .ZN(new_n392));
  OAI211_X1 g191(.A(G228gat), .B(G233gat), .C1(new_n392), .C2(new_n255), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT85), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n350), .A2(new_n292), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n237), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n397), .B2(new_n249), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT29), .B1(new_n250), .B2(new_n252), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n398), .B(new_n399), .C1(new_n350), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n394), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n237), .B1(new_n391), .B2(KEYINPUT84), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n350), .A2(KEYINPUT84), .A3(new_n292), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n249), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n350), .B2(new_n400), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n395), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT86), .B(G22gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(G78gat), .B(G106gat), .Z(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT31), .B(G50gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n413), .B(KEYINPUT83), .Z(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n413), .B1(new_n408), .B2(G22gat), .ZN(new_n417));
  AND4_X1   g216(.A1(KEYINPUT87), .A2(new_n402), .A3(new_n407), .A4(new_n409), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n394), .A2(new_n401), .B1(new_n406), .B2(new_n395), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT87), .B1(new_n419), .B2(new_n409), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n417), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n417), .B(KEYINPUT88), .C1(new_n418), .C2(new_n420), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n416), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n368), .A2(KEYINPUT30), .A3(new_n364), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT77), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n366), .A2(new_n367), .A3(new_n374), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  XOR2_X1   g229(.A(KEYINPUT78), .B(KEYINPUT30), .Z(new_n431));
  NOR2_X1   g230(.A1(new_n375), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n428), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT40), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n236), .A2(new_n253), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n258), .A2(new_n264), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n203), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n236), .A2(new_n249), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(new_n256), .A3(new_n202), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n438), .A2(KEYINPUT39), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT39), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n437), .A2(new_n442), .A3(new_n203), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n282), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n435), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n438), .A2(KEYINPUT39), .A3(new_n440), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n446), .A2(KEYINPUT40), .A3(new_n282), .A4(new_n443), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n287), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n449), .A3(KEYINPUT89), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n452));
  OAI22_X1  g251(.A1(new_n452), .A2(new_n432), .B1(new_n427), .B2(new_n426), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n451), .B1(new_n453), .B2(new_n448), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n425), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n388), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT36), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n318), .A2(new_n330), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n236), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n263), .B(new_n215), .C1(new_n318), .C2(new_n330), .ZN(new_n460));
  NAND2_X1  g259(.A1(G227gat), .A2(G233gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(KEYINPUT64), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT32), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT73), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(KEYINPUT73), .A3(KEYINPUT32), .ZN(new_n467));
  XNOR2_X1  g266(.A(G15gat), .B(G43gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(G71gat), .B(G99gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT33), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n470), .B1(new_n463), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n466), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n463), .B(KEYINPUT32), .C1(new_n471), .C2(new_n470), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT75), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(KEYINPUT75), .A3(new_n474), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n459), .A2(new_n460), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n479), .A2(KEYINPUT34), .A3(new_n462), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT74), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n459), .A2(new_n460), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT74), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n461), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n480), .B1(new_n485), .B2(KEYINPUT34), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n477), .A2(new_n478), .A3(new_n486), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n475), .A2(new_n486), .A3(new_n476), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n457), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OR3_X1    g288(.A1(new_n475), .A2(new_n486), .A3(new_n476), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n477), .A2(new_n478), .A3(new_n486), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT36), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT82), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n384), .A2(new_n494), .A3(new_n453), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n384), .B2(new_n453), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n493), .B1(new_n497), .B2(new_n425), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n423), .A2(new_n424), .ZN(new_n499));
  INV_X1    g298(.A(new_n416), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n490), .A2(new_n491), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n495), .B2(new_n496), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n290), .A2(KEYINPUT35), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n501), .A2(new_n504), .A3(new_n453), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n456), .A2(new_n498), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT94), .ZN(new_n507));
  XOR2_X1   g306(.A(G15gat), .B(G22gat), .Z(new_n508));
  INV_X1    g307(.A(G1gat), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT16), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(G1gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n514), .A2(G8gat), .ZN(new_n515));
  INV_X1    g314(.A(G8gat), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n510), .B2(new_n513), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G29gat), .ZN(new_n519));
  INV_X1    g318(.A(G36gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT14), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT14), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(G29gat), .A2(G36gat), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n521), .A2(new_n523), .A3(KEYINPUT15), .A4(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G43gat), .B(G50gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT15), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n525), .A2(new_n526), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n528), .B(new_n529), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n525), .A2(new_n526), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n532), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n529), .B1(new_n538), .B2(new_n528), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n518), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n514), .B(G8gat), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n527), .B1(new_n537), .B2(new_n532), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT18), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(G197gat), .ZN(new_n550));
  XOR2_X1   g349(.A(KEYINPUT11), .B(G169gat), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT12), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n540), .A2(new_n545), .A3(KEYINPUT18), .A4(new_n541), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n541), .B(KEYINPUT13), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n518), .A2(new_n543), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n518), .A2(new_n543), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n548), .A2(new_n553), .A3(new_n554), .A4(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n556), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n546), .A2(new_n547), .B1(new_n562), .B2(new_n555), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n553), .B1(new_n563), .B2(new_n554), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT95), .B1(new_n506), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n567));
  INV_X1    g366(.A(new_n564), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n560), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n499), .A2(new_n500), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT89), .B1(new_n434), .B2(new_n449), .ZN(new_n571));
  NOR3_X1   g370(.A1(new_n453), .A2(new_n448), .A3(new_n451), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n373), .A2(new_n375), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n574), .A2(new_n289), .A3(new_n288), .A4(new_n381), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n575), .A2(new_n378), .B1(KEYINPUT38), .B2(new_n386), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n573), .B1(new_n377), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n489), .A2(new_n492), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n384), .A2(new_n453), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT82), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n384), .A2(new_n494), .A3(new_n453), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n425), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n501), .A2(new_n453), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n586), .A2(new_n504), .B1(new_n502), .B2(KEYINPUT35), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n567), .B(new_n569), .C1(new_n584), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n566), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(new_n384), .ZN(new_n591));
  XNOR2_X1  g390(.A(G57gat), .B(G64gat), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OR2_X1    g393(.A1(G71gat), .A2(G78gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(G71gat), .A2(G78gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT96), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n595), .A2(KEYINPUT96), .A3(new_n596), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n594), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n597), .B(new_n598), .C1(new_n592), .C2(new_n593), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n542), .B1(KEYINPUT21), .B2(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n601), .A2(new_n602), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(G127gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n608), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n610), .B1(new_n609), .B2(new_n611), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n604), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n614), .ZN(new_n616));
  INV_X1    g415(.A(new_n604), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n617), .A3(new_n612), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT97), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G155gat), .ZN(new_n621));
  XOR2_X1   g420(.A(G183gat), .B(G211gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n615), .A2(new_n618), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n623), .B1(new_n615), .B2(new_n618), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(G85gat), .A2(G92gat), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT7), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(KEYINPUT98), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G99gat), .A2(G106gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT8), .ZN(new_n632));
  INV_X1    g431(.A(G85gat), .ZN(new_n633));
  INV_X1    g432(.A(G92gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n630), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n637));
  OR2_X1    g436(.A1(G99gat), .A2(G106gat), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n638), .B2(new_n631), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n637), .A3(new_n631), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT98), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT7), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n629), .A2(KEYINPUT98), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n643), .A2(new_n644), .A3(G85gat), .A4(G92gat), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n636), .A2(new_n640), .A3(new_n641), .A4(new_n645), .ZN(new_n646));
  AND4_X1   g445(.A1(G85gat), .A2(new_n643), .A3(new_n644), .A4(G92gat), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n630), .A2(new_n632), .A3(new_n635), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n638), .A2(new_n637), .A3(new_n631), .ZN(new_n649));
  OAI22_X1  g448(.A1(new_n647), .A2(new_n648), .B1(new_n649), .B2(new_n639), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n627), .B1(new_n651), .B2(new_n543), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(KEYINPUT100), .B(new_n627), .C1(new_n651), .C2(new_n543), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n651), .B1(new_n536), .B2(new_n539), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(G190gat), .B(G218gat), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n659), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n656), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(G134gat), .B(G162gat), .Z(new_n664));
  AOI21_X1  g463(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(KEYINPUT101), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n666), .A2(KEYINPUT101), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n660), .A2(new_n669), .A3(new_n662), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n605), .A2(new_n651), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT10), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n603), .A2(new_n646), .A3(new_n650), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n603), .A2(KEYINPUT10), .A3(new_n646), .A4(new_n650), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(G230gat), .A2(G233gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(G120gat), .B(G148gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(G176gat), .B(G204gat), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n680), .B(new_n681), .Z(new_n682));
  AND2_X1   g481(.A1(new_n672), .A2(new_n674), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n679), .B(new_n682), .C1(new_n683), .C2(new_n678), .ZN(new_n684));
  INV_X1    g483(.A(new_n682), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n683), .A2(new_n678), .ZN(new_n686));
  INV_X1    g485(.A(new_n678), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n675), .B2(new_n676), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n685), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n626), .A2(new_n671), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n591), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g494(.A(new_n453), .B1(new_n566), .B2(new_n588), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT16), .B(G8gat), .Z(new_n697));
  NAND4_X1  g496(.A1(new_n696), .A2(KEYINPUT42), .A3(new_n693), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT103), .ZN(new_n699));
  AOI211_X1 g498(.A(new_n692), .B(new_n453), .C1(new_n566), .C2(new_n588), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n700), .A2(new_n701), .A3(KEYINPUT42), .A4(new_n697), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n700), .A2(new_n516), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n696), .A2(new_n693), .A3(new_n697), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n706), .A2(new_n705), .A3(new_n707), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n703), .B(new_n704), .C1(new_n708), .C2(new_n709), .ZN(G1325gat));
  INV_X1    g509(.A(G15gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n490), .A2(new_n491), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n589), .A2(new_n711), .A3(new_n693), .A4(new_n712), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n590), .A2(new_n692), .A3(new_n578), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(new_n711), .ZN(G1326gat));
  NAND3_X1  g514(.A1(new_n589), .A2(new_n693), .A3(new_n425), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n589), .A2(KEYINPUT104), .A3(new_n693), .A4(new_n425), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT43), .B(G22gat), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n718), .B2(new_n719), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(G1327gat));
  NOR2_X1   g522(.A1(new_n626), .A2(new_n690), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n660), .A2(new_n669), .A3(new_n662), .ZN(new_n725));
  INV_X1    g524(.A(new_n667), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n726), .B1(new_n660), .B2(new_n662), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n591), .A2(new_n519), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n591), .A2(KEYINPUT45), .A3(new_n519), .A4(new_n730), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(new_n506), .B2(new_n671), .ZN(new_n736));
  OAI211_X1 g535(.A(KEYINPUT44), .B(new_n728), .C1(new_n584), .C2(new_n587), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n626), .A2(new_n690), .A3(new_n565), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G29gat), .B1(new_n740), .B2(new_n384), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n733), .A2(new_n734), .A3(new_n741), .ZN(G1328gat));
  NAND3_X1  g541(.A1(new_n696), .A2(new_n520), .A3(new_n730), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n743), .A2(KEYINPUT46), .ZN(new_n744));
  OAI21_X1  g543(.A(G36gat), .B1(new_n740), .B2(new_n453), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(KEYINPUT46), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(G1329gat));
  NAND4_X1  g546(.A1(new_n736), .A2(new_n737), .A3(new_n493), .A4(new_n739), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G43gat), .ZN(new_n749));
  INV_X1    g548(.A(G43gat), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n730), .A2(new_n750), .A3(new_n712), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n590), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1330gat));
  NAND4_X1  g553(.A1(new_n736), .A2(new_n737), .A3(new_n425), .A4(new_n739), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G50gat), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n570), .A2(G50gat), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT105), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n730), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n756), .B1(new_n590), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT48), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1331gat));
  NAND3_X1  g563(.A1(new_n626), .A2(new_n671), .A3(new_n690), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n506), .A2(new_n569), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n290), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n434), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT49), .B(G64gat), .Z(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n769), .B2(new_n771), .ZN(G1333gat));
  XOR2_X1   g571(.A(new_n712), .B(KEYINPUT106), .Z(new_n773));
  AOI21_X1  g572(.A(G71gat), .B1(new_n766), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n493), .A2(G71gat), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n774), .B1(new_n766), .B2(new_n775), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n776), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g576(.A1(new_n766), .A2(new_n425), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g578(.A1(new_n626), .A2(new_n569), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n691), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n738), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783), .B2(new_n384), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n456), .A2(new_n582), .A3(new_n578), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n570), .A2(new_n712), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n580), .B2(new_n581), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT35), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n505), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n671), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT51), .B1(new_n790), .B2(new_n780), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(KEYINPUT51), .A3(new_n780), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(KEYINPUT107), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n290), .A2(new_n633), .A3(new_n690), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n784), .B1(new_n797), .B2(new_n798), .ZN(G1336gat));
  XOR2_X1   g598(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n800));
  NAND4_X1  g599(.A1(new_n736), .A2(new_n737), .A3(new_n434), .A4(new_n782), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n801), .B2(G92gat), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n434), .A2(new_n634), .A3(new_n690), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n801), .A2(KEYINPUT108), .A3(G92gat), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT108), .B1(new_n801), .B2(G92gat), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n803), .B1(new_n792), .B2(new_n793), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n804), .B1(new_n808), .B2(new_n809), .ZN(G1337gat));
  NOR2_X1   g609(.A1(new_n783), .A2(new_n578), .ZN(new_n811));
  XNOR2_X1  g610(.A(KEYINPUT110), .B(G99gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n712), .A2(new_n690), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT111), .ZN(new_n814));
  OAI22_X1  g613(.A1(new_n811), .A2(new_n812), .B1(new_n797), .B2(new_n814), .ZN(G1338gat));
  NOR3_X1   g614(.A1(new_n570), .A2(G106gat), .A3(new_n691), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n794), .A2(new_n796), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n736), .A2(new_n737), .A3(new_n425), .A4(new_n782), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(G106gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n823));
  NOR4_X1   g622(.A1(new_n506), .A2(new_n823), .A3(new_n671), .A4(new_n781), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n816), .B1(new_n824), .B2(new_n791), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n820), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n822), .B1(new_n826), .B2(KEYINPUT53), .ZN(new_n827));
  AOI211_X1 g626(.A(KEYINPUT112), .B(new_n818), .C1(new_n820), .C2(new_n825), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n821), .B1(new_n827), .B2(new_n828), .ZN(G1339gat));
  NOR2_X1   g628(.A1(new_n692), .A2(new_n569), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n562), .A2(new_n555), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n541), .B1(new_n540), .B2(new_n545), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n552), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n668), .A2(new_n670), .A3(new_n560), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n675), .A2(new_n676), .A3(new_n687), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n679), .A2(KEYINPUT54), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n682), .B1(new_n688), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n836), .A2(KEYINPUT55), .A3(new_n838), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n684), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT113), .B1(new_n834), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n684), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT55), .B1(new_n836), .B2(new_n838), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n560), .A2(new_n833), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n847), .A2(new_n848), .A3(new_n728), .A4(new_n849), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n690), .A2(new_n560), .A3(new_n833), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n851), .B1(new_n847), .B2(new_n569), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n844), .B(new_n850), .C1(new_n852), .C2(new_n728), .ZN(new_n853));
  INV_X1    g652(.A(new_n626), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n830), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n384), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n586), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(G113gat), .B1(new_n858), .B2(new_n569), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n855), .A2(new_n425), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n384), .A2(new_n434), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n712), .A3(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(G113gat), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n862), .A2(new_n863), .A3(new_n565), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n859), .A2(new_n864), .ZN(G1340gat));
  OAI21_X1  g664(.A(G120gat), .B1(new_n862), .B2(new_n691), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n690), .A2(new_n232), .ZN(new_n867));
  XOR2_X1   g666(.A(new_n867), .B(KEYINPUT114), .Z(new_n868));
  OAI21_X1  g667(.A(new_n866), .B1(new_n857), .B2(new_n868), .ZN(G1341gat));
  NAND3_X1  g668(.A1(new_n858), .A2(new_n626), .A3(new_n206), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n862), .A2(new_n854), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n206), .B2(new_n871), .ZN(G1342gat));
  NOR3_X1   g671(.A1(new_n857), .A2(G134gat), .A3(new_n671), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n862), .B2(new_n671), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n878), .A2(KEYINPUT115), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(KEYINPUT115), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n875), .B(new_n876), .C1(new_n879), .C2(new_n880), .ZN(G1343gat));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n493), .A2(new_n570), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n453), .ZN(new_n884));
  INV_X1    g683(.A(new_n856), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(G141gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n569), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT118), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n855), .A2(new_n891), .A3(new_n570), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n855), .B2(new_n570), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT116), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n895), .B(new_n891), .C1(new_n855), .C2(new_n570), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n892), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n578), .A2(new_n861), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n897), .A2(new_n565), .A3(new_n898), .ZN(new_n899));
  OAI221_X1 g698(.A(new_n882), .B1(new_n887), .B2(new_n890), .C1(new_n899), .C2(new_n888), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n887), .A2(new_n890), .ZN(new_n901));
  INV_X1    g700(.A(new_n892), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n849), .A2(new_n690), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n903), .B1(new_n843), .B2(new_n565), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n842), .A2(new_n684), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n728), .A2(new_n905), .A3(new_n841), .A4(new_n849), .ZN(new_n906));
  AOI22_X1  g705(.A1(new_n671), .A2(new_n904), .B1(new_n906), .B2(KEYINPUT113), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n626), .B1(new_n907), .B2(new_n850), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n425), .B1(new_n908), .B2(new_n830), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n895), .B1(new_n909), .B2(new_n891), .ZN(new_n910));
  INV_X1    g709(.A(new_n896), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n902), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n898), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(KEYINPUT117), .A3(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(new_n897), .B2(new_n898), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n914), .A2(new_n916), .A3(new_n569), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n901), .B1(new_n917), .B2(G141gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n900), .B1(new_n918), .B2(new_n882), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT119), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g720(.A(KEYINPUT119), .B(new_n900), .C1(new_n918), .C2(new_n882), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1344gat));
  NAND3_X1  g722(.A1(new_n914), .A2(new_n916), .A3(new_n690), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(new_n925), .A3(G148gat), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n913), .A2(new_n690), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n906), .B1(new_n852), .B2(new_n728), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n928), .A2(new_n854), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n425), .B1(new_n929), .B2(new_n830), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n892), .B1(new_n891), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G148gat), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT59), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n926), .A2(KEYINPUT120), .A3(new_n933), .ZN(new_n934));
  OR3_X1    g733(.A1(new_n887), .A2(G148gat), .A3(new_n691), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n934), .B(new_n935), .C1(KEYINPUT120), .C2(new_n926), .ZN(G1345gat));
  NAND3_X1  g735(.A1(new_n886), .A2(new_n239), .A3(new_n626), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n914), .A2(new_n626), .A3(new_n916), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n239), .ZN(G1346gat));
  NAND4_X1  g738(.A1(new_n914), .A2(new_n916), .A3(G162gat), .A4(new_n728), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n240), .B1(new_n887), .B2(new_n671), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n940), .A2(new_n941), .ZN(G1347gat));
  NOR2_X1   g741(.A1(new_n290), .A2(new_n453), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n773), .A2(new_n860), .A3(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(G169gat), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n944), .A2(new_n945), .A3(new_n565), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n384), .B1(new_n908), .B2(new_n830), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT121), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n434), .A3(new_n501), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n569), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n946), .B1(new_n951), .B2(new_n945), .ZN(G1348gat));
  OAI21_X1  g751(.A(G176gat), .B1(new_n944), .B2(new_n691), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n691), .A2(G176gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n949), .B2(new_n954), .ZN(G1349gat));
  OAI21_X1  g754(.A(G183gat), .B1(new_n944), .B2(new_n854), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n626), .A2(new_n324), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n949), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g758(.A(G190gat), .B1(new_n944), .B2(new_n671), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT61), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n728), .A2(new_n307), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n949), .B2(new_n962), .ZN(G1351gat));
  NAND3_X1  g762(.A1(new_n948), .A2(new_n434), .A3(new_n883), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(G197gat), .B1(new_n965), .B2(new_n569), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n931), .B(KEYINPUT122), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n578), .A2(new_n943), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(G197gat), .A3(new_n569), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n966), .B1(new_n967), .B2(new_n970), .ZN(G1352gat));
  NOR3_X1   g770(.A1(new_n964), .A2(G204gat), .A3(new_n691), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT62), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n967), .A2(new_n690), .A3(new_n969), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT123), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(G204gat), .B1(new_n974), .B2(new_n975), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(G1353gat));
  NAND2_X1  g777(.A1(new_n969), .A2(new_n626), .ZN(new_n979));
  OAI21_X1  g778(.A(G211gat), .B1(new_n979), .B2(new_n931), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT63), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  OAI221_X1 g782(.A(G211gat), .B1(KEYINPUT124), .B2(KEYINPUT63), .C1(new_n979), .C2(new_n931), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n983), .B(new_n984), .C1(new_n981), .C2(new_n982), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n626), .A2(new_n342), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n985), .B1(new_n964), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(KEYINPUT125), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n985), .B(new_n989), .C1(new_n964), .C2(new_n986), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n988), .A2(new_n990), .ZN(G1354gat));
  AOI21_X1  g790(.A(G218gat), .B1(new_n965), .B2(new_n728), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n671), .A2(new_n343), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n993), .B(KEYINPUT126), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n968), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n992), .B1(new_n967), .B2(new_n995), .ZN(G1355gat));
endmodule


