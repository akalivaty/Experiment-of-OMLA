//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n521,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  AND2_X1   g048(.A1(new_n461), .A2(new_n463), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(new_n471), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n477), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND3_X1  g059(.A1(new_n461), .A2(new_n463), .A3(G126), .ZN(new_n485));
  NAND2_X1  g060(.A1(G114), .A2(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n471), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  OAI22_X1  g064(.A1(new_n487), .A2(new_n488), .B1(new_n478), .B2(new_n489), .ZN(new_n490));
  NOR3_X1   g065(.A1(new_n464), .A2(new_n488), .A3(new_n489), .ZN(new_n491));
  AND2_X1   g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n471), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n496));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(KEYINPUT6), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(KEYINPUT67), .A3(G651), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n498), .A2(new_n500), .B1(KEYINPUT6), .B2(new_n497), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(G62), .A3(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n498), .A2(new_n500), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n497), .A2(KEYINPUT6), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(new_n505), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n504), .A2(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  NAND3_X1  g088(.A1(new_n501), .A2(G51), .A3(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n501), .A2(G89), .A3(new_n505), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n514), .A2(new_n515), .A3(new_n516), .A4(new_n518), .ZN(G286));
  INV_X1    g094(.A(G286), .ZN(G168));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G543), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n522), .A2(new_n524), .A3(G64), .ZN(new_n525));
  NAND2_X1  g100(.A1(G77), .A2(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n497), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n507), .A2(G543), .A3(new_n508), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(G52), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n501), .A2(G90), .A3(new_n505), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n521), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n527), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n501), .A2(G52), .A3(G543), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n532), .A2(new_n530), .A3(new_n533), .A4(new_n521), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n531), .A2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  NAND2_X1  g112(.A1(new_n522), .A2(new_n524), .ZN(new_n538));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  INV_X1    g114(.A(G68), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n538), .A2(new_n539), .B1(new_n540), .B2(new_n503), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT69), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI221_X1 g118(.A(KEYINPUT69), .B1(new_n540), .B2(new_n503), .C1(new_n538), .C2(new_n539), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n543), .A2(G651), .A3(new_n544), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n507), .A2(G43), .A3(G543), .A4(new_n508), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n507), .A2(G81), .A3(new_n508), .A4(new_n505), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT70), .ZN(new_n548));
  AOI21_X1  g123(.A(KEYINPUT70), .B1(new_n546), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT71), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT72), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n559), .B(KEYINPUT73), .Z(G188));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n509), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n501), .A2(KEYINPUT75), .A3(new_n505), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G91), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n501), .A2(G53), .A3(G543), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n569));
  OR3_X1    g144(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n538), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n566), .A2(new_n568), .B1(G651), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n565), .A2(new_n570), .A3(new_n574), .ZN(G299));
  NAND2_X1  g150(.A1(new_n564), .A2(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n528), .A2(G49), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n564), .A2(G87), .B1(G49), .B2(new_n528), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n582), .A2(KEYINPUT76), .A3(new_n577), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(G288));
  NAND3_X1  g159(.A1(new_n501), .A2(G48), .A3(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n538), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n501), .A2(new_n591), .A3(G48), .A4(G543), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n586), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n562), .B2(new_n563), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n593), .A2(new_n595), .ZN(G305));
  INV_X1    g171(.A(new_n509), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G85), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  INV_X1    g174(.A(new_n528), .ZN(new_n600));
  XOR2_X1   g175(.A(KEYINPUT78), .B(G47), .Z(new_n601));
  OAI221_X1 g176(.A(new_n598), .B1(new_n497), .B2(new_n599), .C1(new_n600), .C2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n538), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n528), .A2(G54), .B1(new_n606), .B2(G651), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT10), .B1(new_n564), .B2(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  AOI211_X1 g185(.A(new_n609), .B(new_n610), .C1(new_n562), .C2(new_n563), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n607), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT79), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(KEYINPUT80), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(KEYINPUT80), .ZN(new_n615));
  AND2_X1   g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n603), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n603), .B1(new_n616), .B2(G868), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  AND3_X1   g194(.A1(new_n565), .A2(new_n570), .A3(new_n574), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n614), .A2(new_n615), .ZN(new_n625));
  OR3_X1    g200(.A1(new_n625), .A2(KEYINPUT81), .A3(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(KEYINPUT81), .B1(new_n625), .B2(G559), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g206(.A1(new_n460), .A2(G2105), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n474), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT82), .B(G2100), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n638), .B(G2104), .C1(G111), .C2(new_n471), .ZN(new_n639));
  INV_X1    g214(.A(G123), .ZN(new_n640));
  INV_X1    g215(.A(G135), .ZN(new_n641));
  OAI221_X1 g216(.A(new_n639), .B1(new_n475), .B2(new_n640), .C1(new_n641), .C2(new_n478), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n637), .A2(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2435), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2438), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT14), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2451), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n655), .B(new_n656), .Z(new_n657));
  AND2_X1   g232(.A1(new_n657), .A2(G14), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2067), .B(G2678), .Z(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(new_n663), .A3(KEYINPUT17), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n662), .B2(KEYINPUT18), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT84), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n673), .A2(new_n674), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n678), .A3(new_n680), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n683), .B(new_n684), .C1(new_n682), .C2(new_n681), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(G1986), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT22), .B(G1981), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n689), .B(new_n690), .Z(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G35), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G162), .B2(new_n693), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT29), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n696), .A2(G2090), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT28), .ZN(new_n698));
  INV_X1    g273(.A(G26), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(G29), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(G29), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n476), .A2(G128), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n479), .A2(G140), .ZN(new_n703));
  NOR2_X1   g278(.A1(G104), .A2(G2105), .ZN(new_n704));
  OAI21_X1  g279(.A(G2104), .B1(new_n471), .B2(G116), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n702), .B(new_n703), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n701), .B1(new_n706), .B2(G29), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n700), .B1(new_n707), .B2(new_n698), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n696), .A2(G2090), .B1(G2067), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G21), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G168), .B2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G1966), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(KEYINPUT24), .A2(G34), .ZN(new_n715));
  NAND2_X1  g290(.A1(KEYINPUT24), .A2(G34), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n715), .A2(new_n693), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G160), .B2(new_n693), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT89), .Z(new_n719));
  INV_X1    g294(.A(G2084), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n697), .A2(new_n709), .A3(new_n714), .A4(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(G5), .A2(G16), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G171), .B2(G16), .ZN(new_n724));
  INV_X1    g299(.A(G1961), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G1341), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n551), .A2(G16), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G16), .B2(G19), .ZN(new_n729));
  OAI221_X1 g304(.A(new_n726), .B1(new_n727), .B2(new_n729), .C1(new_n720), .C2(new_n719), .ZN(new_n730));
  INV_X1    g305(.A(G2072), .ZN(new_n731));
  OR2_X1    g306(.A1(G29), .A2(G33), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT25), .Z(new_n734));
  INV_X1    g309(.A(G139), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n736));
  OAI221_X1 g311(.A(new_n734), .B1(new_n478), .B2(new_n735), .C1(new_n736), .C2(new_n471), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT88), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n732), .B1(new_n738), .B2(new_n693), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n722), .B(new_n730), .C1(new_n731), .C2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G4), .B2(G16), .ZN(new_n742));
  OR3_X1    g317(.A1(new_n741), .A2(G4), .A3(G16), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n742), .B(new_n743), .C1(new_n625), .C2(new_n710), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1348), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n693), .A2(G27), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G164), .B2(new_n693), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2078), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(G28), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(G28), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n750), .A2(new_n751), .A3(new_n693), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n752), .B1(new_n693), .B2(new_n642), .C1(new_n739), .C2(new_n731), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n748), .B(new_n753), .C1(new_n727), .C2(new_n729), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n710), .A2(KEYINPUT23), .A3(G20), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT23), .ZN(new_n756));
  INV_X1    g331(.A(G20), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(G16), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n755), .B(new_n758), .C1(new_n620), .C2(new_n710), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT91), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1956), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n740), .A2(new_n745), .A3(new_n754), .A4(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  MUX2_X1   g338(.A(G23), .B(new_n579), .S(G16), .Z(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT33), .B(G1976), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n710), .A2(G6), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n593), .A2(new_n595), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(new_n710), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT32), .B(G1981), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT86), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n769), .B(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G16), .A2(G22), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G166), .B2(G16), .ZN(new_n774));
  INV_X1    g349(.A(G1971), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n766), .A2(new_n772), .A3(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT34), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n476), .A2(G119), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n479), .A2(G131), .ZN(new_n780));
  NOR2_X1   g355(.A1(G95), .A2(G2105), .ZN(new_n781));
  OAI21_X1  g356(.A(G2104), .B1(new_n471), .B2(G107), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n779), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  MUX2_X1   g358(.A(G25), .B(new_n783), .S(G29), .Z(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT35), .B(G1991), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT85), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n784), .B(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(G1986), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n710), .A2(G24), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G290), .B2(G16), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n787), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n788), .B2(new_n790), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n778), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT36), .ZN(new_n794));
  NOR2_X1   g369(.A1(G29), .A2(G32), .ZN(new_n795));
  AOI22_X1  g370(.A1(G129), .A2(new_n476), .B1(new_n479), .B2(G141), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n632), .A2(G105), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT90), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT26), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n795), .B1(new_n803), .B2(G29), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT27), .B(G1996), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT31), .B(G11), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n763), .A2(new_n794), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n708), .A2(G2067), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n808), .A2(new_n810), .ZN(G311));
  INV_X1    g386(.A(G311), .ZN(G150));
  NAND2_X1  g387(.A1(new_n616), .A2(G559), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT38), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n550), .A2(KEYINPUT92), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n597), .A2(G93), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(new_n497), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n528), .A2(G55), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT92), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n545), .B(new_n822), .C1(new_n548), .C2(new_n549), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n815), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n821), .B1(new_n815), .B2(new_n823), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n814), .B(new_n827), .ZN(new_n828));
  OR3_X1    g403(.A1(new_n828), .A2(KEYINPUT93), .A3(KEYINPUT39), .ZN(new_n829));
  AOI21_X1  g404(.A(G860), .B1(new_n828), .B2(KEYINPUT39), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT93), .B1(new_n828), .B2(KEYINPUT39), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n820), .A2(G860), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT37), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(G145));
  XNOR2_X1  g410(.A(new_n802), .B(new_n783), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n471), .A2(G118), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT94), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n838), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n479), .A2(G142), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n476), .A2(G130), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n836), .B(new_n842), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n738), .B(new_n494), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n642), .B(G160), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n483), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n844), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n843), .B(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n706), .B(new_n634), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(G37), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n620), .ZN(new_n854));
  OAI211_X1 g429(.A(G299), .B(new_n607), .C1(new_n608), .C2(new_n611), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT41), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n855), .A3(KEYINPUT95), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n608), .A2(new_n611), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT95), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n858), .A2(new_n859), .A3(G299), .A4(new_n607), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n856), .B1(new_n861), .B2(KEYINPUT41), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n626), .A2(new_n627), .A3(new_n826), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n826), .B1(new_n626), .B2(new_n627), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n865), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(new_n861), .A3(new_n863), .ZN(new_n868));
  XNOR2_X1  g443(.A(G305), .B(G303), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n579), .B(G290), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n871), .A2(KEYINPUT96), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT42), .Z(new_n873));
  NAND3_X1  g448(.A1(new_n866), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n873), .B1(new_n866), .B2(new_n868), .ZN(new_n876));
  OAI21_X1  g451(.A(G868), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n821), .A2(G868), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(G295));
  INV_X1    g455(.A(G868), .ZN(new_n881));
  INV_X1    g456(.A(new_n873), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n867), .A2(new_n861), .A3(new_n863), .ZN(new_n883));
  INV_X1    g458(.A(new_n862), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n867), .B2(new_n863), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n882), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n881), .B1(new_n886), .B2(new_n874), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT97), .B1(new_n887), .B2(new_n878), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT97), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n877), .A2(new_n889), .A3(new_n879), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(G331));
  OAI21_X1  g466(.A(G168), .B1(new_n531), .B2(new_n535), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n532), .A2(new_n530), .A3(new_n533), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT68), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(G286), .A3(new_n534), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n824), .A2(new_n825), .A3(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n894), .A2(G286), .A3(new_n534), .ZN(new_n898));
  AOI21_X1  g473(.A(G286), .B1(new_n894), .B2(new_n534), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n546), .A2(new_n547), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT70), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT70), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n822), .B1(new_n905), .B2(new_n545), .ZN(new_n906));
  INV_X1    g481(.A(new_n823), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n820), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n815), .A2(new_n821), .A3(new_n823), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n900), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n860), .B(new_n857), .C1(new_n897), .C2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n896), .B1(new_n824), .B2(new_n825), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(new_n900), .A3(new_n909), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n911), .B(new_n871), .C1(new_n862), .C2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(KEYINPUT41), .A3(new_n913), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n861), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n869), .A2(new_n870), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n869), .A2(new_n870), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n854), .A2(new_n855), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n912), .A2(new_n921), .A3(new_n913), .A4(KEYINPUT41), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n915), .A2(new_n923), .A3(new_n851), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT98), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT98), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n915), .A2(new_n923), .A3(new_n926), .A4(new_n851), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(KEYINPUT43), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT99), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n862), .A2(new_n914), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n871), .B1(new_n931), .B2(new_n911), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n915), .A2(new_n851), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n932), .A2(new_n933), .A3(KEYINPUT43), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n925), .A2(KEYINPUT99), .A3(KEYINPUT43), .A4(new_n927), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n930), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT100), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n930), .A2(new_n936), .A3(KEYINPUT100), .A4(new_n937), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT43), .B1(new_n932), .B2(new_n933), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(KEYINPUT43), .B2(new_n924), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n935), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT101), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n942), .A2(new_n948), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(G397));
  INV_X1    g525(.A(G8), .ZN(new_n951));
  NOR2_X1   g526(.A1(G168), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n467), .A2(new_n472), .A3(G40), .ZN(new_n953));
  AOI21_X1  g528(.A(G1384), .B1(new_n490), .B2(new_n493), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n953), .B1(new_n954), .B2(KEYINPUT45), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT112), .B1(new_n954), .B2(KEYINPUT45), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(KEYINPUT112), .A3(KEYINPUT45), .ZN(new_n958));
  AOI21_X1  g533(.A(G1966), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G1384), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n494), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(KEYINPUT50), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n953), .B1(new_n954), .B2(new_n963), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n962), .A2(new_n964), .A3(G2084), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n959), .A2(KEYINPUT118), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT118), .ZN(new_n967));
  INV_X1    g542(.A(new_n953), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n968), .B1(new_n961), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n954), .A2(KEYINPUT45), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n970), .A2(new_n973), .A3(new_n958), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n713), .ZN(new_n975));
  INV_X1    g550(.A(new_n965), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n967), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n952), .B1(new_n966), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT118), .B1(new_n959), .B2(new_n965), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n975), .A2(new_n976), .A3(new_n967), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n951), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT119), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n952), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(G8), .B1(new_n966), .B2(new_n977), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT119), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n979), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  AOI211_X1 g562(.A(new_n951), .B(G286), .C1(new_n975), .C2(new_n976), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n988), .A2(KEYINPUT51), .A3(new_n952), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n978), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n501), .A2(G86), .A3(new_n505), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n586), .A2(new_n590), .A3(new_n592), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(G1981), .ZN(new_n993));
  OAI211_X1 g568(.A(KEYINPUT49), .B(new_n993), .C1(G305), .C2(G1981), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n995));
  INV_X1    g570(.A(new_n993), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n593), .A2(new_n595), .A3(G1981), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n951), .B1(new_n954), .B2(new_n953), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n994), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n576), .A2(G1976), .A3(new_n577), .A4(new_n578), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT104), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT104), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n582), .A2(new_n1003), .A3(G1976), .A4(new_n577), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n999), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT52), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1000), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1976), .B1(new_n581), .B2(new_n583), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1008), .A2(new_n1005), .A3(KEYINPUT52), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT111), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1976), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G288), .A2(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n999), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(new_n1006), .A4(new_n1000), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1010), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT102), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n971), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n954), .A2(KEYINPUT102), .A3(KEYINPUT45), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n970), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n775), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n962), .A2(new_n964), .ZN(new_n1024));
  INV_X1    g599(.A(G2090), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G303), .A2(G8), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT103), .B(KEYINPUT55), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  OR3_X1    g605(.A1(new_n1027), .A2(new_n951), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1018), .A2(new_n1031), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n954), .A2(KEYINPUT108), .A3(new_n963), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT108), .B1(new_n954), .B2(new_n963), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT107), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n964), .A2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT107), .B(new_n953), .C1(new_n954), .C2(new_n963), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1035), .A2(new_n1025), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(new_n1023), .A3(KEYINPUT109), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G8), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT109), .B1(new_n1039), .B2(new_n1023), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1030), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT110), .B(new_n1030), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1032), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n1048));
  INV_X1    g623(.A(G2078), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n970), .A2(new_n1020), .A3(new_n1049), .A4(new_n1021), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n962), .A2(new_n964), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n725), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT102), .B1(new_n954), .B2(KEYINPUT45), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n955), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1056), .A2(KEYINPUT53), .A3(new_n1049), .A4(new_n1021), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(G171), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1050), .A2(new_n1051), .B1(new_n1053), .B2(new_n725), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n957), .A2(KEYINPUT53), .A3(new_n1049), .A4(new_n958), .ZN(new_n1061));
  AOI21_X1  g636(.A(G301), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1048), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(KEYINPUT120), .B(new_n1048), .C1(new_n1059), .C2(new_n1062), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1058), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1060), .A2(KEYINPUT121), .A3(new_n1057), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(G171), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1060), .A2(G301), .A3(new_n1061), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1072), .A3(KEYINPUT54), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT122), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1071), .A2(new_n1072), .A3(new_n1075), .A4(KEYINPUT54), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n990), .A2(new_n1047), .A3(new_n1067), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT123), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n620), .B(KEYINPUT57), .ZN(new_n1080));
  XOR2_X1   g655(.A(new_n1080), .B(KEYINPUT115), .Z(new_n1081));
  INV_X1    g656(.A(G1956), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1022), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT56), .B(G2072), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1082), .A2(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1081), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1348), .ZN(new_n1088));
  INV_X1    g663(.A(G2067), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n961), .A2(new_n968), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1053), .A2(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1086), .B2(new_n1080), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1087), .B1(new_n1092), .B2(new_n613), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1091), .A2(KEYINPUT60), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n613), .B1(new_n1091), .B2(KEYINPUT60), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1097));
  AND2_X1   g672(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1090), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1996), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n970), .A2(new_n1020), .A3(new_n1100), .A4(new_n1021), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1056), .A2(KEYINPUT116), .A3(new_n1100), .A4(new_n1021), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1099), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI211_X1 g682(.A(KEYINPUT117), .B(new_n1099), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n551), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT59), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1111), .B(new_n551), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1096), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1086), .A2(new_n1080), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1114), .B(KEYINPUT61), .Z(new_n1115));
  INV_X1    g690(.A(new_n613), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1094), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1086), .A2(new_n1080), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1093), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1047), .A2(new_n1067), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1121), .A2(new_n1122), .A3(new_n990), .A4(new_n1077), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1079), .A2(new_n1120), .A3(new_n1123), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(new_n1047), .A4(new_n1062), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1027), .A2(new_n951), .A3(new_n1030), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n997), .B(KEYINPUT106), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1000), .A2(new_n1011), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1132), .B2(G288), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n999), .B(KEYINPUT105), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT63), .B1(new_n1047), .B2(new_n988), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1031), .A2(KEYINPUT63), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1030), .B1(new_n1027), .B2(new_n951), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(new_n988), .A3(new_n1129), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT113), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1140), .A2(new_n988), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT63), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1128), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT113), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1143), .A2(new_n1145), .A3(new_n1146), .A4(new_n1129), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1137), .B1(new_n1138), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT114), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g726(.A(KEYINPUT114), .B(new_n1137), .C1(new_n1138), .C2(new_n1148), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1124), .A2(new_n1127), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n803), .A2(new_n1100), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n706), .B(new_n1089), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n783), .A2(new_n785), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n802), .A2(G1996), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1158), .B1(new_n783), .B2(new_n785), .ZN(new_n1159));
  OR2_X1    g734(.A1(G290), .A2(G1986), .ZN(new_n1160));
  NAND2_X1  g735(.A1(G290), .A2(G1986), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n961), .A2(new_n969), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1163), .A2(new_n968), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1153), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1164), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n1155), .B2(new_n803), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT124), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT46), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI22_X1  g746(.A1(new_n1167), .A2(G1996), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1164), .A2(KEYINPUT124), .A3(KEYINPUT46), .A4(new_n1100), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT47), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n1176), .A2(new_n1156), .B1(G2067), .B2(new_n706), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n1164), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1167), .A2(new_n1160), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT48), .Z(new_n1180));
  OAI21_X1  g755(.A(new_n1180), .B1(new_n1159), .B2(new_n1167), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1175), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT125), .Z(new_n1183));
  NAND2_X1  g758(.A1(new_n1166), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g759(.A1(new_n944), .A2(G319), .ZN(new_n1186));
  NOR2_X1   g760(.A1(G401), .A2(G227), .ZN(new_n1187));
  NAND4_X1  g761(.A1(new_n1186), .A2(new_n691), .A3(new_n852), .A4(new_n1187), .ZN(G225));
  XOR2_X1   g762(.A(G225), .B(KEYINPUT126), .Z(G308));
endmodule


