//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  AND2_X1   g000(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n187));
  NOR2_X1   g001(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G143), .B(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G128), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(G143), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n191), .A2(new_n195), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G104), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(G107), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n204), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n206), .A2(G104), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n203), .A2(G107), .ZN(new_n212));
  OAI21_X1  g026(.A(G101), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n202), .A2(new_n214), .A3(KEYINPUT10), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT79), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT79), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n202), .A2(new_n214), .A3(new_n217), .A4(KEYINPUT10), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n190), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AND4_X1   g035(.A1(KEYINPUT0), .A2(new_n196), .A3(new_n198), .A4(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n204), .A2(new_n207), .A3(new_n209), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(G101), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n224), .A2(G101), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n210), .A2(KEYINPUT4), .ZN(new_n229));
  OR2_X1    g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n216), .A2(new_n218), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT76), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n196), .A2(new_n198), .A3(G128), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(new_n192), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n193), .A2(G143), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n199), .A2(new_n200), .B1(KEYINPUT1), .B2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n189), .A2(new_n190), .A3(KEYINPUT76), .A4(G128), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT77), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n240), .A2(new_n241), .A3(new_n214), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(new_n240), .B2(new_n214), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n233), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT11), .ZN(new_n245));
  INV_X1    g059(.A(G134), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n245), .B1(new_n246), .B2(G137), .ZN(new_n247));
  INV_X1    g061(.A(G137), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT11), .A3(G134), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(G137), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n247), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G131), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(KEYINPUT64), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n251), .B(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n231), .A2(new_n244), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G227), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n258), .B(KEYINPUT75), .ZN(new_n259));
  XNOR2_X1  g073(.A(G110), .B(G140), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n259), .B(new_n260), .ZN(new_n261));
  OAI22_X1  g075(.A1(new_n242), .A2(new_n243), .B1(new_n202), .B2(new_n214), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n262), .A2(KEYINPUT12), .A3(new_n254), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT12), .B1(new_n262), .B2(new_n254), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n256), .B(new_n261), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n261), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n231), .A2(new_n255), .A3(new_n244), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n255), .B1(new_n231), .B2(new_n244), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G469), .ZN(new_n271));
  INV_X1    g085(.A(G902), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(G469), .A2(G902), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n256), .B1(new_n263), .B2(new_n264), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n266), .ZN(new_n276));
  OR3_X1    g090(.A1(new_n267), .A2(new_n268), .A3(new_n266), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(G469), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n273), .A2(new_n274), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT9), .B(G234), .ZN(new_n280));
  OAI21_X1  g094(.A(G221), .B1(new_n280), .B2(G902), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(KEYINPUT80), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT80), .B1(new_n279), .B2(new_n281), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G217), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(G234), .B2(new_n272), .ZN(new_n287));
  INV_X1    g101(.A(G140), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G125), .ZN(new_n289));
  INV_X1    g103(.A(G125), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G140), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n291), .A3(KEYINPUT16), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT16), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n288), .A3(G125), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n193), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n292), .A2(G146), .A3(new_n294), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n295), .A2(KEYINPUT73), .A3(new_n193), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n301));
  INV_X1    g115(.A(G119), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(G128), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n303), .B(new_n304), .C1(G119), .C2(new_n200), .ZN(new_n305));
  XNOR2_X1  g119(.A(G119), .B(G128), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT24), .B(G110), .Z(new_n307));
  AOI22_X1  g121(.A1(new_n305), .A2(G110), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n299), .A2(new_n300), .A3(new_n308), .ZN(new_n309));
  OAI22_X1  g123(.A1(new_n305), .A2(G110), .B1(new_n306), .B2(new_n307), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n289), .A2(new_n291), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n193), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n298), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT74), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT22), .B(G137), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n314), .B(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT25), .A3(new_n272), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT25), .B1(new_n320), .B2(new_n272), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n287), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n287), .A2(G902), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G237), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n257), .A3(G210), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT27), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT26), .B(G101), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n254), .A2(new_n223), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n252), .B1(G134), .B2(new_n248), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n251), .A2(new_n252), .B1(new_n250), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT65), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n202), .B1(new_n338), .B2(KEYINPUT65), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n336), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n302), .A2(G116), .ZN(new_n343));
  INV_X1    g157(.A(G116), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G119), .ZN(new_n345));
  INV_X1    g159(.A(G113), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n346), .A2(KEYINPUT2), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(KEYINPUT2), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n343), .B(new_n345), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n343), .A2(new_n345), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT2), .B(G113), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n342), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n251), .A2(new_n252), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n337), .A2(new_n250), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT67), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n338), .A2(KEYINPUT67), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(new_n202), .ZN(new_n361));
  INV_X1    g175(.A(new_n353), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n336), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n335), .B1(new_n354), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT28), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n333), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n360), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n202), .B1(new_n338), .B2(KEYINPUT67), .ZN(new_n370));
  OAI211_X1 g184(.A(KEYINPUT30), .B(new_n336), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT65), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n200), .A2(new_n199), .B1(new_n192), .B2(new_n194), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n357), .A2(new_n372), .B1(new_n191), .B2(new_n373), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n374), .A2(new_n339), .B1(new_n254), .B2(new_n223), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n353), .B(new_n371), .C1(new_n375), .C2(KEYINPUT30), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT31), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n376), .A2(new_n377), .A3(new_n363), .A4(new_n332), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n368), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n363), .A3(new_n332), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT68), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n376), .A2(KEYINPUT68), .A3(new_n363), .A4(new_n332), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(KEYINPUT31), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT72), .ZN(new_n386));
  NOR2_X1   g200(.A1(G472), .A2(G902), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT32), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n385), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n386), .B1(new_n385), .B2(new_n390), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n385), .A2(new_n387), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n376), .A2(new_n363), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n333), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n364), .A2(new_n367), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n395), .B(new_n397), .C1(new_n398), .C2(new_n333), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT71), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n366), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n363), .A2(KEYINPUT71), .A3(new_n365), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT70), .ZN(new_n404));
  INV_X1    g218(.A(new_n363), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n362), .B1(new_n361), .B2(new_n336), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n404), .B1(new_n407), .B2(new_n365), .ZN(new_n408));
  OAI211_X1 g222(.A(KEYINPUT70), .B(KEYINPUT28), .C1(new_n405), .C2(new_n406), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n333), .A2(new_n395), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n403), .A2(new_n408), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n399), .A2(new_n272), .A3(new_n411), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n394), .A2(new_n389), .B1(new_n412), .B2(G472), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n327), .B1(new_n393), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT20), .ZN(new_n415));
  XNOR2_X1  g229(.A(G113), .B(G122), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(new_n203), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n328), .A2(new_n257), .A3(G214), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(G143), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n420));
  OR3_X1    g234(.A1(new_n419), .A2(new_n420), .A3(new_n252), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n311), .B(new_n193), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n419), .B1(new_n420), .B2(new_n252), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n299), .A2(KEYINPUT85), .A3(new_n300), .ZN(new_n425));
  INV_X1    g239(.A(new_n419), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(KEYINPUT17), .A3(G131), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n298), .A2(new_n297), .ZN(new_n430));
  AOI21_X1  g244(.A(G146), .B1(new_n292), .B2(new_n294), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n300), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n429), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT86), .B1(new_n428), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n434), .A2(KEYINPUT86), .A3(new_n425), .A4(new_n427), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n419), .B(new_n252), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n437), .A2(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n417), .B(new_n424), .C1(new_n435), .C2(new_n439), .ZN(new_n440));
  XOR2_X1   g254(.A(new_n311), .B(KEYINPUT19), .Z(new_n441));
  OAI211_X1 g255(.A(new_n437), .B(new_n298), .C1(G146), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n424), .ZN(new_n443));
  INV_X1    g257(.A(new_n417), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(G475), .A2(G902), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n415), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n447), .ZN(new_n449));
  AOI211_X1 g263(.A(KEYINPUT20), .B(new_n449), .C1(new_n440), .C2(new_n445), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n424), .B1(new_n435), .B2(new_n439), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n444), .ZN(new_n452));
  AOI21_X1  g266(.A(G902), .B1(new_n452), .B2(new_n440), .ZN(new_n453));
  INV_X1    g267(.A(G475), .ZN(new_n454));
  OAI22_X1  g268(.A1(new_n448), .A2(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G210), .B1(G237), .B2(G902), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT7), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n257), .A2(G224), .ZN(new_n459));
  OAI21_X1  g273(.A(G125), .B1(new_n221), .B2(new_n222), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT82), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n191), .A2(new_n290), .A3(new_n201), .A4(new_n195), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n373), .A2(KEYINPUT82), .A3(new_n290), .A4(new_n191), .ZN(new_n464));
  AOI211_X1 g278(.A(new_n458), .B(new_n459), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT83), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n459), .B1(new_n466), .B2(new_n458), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n466), .B2(new_n458), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n463), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  XOR2_X1   g283(.A(G110), .B(G122), .Z(new_n470));
  XOR2_X1   g284(.A(new_n470), .B(KEYINPUT8), .Z(new_n471));
  INV_X1    g285(.A(KEYINPUT5), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n302), .A3(G116), .ZN(new_n473));
  OAI211_X1 g287(.A(G113), .B(new_n473), .C1(new_n350), .C2(new_n472), .ZN(new_n474));
  AND4_X1   g288(.A1(new_n349), .A2(new_n474), .A3(new_n213), .A4(new_n210), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n474), .A2(new_n349), .B1(new_n213), .B2(new_n210), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n471), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT84), .B1(new_n465), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n353), .B(new_n226), .C1(new_n228), .C2(new_n229), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n214), .A2(new_n349), .A3(new_n474), .ZN(new_n481));
  INV_X1    g295(.A(new_n470), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n463), .A2(new_n464), .ZN(new_n484));
  INV_X1    g298(.A(new_n459), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(KEYINPUT7), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT84), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n469), .A4(new_n477), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n479), .A2(new_n483), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n484), .A2(new_n485), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n463), .A2(new_n459), .A3(new_n464), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n480), .A2(new_n481), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n470), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(KEYINPUT6), .A3(new_n483), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n496));
  AND4_X1   g310(.A1(KEYINPUT81), .A2(new_n493), .A3(new_n496), .A4(new_n470), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n482), .B1(new_n480), .B2(new_n481), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT81), .B1(new_n498), .B2(new_n496), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n492), .B(new_n495), .C1(new_n497), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n272), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n457), .B1(new_n489), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n479), .A2(new_n483), .A3(new_n488), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n503), .A2(new_n272), .A3(new_n456), .A4(new_n500), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  XOR2_X1   g320(.A(G116), .B(G122), .Z(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G107), .ZN(new_n508));
  XNOR2_X1  g322(.A(G116), .B(G122), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n206), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n200), .A2(G143), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT13), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n246), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G128), .B(G143), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n508), .A2(new_n510), .A3(KEYINPUT87), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n513), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n280), .A2(new_n286), .A3(G953), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(KEYINPUT88), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n344), .A2(KEYINPUT14), .A3(G122), .ZN(new_n523));
  OAI211_X1 g337(.A(G107), .B(new_n523), .C1(new_n507), .C2(KEYINPUT14), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n517), .A2(G134), .ZN(new_n525));
  OR2_X1    g339(.A1(new_n517), .A2(G134), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n524), .A2(new_n510), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n520), .A2(new_n522), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n522), .B1(new_n520), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n272), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT89), .ZN(new_n531));
  INV_X1    g345(.A(G478), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT90), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT89), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n537), .B(new_n272), .C1(new_n528), .C2(new_n529), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n531), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n530), .A2(new_n536), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n257), .A2(G952), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(G234), .B2(G237), .ZN(new_n543));
  AOI211_X1 g357(.A(new_n272), .B(new_n257), .C1(G234), .C2(G237), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT21), .B(G898), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G214), .B1(G237), .B2(G902), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NOR4_X1   g364(.A1(new_n455), .A2(new_n506), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n285), .A2(new_n414), .A3(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(KEYINPUT91), .B(G101), .Z(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(G3));
  INV_X1    g368(.A(G472), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n385), .B2(new_n272), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n394), .ZN(new_n558));
  NOR4_X1   g372(.A1(new_n283), .A2(new_n558), .A3(new_n284), .A4(new_n327), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n531), .A2(new_n532), .A3(new_n538), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT95), .ZN(new_n561));
  INV_X1    g375(.A(new_n529), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n562), .A2(KEYINPUT94), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(KEYINPUT94), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n528), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n565), .B1(new_n528), .B2(new_n529), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT93), .ZN(new_n569));
  OR2_X1    g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n569), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n567), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n532), .A2(G902), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n561), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n455), .ZN(new_n576));
  OAI211_X1 g390(.A(KEYINPUT92), .B(new_n457), .C1(new_n489), .C2(new_n501), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n577), .A2(new_n549), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT92), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n502), .A2(new_n579), .A3(new_n504), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n576), .A2(new_n546), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n559), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT96), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT34), .B(G104), .Z(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(G6));
  NAND2_X1  g400(.A1(new_n446), .A2(new_n447), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT20), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n446), .A2(new_n415), .A3(new_n447), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT86), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n425), .A2(new_n427), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT85), .B1(new_n299), .B2(new_n300), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(new_n438), .A3(new_n436), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n595), .A2(new_n417), .A3(new_n424), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n417), .B1(new_n595), .B2(new_n424), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n272), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n541), .B1(G475), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n590), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n600), .A2(new_n581), .A3(new_n546), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n559), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT35), .B(G107), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G9));
  NOR2_X1   g418(.A1(new_n318), .A2(KEYINPUT36), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n314), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n325), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n324), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n558), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n285), .A2(new_n610), .A3(new_n551), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT37), .B(G110), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G12));
  AOI21_X1  g427(.A(new_n609), .B1(new_n393), .B2(new_n413), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n448), .A2(new_n450), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n539), .A2(new_n540), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(new_n453), .B2(new_n454), .ZN(new_n617));
  INV_X1    g431(.A(G900), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n543), .B1(new_n544), .B2(new_n618), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n615), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n580), .A2(new_n549), .A3(new_n577), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT97), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n619), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n590), .A2(new_n599), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n624), .A2(new_n581), .A3(new_n625), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n285), .B(new_n614), .C1(new_n622), .C2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G128), .ZN(G30));
  XOR2_X1   g442(.A(new_n619), .B(KEYINPUT39), .Z(new_n629));
  NAND2_X1  g443(.A1(new_n285), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n630), .A2(KEYINPUT40), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(KEYINPUT40), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT32), .B1(new_n385), .B2(new_n387), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n382), .A2(new_n383), .ZN(new_n635));
  INV_X1    g449(.A(new_n406), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n363), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n635), .B1(new_n333), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(G472), .B1(new_n638), .B2(G902), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n393), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n455), .A2(new_n616), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n505), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n549), .A3(new_n609), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n641), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n631), .A2(new_n632), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G143), .ZN(G45));
  NAND3_X1  g462(.A1(new_n575), .A2(new_n455), .A3(new_n623), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n581), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n285), .A2(new_n614), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G146), .ZN(G48));
  AOI21_X1  g466(.A(new_n271), .B1(new_n270), .B2(new_n272), .ZN(new_n653));
  AOI211_X1 g467(.A(G469), .B(G902), .C1(new_n265), .C2(new_n269), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n281), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n582), .A2(new_n414), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT41), .B(G113), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G15));
  NAND3_X1  g474(.A1(new_n414), .A2(new_n601), .A3(new_n657), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT99), .B(G116), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G18));
  NAND4_X1  g477(.A1(new_n655), .A2(new_n281), .A3(new_n578), .A4(new_n580), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n664), .A2(new_n455), .A3(new_n548), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n614), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G119), .ZN(G21));
  NOR4_X1   g481(.A1(new_n642), .A2(new_n656), .A3(new_n581), .A4(new_n546), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n409), .A2(new_n402), .A3(new_n401), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT70), .B1(new_n637), .B2(KEYINPUT28), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n333), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n384), .A3(new_n378), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(KEYINPUT100), .A3(new_n387), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT100), .B1(new_n672), .B2(new_n387), .ZN(new_n675));
  NOR4_X1   g489(.A1(new_n674), .A2(new_n675), .A3(new_n556), .A4(new_n327), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n668), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT101), .B(G122), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G24));
  INV_X1    g493(.A(new_n675), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n680), .A2(new_n557), .A3(new_n608), .A4(new_n673), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n681), .A2(new_n649), .A3(new_n664), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n290), .ZN(G27));
  INV_X1    g497(.A(new_n649), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n505), .A2(new_n550), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n279), .A2(new_n281), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n414), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT102), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n689), .A2(new_n693), .A3(new_n690), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n633), .A2(KEYINPUT103), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n385), .A2(new_n390), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n412), .A2(G472), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n633), .A2(KEYINPUT103), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n696), .A2(new_n697), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n327), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n649), .A2(new_n687), .A3(new_n686), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(KEYINPUT42), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n695), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G131), .ZN(G33));
  NAND3_X1  g521(.A1(new_n414), .A2(new_n620), .A3(new_n688), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G134), .ZN(G36));
  NOR3_X1   g523(.A1(new_n267), .A2(new_n268), .A3(new_n266), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n266), .B2(new_n275), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n711), .A2(KEYINPUT45), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(KEYINPUT45), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(G469), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n274), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n273), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n715), .A2(new_n716), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n281), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  INV_X1    g535(.A(new_n629), .ZN(new_n722));
  OR3_X1    g536(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n721), .B1(new_n720), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n726));
  INV_X1    g540(.A(new_n575), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n726), .B1(new_n727), .B2(new_n455), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n727), .A2(new_n726), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n455), .A2(KEYINPUT105), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n455), .A2(KEYINPUT105), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n730), .A2(KEYINPUT106), .A3(new_n731), .A4(new_n732), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n729), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n738), .A2(new_n558), .A3(new_n608), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n725), .B(new_n685), .C1(new_n739), .C2(KEYINPUT44), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(KEYINPUT44), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n741), .A2(KEYINPUT107), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(KEYINPUT107), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n740), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n248), .ZN(G39));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n720), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g561(.A(KEYINPUT47), .B(new_n281), .C1(new_n718), .C2(new_n719), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n393), .A2(new_n413), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n750), .A2(new_n701), .A3(new_n686), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n684), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G140), .ZN(G42));
  INV_X1    g567(.A(new_n681), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n704), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n608), .A2(new_n541), .A3(new_n623), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n686), .A2(new_n455), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n285), .A2(new_n757), .A3(new_n750), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n758), .A3(new_n708), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n759), .B1(new_n695), .B2(new_n705), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n576), .A2(new_n600), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n506), .A2(new_n546), .A3(new_n550), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n559), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n552), .A3(new_n611), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n677), .A2(new_n658), .A3(new_n661), .A4(new_n666), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n760), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n649), .A2(new_n664), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n754), .A2(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n687), .A2(new_n608), .A3(new_n619), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n642), .A2(new_n581), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n773), .A3(new_n640), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n627), .A2(new_n651), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n776), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(new_n775), .B2(new_n777), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n651), .A2(new_n774), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n285), .A2(new_n614), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n625), .B1(new_n624), .B2(new_n581), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n615), .A2(new_n617), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n788), .A2(new_n621), .A3(KEYINPUT97), .A4(new_n623), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n682), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n785), .A2(new_n791), .A3(KEYINPUT110), .A4(KEYINPUT52), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n783), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n780), .A2(new_n781), .A3(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n783), .A2(new_n792), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n787), .A2(new_n789), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT80), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n687), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n750), .A2(new_n798), .A3(new_n282), .A4(new_n608), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n771), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n777), .B1(new_n800), .B2(new_n784), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT111), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT112), .B1(new_n795), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n769), .B1(new_n794), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n775), .B(new_n777), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n766), .A2(KEYINPUT109), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n668), .A2(new_n676), .B1(new_n665), .B2(new_n614), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT109), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n811), .A3(new_n658), .A4(new_n661), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n764), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n808), .A2(new_n813), .A3(new_n760), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n765), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n806), .A2(new_n807), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT113), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n781), .B1(new_n780), .B2(new_n793), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n795), .A2(new_n804), .A3(KEYINPUT112), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n760), .A2(new_n813), .A3(new_n765), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n820), .A2(new_n821), .B1(KEYINPUT53), .B2(new_n814), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT54), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n806), .A2(new_n824), .A3(new_n807), .A4(new_n815), .ZN(new_n825));
  INV_X1    g639(.A(new_n664), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n738), .A2(new_n543), .A3(new_n826), .A4(new_n676), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n657), .A2(new_n685), .ZN(new_n828));
  INV_X1    g642(.A(new_n543), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n828), .A2(new_n640), .A3(new_n327), .A4(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n576), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n542), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n827), .A2(KEYINPUT117), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT117), .B1(new_n827), .B2(new_n832), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT48), .ZN(new_n836));
  NOR4_X1   g650(.A1(new_n737), .A2(new_n829), .A3(new_n702), .A4(new_n828), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n836), .B1(new_n837), .B2(KEYINPUT118), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(KEYINPUT118), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n837), .A2(KEYINPUT118), .A3(new_n836), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n835), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n655), .B(KEYINPUT108), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n747), .B(new_n748), .C1(new_n281), .C2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n737), .A2(new_n829), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(new_n846), .A3(new_n676), .A4(new_n685), .ZN(new_n847));
  INV_X1    g661(.A(new_n455), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n830), .A2(new_n848), .A3(new_n727), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT116), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n846), .A2(new_n657), .A3(new_n754), .A4(new_n685), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n847), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT50), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n644), .B1(KEYINPUT115), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n657), .A2(KEYINPUT114), .A3(new_n550), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n857), .B1(new_n656), .B2(new_n549), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n846), .A2(new_n676), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n854), .A2(KEYINPUT115), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n860), .B(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n853), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n860), .B(new_n861), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT51), .B1(new_n866), .B2(new_n852), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n842), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n817), .A2(new_n823), .A3(new_n825), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT119), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n768), .B1(new_n818), .B2(new_n819), .ZN(new_n871));
  INV_X1    g685(.A(new_n815), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT54), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n873), .A2(new_n824), .B1(new_n822), .B2(KEYINPUT54), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n875), .A3(new_n817), .A4(new_n868), .ZN(new_n876));
  OR2_X1    g690(.A1(G952), .A2(G953), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n870), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n575), .A2(new_n701), .A3(new_n281), .A4(new_n549), .ZN(new_n879));
  AOI211_X1 g693(.A(new_n879), .B(new_n644), .C1(new_n844), .C2(KEYINPUT49), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n732), .A2(new_n731), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n844), .A2(KEYINPUT49), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n880), .A2(new_n641), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n878), .A2(new_n883), .ZN(G75));
  AOI21_X1  g698(.A(new_n272), .B1(new_n806), .B2(new_n815), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(G210), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(new_n492), .ZN(new_n889));
  XOR2_X1   g703(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n890));
  XNOR2_X1  g704(.A(new_n889), .B(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n886), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n886), .B2(new_n887), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n257), .A2(G952), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(G51));
  OAI21_X1  g709(.A(KEYINPUT54), .B1(new_n871), .B2(new_n872), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n816), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n806), .A2(new_n815), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n274), .B(KEYINPUT57), .Z(new_n901));
  NAND3_X1  g715(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n270), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n885), .A2(G469), .A3(new_n713), .A4(new_n712), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n894), .B1(new_n903), .B2(new_n904), .ZN(G54));
  NAND3_X1  g719(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n906));
  INV_X1    g720(.A(new_n446), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n909), .A3(new_n894), .ZN(G60));
  INV_X1    g724(.A(new_n572), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n874), .A2(new_n817), .ZN(new_n912));
  XNOR2_X1  g726(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n532), .A2(new_n272), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n898), .A2(new_n911), .A3(new_n900), .A4(new_n915), .ZN(new_n917));
  INV_X1    g731(.A(new_n894), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n916), .A2(new_n919), .ZN(G63));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT60), .Z(new_n922));
  NAND2_X1  g736(.A1(new_n899), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n320), .B(KEYINPUT123), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n899), .A2(new_n606), .A3(new_n922), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n918), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT61), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(G66));
  INV_X1    g743(.A(G224), .ZN(new_n930));
  OAI21_X1  g744(.A(G953), .B1(new_n545), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n813), .B2(G953), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n888), .B1(G898), .B2(new_n257), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(G69));
  OAI21_X1  g748(.A(new_n371), .B1(new_n375), .B2(KEYINPUT30), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n441), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n800), .B1(new_n786), .B2(new_n650), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n647), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n938), .A2(KEYINPUT62), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n414), .A2(new_n685), .A3(new_n761), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n752), .B1(new_n630), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(KEYINPUT62), .B2(new_n938), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n943), .A2(new_n744), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n936), .B1(new_n944), .B2(new_n257), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n257), .B1(G227), .B2(G900), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n936), .B1(new_n618), .B2(new_n257), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n752), .A2(new_n708), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n725), .A2(new_n773), .A3(new_n703), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n948), .A2(new_n706), .A3(new_n937), .A4(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n744), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n947), .B1(new_n951), .B2(new_n257), .ZN(new_n952));
  OR3_X1    g766(.A1(new_n945), .A2(new_n946), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n946), .B1(new_n945), .B2(new_n952), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(G72));
  XOR2_X1   g769(.A(new_n396), .B(KEYINPUT125), .Z(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n333), .ZN(new_n957));
  INV_X1    g771(.A(new_n813), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n943), .A2(new_n744), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(G472), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT63), .Z(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT124), .Z(new_n962));
  OAI21_X1  g776(.A(new_n957), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n744), .A2(new_n950), .A3(new_n958), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n333), .B(new_n956), .C1(new_n964), .C2(new_n962), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n963), .A2(new_n965), .A3(new_n918), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n382), .A2(new_n383), .A3(new_n397), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n961), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT126), .Z(new_n969));
  AND2_X1   g783(.A1(new_n822), .A2(new_n969), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n970), .A2(KEYINPUT127), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(KEYINPUT127), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n966), .B1(new_n971), .B2(new_n972), .ZN(G57));
endmodule


