

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751;

  XNOR2_X1 U368 ( .A(n551), .B(KEYINPUT107), .ZN(n749) );
  BUF_X1 U369 ( .A(G119), .Z(n346) );
  AND2_X4 U370 ( .A1(n381), .A2(n380), .ZN(n695) );
  INV_X2 U371 ( .A(G953), .ZN(n745) );
  BUF_X1 U372 ( .A(n575), .Z(n617) );
  NOR2_X2 U373 ( .A1(n549), .A2(n511), .ZN(n497) );
  NOR2_X2 U374 ( .A1(n574), .A2(n511), .ZN(n521) );
  NAND2_X1 U375 ( .A1(n378), .A2(n384), .ZN(n381) );
  OR2_X1 U376 ( .A1(n520), .A2(n606), .ZN(n533) );
  XNOR2_X1 U377 ( .A(n456), .B(n455), .ZN(n458) );
  NOR2_X1 U378 ( .A1(G953), .A2(G237), .ZN(n459) );
  XNOR2_X1 U379 ( .A(n352), .B(n507), .ZN(n539) );
  AND2_X1 U380 ( .A1(n371), .A2(n348), .ZN(n362) );
  XNOR2_X1 U381 ( .A(n582), .B(KEYINPUT80), .ZN(n594) );
  OR2_X1 U382 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U383 ( .A(KEYINPUT11), .B(KEYINPUT102), .Z(n434) );
  XOR2_X1 U384 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n432) );
  XNOR2_X1 U385 ( .A(G143), .B(G128), .ZN(n423) );
  AND2_X1 U386 ( .A1(n544), .A2(n552), .ZN(n365) );
  INV_X1 U387 ( .A(KEYINPUT30), .ZN(n570) );
  XNOR2_X1 U388 ( .A(n468), .B(G472), .ZN(n504) );
  XOR2_X1 U389 ( .A(G128), .B(KEYINPUT23), .Z(n472) );
  XNOR2_X1 U390 ( .A(n346), .B(G110), .ZN(n474) );
  NAND2_X1 U391 ( .A1(n622), .A2(n623), .ZN(n382) );
  XNOR2_X1 U392 ( .A(G140), .B(G137), .ZN(n487) );
  XNOR2_X1 U393 ( .A(n358), .B(n357), .ZN(n620) );
  INV_X1 U394 ( .A(KEYINPUT39), .ZN(n357) );
  NAND2_X1 U395 ( .A1(n599), .A2(n646), .ZN(n358) );
  BUF_X1 U396 ( .A(n504), .Z(n635) );
  NAND2_X1 U397 ( .A1(n695), .A2(G472), .ZN(n356) );
  XNOR2_X1 U398 ( .A(n627), .B(KEYINPUT94), .ZN(n703) );
  AND2_X1 U399 ( .A1(n533), .A2(n673), .ZN(n532) );
  INV_X1 U400 ( .A(KEYINPUT72), .ZN(n451) );
  NOR2_X1 U401 ( .A1(n671), .A2(n353), .ZN(n352) );
  INV_X1 U402 ( .A(G237), .ZN(n397) );
  XNOR2_X1 U403 ( .A(G137), .B(G101), .ZN(n462) );
  XOR2_X1 U404 ( .A(G146), .B(KEYINPUT74), .Z(n461) );
  INV_X1 U405 ( .A(KEYINPUT71), .ZN(n427) );
  XNOR2_X1 U406 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n391) );
  XNOR2_X1 U407 ( .A(G146), .B(G125), .ZN(n429) );
  XNOR2_X1 U408 ( .A(n372), .B(n611), .ZN(n371) );
  NAND2_X1 U409 ( .A1(G234), .A2(G237), .ZN(n403) );
  INV_X1 U410 ( .A(G902), .ZN(n479) );
  XNOR2_X1 U411 ( .A(n377), .B(n376), .ZN(n465) );
  XNOR2_X1 U412 ( .A(G116), .B(G113), .ZN(n377) );
  XNOR2_X1 U413 ( .A(KEYINPUT3), .B(G119), .ZN(n376) );
  INV_X1 U414 ( .A(G134), .ZN(n422) );
  XOR2_X1 U415 ( .A(G116), .B(KEYINPUT9), .Z(n417) );
  XNOR2_X1 U416 ( .A(G122), .B(G107), .ZN(n419) );
  INV_X1 U417 ( .A(KEYINPUT7), .ZN(n418) );
  XNOR2_X1 U418 ( .A(G113), .B(G143), .ZN(n437) );
  XNOR2_X1 U419 ( .A(G104), .B(G122), .ZN(n438) );
  XNOR2_X1 U420 ( .A(G140), .B(KEYINPUT101), .ZN(n431) );
  NAND2_X1 U421 ( .A1(n631), .A2(KEYINPUT83), .ZN(n384) );
  XNOR2_X1 U422 ( .A(G110), .B(G107), .ZN(n388) );
  INV_X1 U423 ( .A(G104), .ZN(n387) );
  NAND2_X2 U424 ( .A1(n366), .A2(n363), .ZN(n727) );
  AND2_X1 U425 ( .A1(n365), .A2(n374), .ZN(n364) );
  AND2_X1 U426 ( .A1(n371), .A2(n621), .ZN(n743) );
  AND2_X1 U427 ( .A1(n360), .A2(n359), .ZN(n599) );
  XNOR2_X1 U428 ( .A(n571), .B(n570), .ZN(n572) );
  NOR2_X1 U429 ( .A1(n557), .A2(n568), .ZN(n573) );
  XNOR2_X1 U430 ( .A(n504), .B(n503), .ZN(n569) );
  BUF_X1 U431 ( .A(n511), .Z(n637) );
  XNOR2_X1 U432 ( .A(n375), .B(n489), .ZN(n733) );
  XNOR2_X1 U433 ( .A(n465), .B(n386), .ZN(n375) );
  XNOR2_X1 U434 ( .A(KEYINPUT16), .B(G122), .ZN(n386) );
  XNOR2_X1 U435 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X2 U436 ( .A1(n727), .A2(n743), .ZN(n631) );
  XNOR2_X1 U437 ( .A(n602), .B(n601), .ZN(n750) );
  NOR2_X1 U438 ( .A1(n620), .A2(n600), .ZN(n602) );
  XOR2_X1 U439 ( .A(n514), .B(n513), .Z(n722) );
  NOR2_X1 U440 ( .A1(n641), .A2(n524), .ZN(n513) );
  XNOR2_X1 U441 ( .A(n354), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U442 ( .A1(n355), .A2(n628), .ZN(n354) );
  XNOR2_X1 U443 ( .A(n356), .B(n350), .ZN(n355) );
  XNOR2_X1 U444 ( .A(n510), .B(n509), .ZN(n574) );
  INV_X1 U445 ( .A(n574), .ZN(n359) );
  XOR2_X1 U446 ( .A(n497), .B(n496), .Z(n347) );
  AND2_X1 U447 ( .A1(n621), .A2(n623), .ZN(n348) );
  OR2_X1 U448 ( .A1(KEYINPUT47), .A2(n607), .ZN(n349) );
  XNOR2_X1 U449 ( .A(KEYINPUT15), .B(G902), .ZN(n622) );
  XOR2_X1 U450 ( .A(n626), .B(n625), .Z(n350) );
  AND2_X1 U451 ( .A1(n396), .A2(n383), .ZN(n351) );
  INV_X1 U452 ( .A(KEYINPUT2), .ZN(n383) );
  OR2_X2 U453 ( .A1(n539), .A2(KEYINPUT88), .ZN(n541) );
  INV_X1 U454 ( .A(n672), .ZN(n353) );
  XNOR2_X1 U455 ( .A(n502), .B(n501), .ZN(n671) );
  AND2_X1 U456 ( .A1(n572), .A2(n573), .ZN(n360) );
  NAND2_X1 U457 ( .A1(n361), .A2(n351), .ZN(n379) );
  NAND2_X1 U458 ( .A1(n362), .A2(n727), .ZN(n361) );
  XNOR2_X2 U459 ( .A(n485), .B(KEYINPUT97), .ZN(n739) );
  NAND2_X1 U460 ( .A1(n364), .A2(n543), .ZN(n363) );
  AND2_X2 U461 ( .A1(n369), .A2(n367), .ZN(n366) );
  NAND2_X1 U462 ( .A1(n368), .A2(n373), .ZN(n367) );
  NAND2_X1 U463 ( .A1(n374), .A2(n544), .ZN(n368) );
  NAND2_X1 U464 ( .A1(n370), .A2(n373), .ZN(n369) );
  INV_X1 U465 ( .A(n543), .ZN(n370) );
  NAND2_X1 U466 ( .A1(n609), .A2(n610), .ZN(n372) );
  INV_X1 U467 ( .A(n552), .ZN(n373) );
  INV_X1 U468 ( .A(n749), .ZN(n374) );
  NAND2_X1 U469 ( .A1(n379), .A2(n382), .ZN(n378) );
  INV_X1 U470 ( .A(n624), .ZN(n380) );
  INV_X1 U471 ( .A(n584), .ZN(n557) );
  AND2_X1 U472 ( .A1(n595), .A2(n632), .ZN(n385) );
  INV_X1 U473 ( .A(KEYINPUT89), .ZN(n507) );
  NOR2_X1 U474 ( .A1(n558), .A2(n557), .ZN(n559) );
  INV_X1 U475 ( .A(KEYINPUT24), .ZN(n473) );
  AND2_X1 U476 ( .A1(n560), .A2(n559), .ZN(n561) );
  INV_X1 U477 ( .A(KEYINPUT48), .ZN(n611) );
  XNOR2_X1 U478 ( .A(n419), .B(n418), .ZN(n420) );
  OR2_X1 U479 ( .A1(n518), .A2(n527), .ZN(n600) );
  INV_X1 U480 ( .A(KEYINPUT40), .ZN(n601) );
  XNOR2_X1 U481 ( .A(n387), .B(G101), .ZN(n389) );
  XNOR2_X1 U482 ( .A(n389), .B(n388), .ZN(n489) );
  NAND2_X1 U483 ( .A1(n745), .A2(G224), .ZN(n390) );
  XNOR2_X1 U484 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U485 ( .A(n392), .B(n429), .ZN(n394) );
  XNOR2_X2 U486 ( .A(KEYINPUT69), .B(KEYINPUT4), .ZN(n450) );
  XNOR2_X1 U487 ( .A(n423), .B(n450), .ZN(n393) );
  XNOR2_X1 U488 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U489 ( .A(n733), .B(n395), .ZN(n696) );
  INV_X1 U490 ( .A(n622), .ZN(n396) );
  OR2_X2 U491 ( .A1(n696), .A2(n396), .ZN(n399) );
  NAND2_X1 U492 ( .A1(n479), .A2(n397), .ZN(n400) );
  NAND2_X1 U493 ( .A1(n400), .A2(G210), .ZN(n398) );
  XNOR2_X2 U494 ( .A(n399), .B(n398), .ZN(n575) );
  NAND2_X1 U495 ( .A1(n400), .A2(G214), .ZN(n645) );
  INV_X1 U496 ( .A(n645), .ZN(n401) );
  OR2_X2 U497 ( .A1(n575), .A2(n401), .ZN(n402) );
  XNOR2_X2 U498 ( .A(n402), .B(KEYINPUT19), .ZN(n566) );
  XNOR2_X1 U499 ( .A(n403), .B(KEYINPUT14), .ZN(n407) );
  NAND2_X1 U500 ( .A1(n407), .A2(G952), .ZN(n404) );
  XNOR2_X1 U501 ( .A(n404), .B(KEYINPUT95), .ZN(n660) );
  NAND2_X1 U502 ( .A1(n660), .A2(n745), .ZN(n406) );
  INV_X1 U503 ( .A(KEYINPUT96), .ZN(n405) );
  XNOR2_X1 U504 ( .A(n406), .B(n405), .ZN(n555) );
  AND2_X1 U505 ( .A1(G953), .A2(n407), .ZN(n408) );
  NAND2_X1 U506 ( .A1(G902), .A2(n408), .ZN(n553) );
  NOR2_X1 U507 ( .A1(n553), .A2(G898), .ZN(n409) );
  OR2_X1 U508 ( .A1(n555), .A2(n409), .ZN(n410) );
  NAND2_X1 U509 ( .A1(n566), .A2(n410), .ZN(n413) );
  INV_X1 U510 ( .A(KEYINPUT67), .ZN(n411) );
  XNOR2_X1 U511 ( .A(n411), .B(KEYINPUT0), .ZN(n412) );
  XNOR2_X1 U512 ( .A(n413), .B(n412), .ZN(n512) );
  INV_X1 U513 ( .A(n512), .ZN(n448) );
  XOR2_X1 U514 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n415) );
  NAND2_X1 U515 ( .A1(G234), .A2(n745), .ZN(n414) );
  XNOR2_X1 U516 ( .A(n415), .B(n414), .ZN(n470) );
  NAND2_X1 U517 ( .A1(G217), .A2(n470), .ZN(n416) );
  XNOR2_X1 U518 ( .A(n417), .B(n416), .ZN(n421) );
  XNOR2_X1 U519 ( .A(n421), .B(n420), .ZN(n424) );
  XNOR2_X1 U520 ( .A(n423), .B(n422), .ZN(n457) );
  XNOR2_X1 U521 ( .A(n424), .B(n457), .ZN(n679) );
  AND2_X1 U522 ( .A1(n679), .A2(n479), .ZN(n426) );
  XOR2_X1 U523 ( .A(KEYINPUT104), .B(G478), .Z(n425) );
  XNOR2_X1 U524 ( .A(n426), .B(n425), .ZN(n527) );
  XNOR2_X1 U525 ( .A(n427), .B(G131), .ZN(n455) );
  INV_X1 U526 ( .A(KEYINPUT10), .ZN(n428) );
  XNOR2_X1 U527 ( .A(n429), .B(n428), .ZN(n477) );
  XOR2_X1 U528 ( .A(n455), .B(n477), .Z(n430) );
  XNOR2_X1 U529 ( .A(n430), .B(KEYINPUT100), .ZN(n442) );
  XNOR2_X1 U530 ( .A(n432), .B(n431), .ZN(n436) );
  NAND2_X1 U531 ( .A1(G214), .A2(n459), .ZN(n433) );
  XNOR2_X1 U532 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U533 ( .A(n436), .B(n435), .ZN(n440) );
  XNOR2_X1 U534 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U535 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U536 ( .A(n442), .B(n441), .ZN(n684) );
  NAND2_X1 U537 ( .A1(n684), .A2(n479), .ZN(n444) );
  XNOR2_X1 U538 ( .A(KEYINPUT13), .B(G475), .ZN(n443) );
  XNOR2_X1 U539 ( .A(n444), .B(n443), .ZN(n518) );
  INV_X1 U540 ( .A(n518), .ZN(n526) );
  NOR2_X1 U541 ( .A1(n527), .A2(n526), .ZN(n595) );
  NAND2_X1 U542 ( .A1(n622), .A2(G234), .ZN(n445) );
  XNOR2_X1 U543 ( .A(n445), .B(KEYINPUT20), .ZN(n446) );
  XNOR2_X1 U544 ( .A(KEYINPUT98), .B(n446), .ZN(n480) );
  AND2_X1 U545 ( .A1(n480), .A2(G221), .ZN(n447) );
  XNOR2_X1 U546 ( .A(n447), .B(KEYINPUT21), .ZN(n632) );
  NAND2_X1 U547 ( .A1(n448), .A2(n385), .ZN(n449) );
  XNOR2_X1 U548 ( .A(n449), .B(KEYINPUT22), .ZN(n545) );
  NAND2_X1 U549 ( .A1(n450), .A2(KEYINPUT72), .ZN(n454) );
  INV_X1 U550 ( .A(n450), .ZN(n452) );
  NAND2_X1 U551 ( .A1(n452), .A2(n451), .ZN(n453) );
  NAND2_X1 U552 ( .A1(n454), .A2(n453), .ZN(n456) );
  XNOR2_X2 U553 ( .A(n458), .B(n457), .ZN(n485) );
  NAND2_X1 U554 ( .A1(n459), .A2(G210), .ZN(n460) );
  XNOR2_X1 U555 ( .A(n461), .B(n460), .ZN(n464) );
  XNOR2_X1 U556 ( .A(n462), .B(KEYINPUT5), .ZN(n463) );
  XNOR2_X1 U557 ( .A(n464), .B(n463), .ZN(n466) );
  XNOR2_X1 U558 ( .A(n465), .B(n466), .ZN(n467) );
  XNOR2_X1 U559 ( .A(n485), .B(n467), .ZN(n626) );
  NAND2_X1 U560 ( .A1(n626), .A2(n479), .ZN(n468) );
  INV_X1 U561 ( .A(KEYINPUT6), .ZN(n469) );
  XNOR2_X1 U562 ( .A(n635), .B(n469), .ZN(n587) );
  INV_X1 U563 ( .A(n587), .ZN(n498) );
  NAND2_X1 U564 ( .A1(n470), .A2(G221), .ZN(n471) );
  XNOR2_X1 U565 ( .A(n472), .B(n471), .ZN(n476) );
  XNOR2_X1 U566 ( .A(n476), .B(n475), .ZN(n478) );
  XNOR2_X1 U567 ( .A(n477), .B(n487), .ZN(n737) );
  XNOR2_X1 U568 ( .A(n478), .B(n737), .ZN(n675) );
  NAND2_X1 U569 ( .A1(n675), .A2(n479), .ZN(n483) );
  NAND2_X1 U570 ( .A1(G217), .A2(n480), .ZN(n481) );
  XNOR2_X1 U571 ( .A(KEYINPUT25), .B(n481), .ZN(n482) );
  XNOR2_X2 U572 ( .A(n483), .B(n482), .ZN(n583) );
  INV_X1 U573 ( .A(KEYINPUT106), .ZN(n484) );
  XNOR2_X1 U574 ( .A(n583), .B(n484), .ZN(n549) );
  NAND2_X1 U575 ( .A1(n745), .A2(G227), .ZN(n486) );
  XNOR2_X1 U576 ( .A(n486), .B(G146), .ZN(n488) );
  XNOR2_X1 U577 ( .A(n488), .B(n487), .ZN(n491) );
  INV_X1 U578 ( .A(n489), .ZN(n490) );
  XNOR2_X1 U579 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U580 ( .A(n739), .B(n492), .ZN(n689) );
  OR2_X2 U581 ( .A1(n689), .A2(G902), .ZN(n494) );
  XNOR2_X1 U582 ( .A(KEYINPUT73), .B(G469), .ZN(n493) );
  XNOR2_X2 U583 ( .A(n494), .B(n493), .ZN(n515) );
  XNOR2_X1 U584 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n495) );
  XNOR2_X2 U585 ( .A(n515), .B(n495), .ZN(n511) );
  INV_X1 U586 ( .A(KEYINPUT108), .ZN(n496) );
  NAND2_X1 U587 ( .A1(n498), .A2(n347), .ZN(n499) );
  NOR2_X1 U588 ( .A1(n545), .A2(n499), .ZN(n502) );
  XNOR2_X1 U589 ( .A(KEYINPUT77), .B(KEYINPUT32), .ZN(n500) );
  XNOR2_X1 U590 ( .A(n500), .B(KEYINPUT65), .ZN(n501) );
  INV_X1 U591 ( .A(n583), .ZN(n558) );
  INV_X1 U592 ( .A(KEYINPUT109), .ZN(n503) );
  NOR2_X1 U593 ( .A1(n558), .A2(n569), .ZN(n505) );
  NAND2_X1 U594 ( .A1(n505), .A2(n637), .ZN(n506) );
  OR2_X1 U595 ( .A1(n545), .A2(n506), .ZN(n672) );
  XOR2_X1 U596 ( .A(KEYINPUT31), .B(KEYINPUT99), .Z(n514) );
  INV_X1 U597 ( .A(n632), .ZN(n508) );
  NOR2_X1 U598 ( .A1(n583), .A2(n508), .ZN(n510) );
  INV_X1 U599 ( .A(KEYINPUT68), .ZN(n509) );
  NAND2_X1 U600 ( .A1(n521), .A2(n635), .ZN(n641) );
  BUF_X1 U601 ( .A(n512), .Z(n524) );
  INV_X1 U602 ( .A(n515), .ZN(n562) );
  INV_X1 U603 ( .A(n562), .ZN(n568) );
  NOR2_X1 U604 ( .A1(n568), .A2(n635), .ZN(n516) );
  NAND2_X1 U605 ( .A1(n359), .A2(n516), .ZN(n517) );
  NOR2_X1 U606 ( .A1(n517), .A2(n524), .ZN(n707) );
  NOR2_X1 U607 ( .A1(n722), .A2(n707), .ZN(n520) );
  AND2_X1 U608 ( .A1(n527), .A2(n518), .ZN(n721) );
  INV_X1 U609 ( .A(n721), .ZN(n619) );
  NAND2_X1 U610 ( .A1(n619), .A2(n600), .ZN(n519) );
  XNOR2_X1 U611 ( .A(n519), .B(KEYINPUT105), .ZN(n650) );
  XNOR2_X1 U612 ( .A(n650), .B(KEYINPUT82), .ZN(n606) );
  NAND2_X1 U613 ( .A1(n521), .A2(n587), .ZN(n523) );
  XOR2_X1 U614 ( .A(KEYINPUT110), .B(KEYINPUT33), .Z(n522) );
  XNOR2_X1 U615 ( .A(n523), .B(n522), .ZN(n664) );
  NOR2_X1 U616 ( .A1(n664), .A2(n524), .ZN(n525) );
  XNOR2_X1 U617 ( .A(n525), .B(KEYINPUT34), .ZN(n529) );
  NAND2_X1 U618 ( .A1(n527), .A2(n526), .ZN(n576) );
  XOR2_X1 U619 ( .A(KEYINPUT76), .B(n576), .Z(n528) );
  NAND2_X1 U620 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U621 ( .A(KEYINPUT75), .B(KEYINPUT35), .ZN(n530) );
  XNOR2_X2 U622 ( .A(n531), .B(n530), .ZN(n673) );
  NAND2_X1 U623 ( .A1(n539), .A2(n532), .ZN(n536) );
  INV_X1 U624 ( .A(n533), .ZN(n534) );
  OR2_X1 U625 ( .A1(n534), .A2(KEYINPUT44), .ZN(n535) );
  NAND2_X1 U626 ( .A1(n536), .A2(n535), .ZN(n544) );
  INV_X1 U627 ( .A(KEYINPUT88), .ZN(n537) );
  NOR2_X1 U628 ( .A1(n537), .A2(KEYINPUT44), .ZN(n538) );
  NAND2_X1 U629 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U630 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U631 ( .A1(n542), .A2(n673), .ZN(n543) );
  NOR2_X1 U632 ( .A1(n545), .A2(n587), .ZN(n546) );
  XNOR2_X1 U633 ( .A(KEYINPUT86), .B(n546), .ZN(n547) );
  NAND2_X1 U634 ( .A1(n547), .A2(n637), .ZN(n548) );
  XNOR2_X1 U635 ( .A(n548), .B(KEYINPUT87), .ZN(n550) );
  NAND2_X1 U636 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U637 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n552) );
  AND2_X1 U638 ( .A1(n632), .A2(n569), .ZN(n560) );
  NOR2_X1 U639 ( .A1(G900), .A2(n553), .ZN(n554) );
  XNOR2_X1 U640 ( .A(KEYINPUT112), .B(n554), .ZN(n556) );
  OR2_X1 U641 ( .A1(n556), .A2(n555), .ZN(n584) );
  XNOR2_X1 U642 ( .A(n561), .B(KEYINPUT28), .ZN(n563) );
  AND2_X1 U643 ( .A1(n563), .A2(n562), .ZN(n565) );
  INV_X1 U644 ( .A(KEYINPUT115), .ZN(n564) );
  XNOR2_X1 U645 ( .A(n565), .B(n564), .ZN(n597) );
  NAND2_X1 U646 ( .A1(n597), .A2(n566), .ZN(n605) );
  NAND2_X1 U647 ( .A1(n605), .A2(KEYINPUT47), .ZN(n567) );
  XNOR2_X1 U648 ( .A(n567), .B(KEYINPUT81), .ZN(n581) );
  NAND2_X1 U649 ( .A1(KEYINPUT47), .A2(n650), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n569), .A2(n645), .ZN(n571) );
  NOR2_X1 U651 ( .A1(n576), .A2(n617), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n599), .A2(n577), .ZN(n715) );
  NAND2_X1 U653 ( .A1(n578), .A2(n715), .ZN(n579) );
  XNOR2_X1 U654 ( .A(KEYINPUT78), .B(n579), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n583), .A2(n632), .ZN(n589) );
  XOR2_X1 U656 ( .A(KEYINPUT111), .B(n600), .Z(n716) );
  NAND2_X1 U657 ( .A1(n645), .A2(n584), .ZN(n585) );
  NOR2_X1 U658 ( .A1(n716), .A2(n585), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U660 ( .A1(n589), .A2(n588), .ZN(n612) );
  INV_X1 U661 ( .A(n617), .ZN(n590) );
  AND2_X1 U662 ( .A1(n612), .A2(n590), .ZN(n592) );
  XNOR2_X1 U663 ( .A(KEYINPUT36), .B(KEYINPUT90), .ZN(n591) );
  XNOR2_X1 U664 ( .A(n592), .B(n591), .ZN(n593) );
  INV_X1 U665 ( .A(n637), .ZN(n613) );
  AND2_X1 U666 ( .A1(n593), .A2(n613), .ZN(n724) );
  NOR2_X1 U667 ( .A1(n594), .A2(n724), .ZN(n610) );
  INV_X1 U668 ( .A(n595), .ZN(n648) );
  XNOR2_X1 U669 ( .A(n617), .B(KEYINPUT38), .ZN(n646) );
  NAND2_X1 U670 ( .A1(n646), .A2(n645), .ZN(n651) );
  NOR2_X1 U671 ( .A1(n648), .A2(n651), .ZN(n596) );
  XOR2_X1 U672 ( .A(KEYINPUT41), .B(n596), .Z(n662) );
  NAND2_X1 U673 ( .A1(n662), .A2(n597), .ZN(n598) );
  XNOR2_X1 U674 ( .A(KEYINPUT42), .B(n598), .ZN(n751) );
  NAND2_X1 U675 ( .A1(n751), .A2(n750), .ZN(n604) );
  XNOR2_X1 U676 ( .A(KEYINPUT46), .B(KEYINPUT85), .ZN(n603) );
  XNOR2_X1 U677 ( .A(n604), .B(n603), .ZN(n608) );
  OR2_X1 U678 ( .A1(n605), .A2(n606), .ZN(n607) );
  AND2_X1 U679 ( .A1(n608), .A2(n349), .ZN(n609) );
  XNOR2_X1 U680 ( .A(KEYINPUT113), .B(n612), .ZN(n614) );
  NOR2_X1 U681 ( .A1(n614), .A2(n613), .ZN(n616) );
  XOR2_X1 U682 ( .A(KEYINPUT114), .B(KEYINPUT43), .Z(n615) );
  XNOR2_X1 U683 ( .A(n616), .B(n615), .ZN(n618) );
  NAND2_X1 U684 ( .A1(n618), .A2(n617), .ZN(n629) );
  OR2_X1 U685 ( .A1(n620), .A2(n619), .ZN(n726) );
  AND2_X1 U686 ( .A1(n629), .A2(n726), .ZN(n621) );
  INV_X1 U687 ( .A(KEYINPUT83), .ZN(n623) );
  NOR2_X1 U688 ( .A1(n631), .A2(n383), .ZN(n624) );
  XOR2_X1 U689 ( .A(KEYINPUT92), .B(KEYINPUT62), .Z(n625) );
  NOR2_X1 U690 ( .A1(n745), .A2(G952), .ZN(n627) );
  INV_X1 U691 ( .A(n703), .ZN(n628) );
  XNOR2_X1 U692 ( .A(n629), .B(G140), .ZN(G42) );
  XNOR2_X1 U693 ( .A(KEYINPUT2), .B(KEYINPUT84), .ZN(n630) );
  XNOR2_X1 U694 ( .A(n631), .B(n630), .ZN(n669) );
  NOR2_X1 U695 ( .A1(n549), .A2(n632), .ZN(n633) );
  XOR2_X1 U696 ( .A(KEYINPUT49), .B(n633), .Z(n634) );
  NOR2_X1 U697 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U698 ( .A(KEYINPUT118), .B(n636), .ZN(n640) );
  NAND2_X1 U699 ( .A1(n574), .A2(n637), .ZN(n638) );
  XNOR2_X1 U700 ( .A(n638), .B(KEYINPUT50), .ZN(n639) );
  NAND2_X1 U701 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U702 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U703 ( .A(KEYINPUT51), .B(n643), .Z(n644) );
  NAND2_X1 U704 ( .A1(n644), .A2(n662), .ZN(n657) );
  INV_X1 U705 ( .A(n664), .ZN(n655) );
  NOR2_X1 U706 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U707 ( .A(n647), .B(KEYINPUT119), .ZN(n649) );
  NAND2_X1 U708 ( .A1(n649), .A2(n595), .ZN(n653) );
  OR2_X1 U709 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U710 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U711 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U712 ( .A1(n657), .A2(n656), .ZN(n659) );
  XOR2_X1 U713 ( .A(KEYINPUT52), .B(KEYINPUT120), .Z(n658) );
  XOR2_X1 U714 ( .A(n659), .B(n658), .Z(n661) );
  NAND2_X1 U715 ( .A1(n661), .A2(n660), .ZN(n667) );
  INV_X1 U716 ( .A(n662), .ZN(n663) );
  NOR2_X1 U717 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U718 ( .A1(n665), .A2(G953), .ZN(n666) );
  NAND2_X1 U719 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U720 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U721 ( .A(n670), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U722 ( .A(n671), .B(n346), .Z(G21) );
  XNOR2_X1 U723 ( .A(n672), .B(G110), .ZN(G12) );
  XNOR2_X1 U724 ( .A(n673), .B(G122), .ZN(G24) );
  NAND2_X1 U725 ( .A1(n695), .A2(G217), .ZN(n677) );
  XNOR2_X1 U726 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n674) );
  XNOR2_X1 U727 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U728 ( .A(n677), .B(n676), .ZN(n678) );
  NOR2_X1 U729 ( .A1(n678), .A2(n703), .ZN(G66) );
  NAND2_X1 U730 ( .A1(n695), .A2(G478), .ZN(n681) );
  XOR2_X1 U731 ( .A(KEYINPUT122), .B(n679), .Z(n680) );
  XNOR2_X1 U732 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U733 ( .A1(n682), .A2(n703), .ZN(G63) );
  NAND2_X1 U734 ( .A1(n695), .A2(G475), .ZN(n686) );
  XOR2_X1 U735 ( .A(KEYINPUT93), .B(KEYINPUT59), .Z(n683) );
  XNOR2_X1 U736 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U737 ( .A(n686), .B(n685), .ZN(n687) );
  NOR2_X1 U738 ( .A1(n687), .A2(n703), .ZN(n688) );
  XNOR2_X1 U739 ( .A(n688), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U740 ( .A1(n695), .A2(G469), .ZN(n693) );
  XNOR2_X1 U741 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n690) );
  XNOR2_X1 U742 ( .A(n690), .B(KEYINPUT58), .ZN(n691) );
  XNOR2_X1 U743 ( .A(n689), .B(n691), .ZN(n692) );
  XNOR2_X1 U744 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U745 ( .A1(n694), .A2(n703), .ZN(G54) );
  NAND2_X1 U746 ( .A1(n695), .A2(G210), .ZN(n702) );
  BUF_X1 U747 ( .A(n696), .Z(n700) );
  XOR2_X1 U748 ( .A(KEYINPUT79), .B(KEYINPUT91), .Z(n698) );
  XNOR2_X1 U749 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n697) );
  XNOR2_X1 U750 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U751 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U752 ( .A(n702), .B(n701), .ZN(n704) );
  NOR2_X1 U753 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U754 ( .A(n705), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U755 ( .A(n716), .ZN(n718) );
  NAND2_X1 U756 ( .A1(n707), .A2(n718), .ZN(n706) );
  XNOR2_X1 U757 ( .A(n706), .B(G104), .ZN(G6) );
  XNOR2_X1 U758 ( .A(G107), .B(KEYINPUT116), .ZN(n711) );
  XOR2_X1 U759 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n709) );
  NAND2_X1 U760 ( .A1(n707), .A2(n721), .ZN(n708) );
  XNOR2_X1 U761 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U762 ( .A(n711), .B(n710), .ZN(G9) );
  XOR2_X1 U763 ( .A(G128), .B(KEYINPUT29), .Z(n714) );
  INV_X1 U764 ( .A(n605), .ZN(n712) );
  NAND2_X1 U765 ( .A1(n712), .A2(n721), .ZN(n713) );
  XNOR2_X1 U766 ( .A(n714), .B(n713), .ZN(G30) );
  XNOR2_X1 U767 ( .A(G143), .B(n715), .ZN(G45) );
  OR2_X1 U768 ( .A1(n605), .A2(n716), .ZN(n717) );
  XNOR2_X1 U769 ( .A(n717), .B(G146), .ZN(G48) );
  XOR2_X1 U770 ( .A(G113), .B(KEYINPUT117), .Z(n720) );
  NAND2_X1 U771 ( .A1(n722), .A2(n718), .ZN(n719) );
  XNOR2_X1 U772 ( .A(n720), .B(n719), .ZN(G15) );
  NAND2_X1 U773 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U774 ( .A(n723), .B(G116), .ZN(G18) );
  XNOR2_X1 U775 ( .A(n724), .B(G125), .ZN(n725) );
  XNOR2_X1 U776 ( .A(n725), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U777 ( .A(G134), .B(n726), .ZN(G36) );
  NAND2_X1 U778 ( .A1(n727), .A2(n745), .ZN(n731) );
  NAND2_X1 U779 ( .A1(G953), .A2(G224), .ZN(n728) );
  XNOR2_X1 U780 ( .A(KEYINPUT61), .B(n728), .ZN(n729) );
  NAND2_X1 U781 ( .A1(n729), .A2(G898), .ZN(n730) );
  NAND2_X1 U782 ( .A1(n731), .A2(n730), .ZN(n736) );
  OR2_X1 U783 ( .A1(G898), .A2(n745), .ZN(n732) );
  NAND2_X1 U784 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U785 ( .A(n734), .B(KEYINPUT125), .ZN(n735) );
  XNOR2_X1 U786 ( .A(n736), .B(n735), .ZN(G69) );
  XNOR2_X1 U787 ( .A(n737), .B(KEYINPUT126), .ZN(n738) );
  XNOR2_X1 U788 ( .A(n739), .B(n738), .ZN(n744) );
  XOR2_X1 U789 ( .A(G227), .B(n744), .Z(n740) );
  NAND2_X1 U790 ( .A1(n740), .A2(G900), .ZN(n741) );
  NAND2_X1 U791 ( .A1(n741), .A2(G953), .ZN(n742) );
  XOR2_X1 U792 ( .A(KEYINPUT127), .B(n742), .Z(n748) );
  XNOR2_X1 U793 ( .A(n744), .B(n743), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n748), .A2(n747), .ZN(G72) );
  XOR2_X1 U796 ( .A(G101), .B(n749), .Z(G3) );
  XNOR2_X1 U797 ( .A(n750), .B(G131), .ZN(G33) );
  XNOR2_X1 U798 ( .A(G137), .B(n751), .ZN(G39) );
endmodule

