//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1157, new_n1158, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n454), .A2(new_n458), .B1(new_n449), .B2(new_n455), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT66), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n465), .A2(new_n468), .B1(G101), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n472), .B1(new_n463), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT67), .B(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n471), .A2(new_n476), .ZN(G160));
  XNOR2_X1  g052(.A(new_n463), .B(KEYINPUT68), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n469), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n478), .A2(new_n475), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n468), .C2(G112), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n481), .A2(new_n484), .A3(new_n485), .ZN(G162));
  OAI21_X1  g061(.A(G138), .B1(new_n461), .B2(new_n462), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT4), .B1(new_n487), .B2(new_n475), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(KEYINPUT3), .B(G2104), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n468), .A2(new_n491), .A3(new_n492), .A4(G138), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  INV_X1    g071(.A(new_n462), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n499), .A2(KEYINPUT70), .A3(new_n492), .A4(new_n468), .ZN(new_n500));
  OAI211_X1 g075(.A(KEYINPUT69), .B(KEYINPUT4), .C1(new_n487), .C2(new_n475), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n490), .A2(new_n495), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n469), .A2(G114), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n491), .A2(new_n503), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT72), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(new_n512), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n520), .A2(KEYINPUT71), .A3(G50), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  INV_X1    g100(.A(new_n519), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n510), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n523), .A2(new_n524), .B1(new_n528), .B2(G88), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n514), .A2(new_n529), .ZN(G166));
  NAND2_X1  g105(.A1(new_n520), .A2(G51), .ZN(new_n531));
  XOR2_X1   g106(.A(KEYINPUT73), .B(G89), .Z(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n533), .A2(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(new_n520), .A2(G52), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n527), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n512), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(G171));
  NAND2_X1  g119(.A1(new_n520), .A2(G43), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n527), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n512), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g127(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n553));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND3_X1  g131(.A1(new_n520), .A2(KEYINPUT75), .A3(G53), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT9), .Z(new_n558));
  AOI22_X1  g133(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n559), .A2(new_n512), .B1(new_n527), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND2_X1  g140(.A1(new_n514), .A2(new_n529), .ZN(G303));
  NAND2_X1  g141(.A1(new_n528), .A2(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n520), .A2(G49), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  NAND2_X1  g145(.A1(new_n520), .A2(G48), .ZN(new_n571));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n527), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n510), .A2(G61), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n512), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G305));
  NAND2_X1  g153(.A1(new_n520), .A2(G47), .ZN(new_n579));
  INV_X1    g154(.A(G85), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n527), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n512), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  INV_X1    g161(.A(G92), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n527), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT10), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n510), .A2(G66), .ZN(new_n590));
  INV_X1    g165(.A(G79), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n516), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(G54), .B2(new_n520), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n586), .B1(new_n594), .B2(G868), .ZN(G321));
  XOR2_X1   g170(.A(G321), .B(KEYINPUT76), .Z(G284));
  NAND2_X1  g171(.A1(G286), .A2(G868), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n562), .B2(G868), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(new_n562), .B2(G868), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n594), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n594), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI221_X1 g180(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n468), .C2(G111), .ZN(new_n606));
  INV_X1    g181(.A(G123), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n482), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(G135), .B2(new_n480), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT77), .Z(new_n610));
  XOR2_X1   g185(.A(KEYINPUT78), .B(G2096), .Z(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n491), .A2(new_n470), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(G156));
  XNOR2_X1  g192(.A(KEYINPUT15), .B(G2435), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT79), .B(G2438), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(G2427), .B(G2430), .Z(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n622), .A2(KEYINPUT14), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2451), .B(G2454), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n624), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  AND3_X1   g207(.A1(new_n631), .A2(new_n632), .A3(G14), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT80), .Z(G401));
  INV_X1    g209(.A(KEYINPUT18), .ZN(new_n635));
  XOR2_X1   g210(.A(G2084), .B(G2090), .Z(new_n636));
  XNOR2_X1  g211(.A(G2067), .B(G2678), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT17), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n636), .A2(new_n637), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n635), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n638), .B2(KEYINPUT18), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2096), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(G227));
  XOR2_X1   g221(.A(G1971), .B(G1976), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT19), .ZN(new_n648));
  XOR2_X1   g223(.A(G1956), .B(G2474), .Z(new_n649));
  XOR2_X1   g224(.A(G1961), .B(G1966), .Z(new_n650));
  AND2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT20), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n649), .A2(new_n650), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n648), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n648), .B2(new_n654), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n657), .B(new_n658), .Z(new_n659));
  XNOR2_X1  g234(.A(G1991), .B(G1996), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1981), .B(G1986), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G229));
  INV_X1    g239(.A(G16), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G22), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(G166), .B2(new_n665), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT83), .Z(new_n668));
  INV_X1    g243(.A(G1971), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(KEYINPUT83), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G1971), .ZN(new_n672));
  NOR2_X1   g247(.A1(G6), .A2(G16), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n577), .B2(G16), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT32), .ZN(new_n675));
  INV_X1    g250(.A(G1981), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n665), .A2(G23), .ZN(new_n678));
  INV_X1    g253(.A(G288), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(new_n665), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT82), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT33), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND4_X1  g258(.A1(new_n670), .A2(new_n672), .A3(new_n677), .A4(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n684), .A2(KEYINPUT34), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(KEYINPUT34), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n483), .A2(G119), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n468), .A2(G107), .ZN(new_n688));
  OAI21_X1  g263(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT81), .ZN(new_n690));
  AND3_X1   g265(.A1(new_n480), .A2(new_n690), .A3(G131), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(new_n480), .B2(G131), .ZN(new_n692));
  OAI221_X1 g267(.A(new_n687), .B1(new_n688), .B2(new_n689), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(G25), .B(new_n693), .S(G29), .Z(new_n694));
  XOR2_X1   g269(.A(KEYINPUT35), .B(G1991), .Z(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n694), .A2(new_n696), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n665), .A2(G24), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n584), .B2(new_n665), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1986), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g277(.A1(new_n685), .A2(new_n686), .A3(new_n697), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT36), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G33), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT86), .B(KEYINPUT25), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT87), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(G115), .A2(G2104), .ZN(new_n711));
  INV_X1    g286(.A(G127), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n463), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n710), .B1(new_n475), .B2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G139), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n479), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n706), .B1(new_n717), .B2(new_n705), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G2072), .ZN(new_n719));
  INV_X1    g294(.A(G35), .ZN(new_n720));
  OR3_X1    g295(.A1(new_n720), .A2(KEYINPUT93), .A3(G29), .ZN(new_n721));
  OAI21_X1  g296(.A(KEYINPUT93), .B1(new_n720), .B2(G29), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n721), .B(new_n722), .C1(G162), .C2(new_n705), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT29), .B(G2090), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n665), .A2(G19), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n550), .B2(new_n665), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT84), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1341), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n665), .A2(G4), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n594), .B2(new_n665), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(G1348), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n665), .A2(G20), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT94), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT23), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n562), .B2(new_n665), .ZN(new_n737));
  INV_X1    g312(.A(G1956), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n705), .A2(G26), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT85), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  OAI221_X1 g318(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n468), .C2(G116), .ZN(new_n744));
  INV_X1    g319(.A(G140), .ZN(new_n745));
  INV_X1    g320(.A(G128), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n744), .B1(new_n479), .B2(new_n745), .C1(new_n746), .C2(new_n482), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n743), .B1(new_n747), .B2(G29), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2067), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n665), .A2(G5), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G171), .B2(new_n665), .ZN(new_n751));
  INV_X1    g326(.A(G1961), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G34), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(KEYINPUT24), .ZN(new_n755));
  AOI21_X1  g330(.A(G29), .B1(new_n754), .B2(KEYINPUT24), .ZN(new_n756));
  AOI22_X1  g331(.A1(G160), .A2(G29), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(G2084), .ZN(new_n758));
  INV_X1    g333(.A(G1966), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n665), .A2(G21), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G168), .B2(new_n665), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n758), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n757), .A2(G2084), .B1(new_n761), .B2(G1966), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n749), .A2(new_n753), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n719), .A2(new_n730), .A3(new_n740), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT27), .B(G1996), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n480), .A2(G141), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n483), .A2(G129), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT26), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n773), .A2(new_n774), .B1(G105), .B2(new_n470), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n769), .A2(new_n770), .A3(new_n775), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT88), .Z(new_n777));
  MUX2_X1   g352(.A(G32), .B(new_n777), .S(G29), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT89), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n766), .B1(new_n768), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT31), .B(G11), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT90), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT30), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n783), .A2(G28), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n705), .B1(new_n783), .B2(G28), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n782), .B1(new_n784), .B2(new_n785), .C1(new_n610), .C2(new_n705), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT91), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n705), .A2(G27), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G164), .B2(new_n705), .ZN(new_n789));
  INV_X1    g364(.A(G2078), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(KEYINPUT92), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(KEYINPUT92), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n787), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n780), .B(new_n794), .C1(new_n768), .C2(new_n779), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n704), .A2(new_n795), .ZN(G311));
  NAND2_X1  g371(.A1(new_n704), .A2(new_n795), .ZN(G150));
  XNOR2_X1  g372(.A(KEYINPUT95), .B(G55), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n520), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G93), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n801));
  OAI221_X1 g376(.A(new_n799), .B1(new_n527), .B2(new_n800), .C1(new_n801), .C2(new_n512), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G860), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT37), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n594), .A2(G559), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT38), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n802), .B1(new_n550), .B2(KEYINPUT96), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT97), .B1(new_n550), .B2(KEYINPUT96), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT96), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT97), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n809), .B(new_n810), .C1(new_n547), .C2(new_n549), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n807), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n807), .B1(new_n808), .B2(new_n811), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n806), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n817), .A2(KEYINPUT39), .ZN(new_n818));
  INV_X1    g393(.A(G860), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n817), .B2(KEYINPUT39), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n804), .B1(new_n818), .B2(new_n820), .ZN(G145));
  NAND2_X1  g396(.A1(new_n483), .A2(G130), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT100), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n480), .A2(G142), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT99), .ZN(new_n825));
  OR3_X1    g400(.A1(new_n468), .A2(KEYINPUT101), .A3(G118), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT101), .B1(new_n468), .B2(G118), .ZN(new_n827));
  OR2_X1    g402(.A1(G106), .A2(G2105), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n826), .A2(G2104), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n823), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n747), .B(new_n508), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n693), .B(new_n614), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n835), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n837), .A2(new_n833), .A3(new_n832), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n777), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n717), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n716), .A2(new_n776), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n836), .A2(new_n842), .A3(new_n843), .A4(new_n838), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n610), .B(G160), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G162), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G37), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n849), .A2(new_n845), .A3(new_n846), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g430(.A1(G166), .A2(G290), .ZN(new_n856));
  NAND2_X1  g431(.A1(G303), .A2(new_n584), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(G288), .B(new_n577), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT42), .ZN(new_n861));
  INV_X1    g436(.A(new_n859), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n856), .A2(new_n862), .A3(new_n857), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n865));
  INV_X1    g440(.A(new_n863), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n862), .B1(new_n856), .B2(new_n857), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n860), .A2(KEYINPUT104), .A3(new_n863), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n864), .B1(new_n870), .B2(new_n861), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT105), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n602), .B(KEYINPUT102), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n873), .A2(new_n815), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n815), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n589), .A2(new_n593), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT103), .B1(new_n562), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(G299), .A2(new_n594), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n562), .A2(new_n877), .A3(KEYINPUT103), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT41), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n879), .A2(new_n884), .A3(new_n880), .A4(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n876), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(new_n882), .B2(new_n876), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n889), .B(new_n864), .C1(new_n870), .C2(new_n861), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n872), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(G868), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n888), .B1(new_n872), .B2(new_n890), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n892), .A2(KEYINPUT106), .A3(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n896));
  INV_X1    g471(.A(G868), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n896), .B1(new_n802), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n894), .B1(new_n895), .B2(new_n898), .ZN(G295));
  AOI21_X1  g474(.A(new_n894), .B1(new_n895), .B2(new_n898), .ZN(G331));
  XNOR2_X1  g475(.A(G171), .B(G168), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n813), .B2(new_n814), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n808), .A2(new_n811), .ZN(new_n904));
  INV_X1    g479(.A(new_n807), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(new_n812), .A3(new_n901), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n903), .A2(KEYINPUT107), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n909), .B(new_n902), .C1(new_n813), .C2(new_n814), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n883), .A2(new_n908), .A3(new_n885), .A4(new_n910), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n903), .A2(new_n907), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n882), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n870), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n868), .A2(new_n869), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(new_n911), .A3(new_n913), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n915), .A2(new_n916), .A3(new_n852), .A4(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n919), .A2(KEYINPUT44), .ZN(new_n920));
  INV_X1    g495(.A(new_n882), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(new_n908), .B2(new_n910), .ZN(new_n922));
  OAI22_X1  g497(.A1(new_n922), .A2(KEYINPUT108), .B1(new_n886), .B2(new_n912), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n922), .A2(KEYINPUT108), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n870), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n918), .A2(new_n852), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n920), .B(KEYINPUT110), .C1(new_n928), .C2(new_n916), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n916), .B1(new_n925), .B2(new_n927), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n919), .A2(KEYINPUT44), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n925), .A2(new_n927), .A3(new_n916), .ZN(new_n935));
  INV_X1    g510(.A(new_n915), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT43), .B1(new_n936), .B2(new_n926), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n938), .A2(KEYINPUT109), .A3(new_n939), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n934), .A2(new_n942), .A3(new_n943), .ZN(G397));
  INV_X1    g519(.A(G1384), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n508), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g521(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n471), .A2(G40), .A3(new_n476), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  OR3_X1    g527(.A1(new_n952), .A2(G1986), .A3(G290), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(G1986), .A3(G290), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT112), .Z(new_n956));
  INV_X1    g531(.A(G2067), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n747), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n776), .A2(G1996), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n958), .B(new_n959), .C1(new_n777), .C2(G1996), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n693), .B(new_n696), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n951), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n956), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(G1384), .B1(new_n502), .B2(new_n507), .ZN(new_n964));
  INV_X1    g539(.A(new_n947), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n949), .B1(new_n964), .B2(KEYINPUT45), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n759), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n950), .B1(new_n946), .B2(KEYINPUT50), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n964), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n969), .B(G168), .C1(new_n973), .C2(G2084), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(G8), .ZN(new_n975));
  INV_X1    g550(.A(new_n972), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n949), .B1(new_n964), .B2(new_n971), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G2084), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G168), .B1(new_n980), .B2(new_n969), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT51), .B1(new_n975), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n974), .A2(new_n983), .A3(G8), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT126), .ZN(new_n987));
  XNOR2_X1  g562(.A(KEYINPUT114), .B(G1971), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(G1384), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n502), .B2(new_n507), .ZN(new_n992));
  OAI22_X1  g567(.A1(KEYINPUT113), .A2(new_n992), .B1(new_n964), .B2(new_n965), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n508), .A2(KEYINPUT113), .A3(new_n990), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n949), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n988), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G2090), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n970), .A2(new_n997), .A3(new_n972), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(G8), .ZN(new_n1000));
  INV_X1    g575(.A(G8), .ZN(new_n1001));
  AND2_X1   g576(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1002));
  NOR2_X1   g577(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR3_X1   g579(.A1(G166), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1002), .B1(G303), .B2(G8), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1000), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1001), .B1(new_n996), .B2(new_n998), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1007), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n1012));
  INV_X1    g587(.A(new_n573), .ZN(new_n1013));
  INV_X1    g588(.A(new_n576), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n676), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n573), .A2(new_n576), .A3(G1981), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1012), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT49), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1001), .B1(new_n964), .B2(new_n949), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1012), .B(new_n1020), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n679), .A2(G1976), .ZN(new_n1023));
  INV_X1    g598(.A(G1976), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT52), .B1(G288), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1019), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  AND4_X1   g605(.A1(new_n987), .A2(new_n1008), .A3(new_n1011), .A4(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1026), .B(new_n1022), .C1(new_n1032), .C2(new_n1028), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n987), .B1(new_n1034), .B2(new_n1011), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n966), .B(new_n949), .C1(KEYINPUT45), .C2(new_n964), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(G2078), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1961), .B1(new_n970), .B2(new_n972), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT123), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n752), .B1(new_n976), .B2(new_n977), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT123), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1044), .B(new_n1045), .C1(new_n1037), .C2(new_n1040), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n508), .A2(new_n990), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT113), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n950), .B1(new_n992), .B2(KEYINPUT113), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n948), .A2(new_n1050), .A3(new_n1051), .A4(new_n790), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n1038), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1052), .A2(KEYINPUT124), .A3(new_n1038), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(G301), .B1(new_n1047), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n986), .A2(new_n1036), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n562), .B(KEYINPUT57), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT56), .B(G2072), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n948), .A2(new_n1050), .A3(new_n1051), .A4(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1064), .A2(new_n1065), .B1(new_n978), .B2(G1956), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n993), .A2(new_n995), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT118), .B1(new_n1067), .B2(new_n1063), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1062), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(KEYINPUT118), .A3(new_n1063), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n973), .A2(new_n738), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1070), .A2(new_n1071), .A3(new_n1061), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1348), .B1(new_n970), .B2(new_n972), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n964), .A2(new_n949), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(G2067), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n594), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1069), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT61), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT122), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n1083));
  AOI211_X1 g658(.A(new_n1083), .B(KEYINPUT61), .C1(new_n1069), .C2(new_n1073), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1069), .A2(KEYINPUT61), .A3(new_n1073), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n948), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT119), .B1(new_n1087), .B2(G1996), .ZN(new_n1088));
  INV_X1    g663(.A(new_n993), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n1090));
  INV_X1    g665(.A(G1996), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .A4(new_n1051), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1093));
  XNOR2_X1  g668(.A(new_n1093), .B(G1341), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1076), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1088), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n550), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1077), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n877), .B(new_n1100), .C1(new_n978), .C2(G1348), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1078), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n877), .A2(KEYINPUT60), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1102), .A2(KEYINPUT60), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1096), .A2(new_n1106), .A3(KEYINPUT59), .A4(new_n550), .ZN(new_n1107));
  AND4_X1   g682(.A1(new_n1086), .A2(new_n1099), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1079), .B1(new_n1085), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1056), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT124), .B1(new_n1052), .B2(new_n1038), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1087), .B2(new_n1040), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1067), .A2(KEYINPUT125), .A3(new_n1039), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(new_n1116), .A3(new_n1044), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1113), .A2(new_n1117), .A3(G171), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1110), .B1(new_n1118), .B2(new_n1058), .ZN(new_n1119));
  OAI21_X1  g694(.A(G171), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1047), .A2(new_n1057), .A3(G301), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(new_n1121), .A3(KEYINPUT54), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1036), .A2(new_n1119), .A3(new_n985), .A4(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1060), .B1(new_n1109), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1022), .A2(new_n1024), .A3(new_n679), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(G1981), .B2(G305), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1019), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1011), .B2(new_n1033), .ZN(new_n1128));
  AOI211_X1 g703(.A(new_n1001), .B(G286), .C1(new_n980), .C2(new_n969), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1008), .A2(new_n1129), .A3(new_n1011), .A4(new_n1030), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT63), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1034), .A2(KEYINPUT63), .A3(new_n1011), .A4(new_n1129), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1128), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(KEYINPUT117), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1136), .B(new_n1128), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n963), .B1(new_n1124), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n958), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n951), .B1(new_n1140), .B2(new_n776), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n952), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT46), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1143), .B1(new_n951), .B2(new_n1091), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1141), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT47), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT48), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n953), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n953), .A2(new_n1147), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(new_n962), .A3(new_n1149), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n960), .A2(new_n693), .A3(new_n696), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n747), .A2(G2067), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n951), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1146), .A2(new_n1150), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1139), .A2(new_n1154), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g730(.A(G319), .ZN(new_n1157));
  NOR3_X1   g731(.A1(new_n633), .A2(new_n1157), .A3(G227), .ZN(new_n1158));
  NAND2_X1  g732(.A1(new_n663), .A2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g733(.A(new_n1159), .B(KEYINPUT127), .ZN(new_n1160));
  AND3_X1   g734(.A1(new_n1160), .A2(new_n854), .A3(new_n938), .ZN(G308));
  NAND3_X1  g735(.A1(new_n1160), .A2(new_n854), .A3(new_n938), .ZN(G225));
endmodule


