

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589;

  NAND2_X1 U321 ( .A1(n472), .A2(n471), .ZN(n487) );
  NOR2_X1 U322 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U323 ( .A(n354), .B(n353), .ZN(n357) );
  XNOR2_X1 U324 ( .A(KEYINPUT101), .B(KEYINPUT37), .ZN(n490) );
  XOR2_X1 U325 ( .A(n308), .B(n307), .Z(n531) );
  XOR2_X1 U326 ( .A(G211GAT), .B(G218GAT), .Z(n289) );
  XOR2_X1 U327 ( .A(KEYINPUT40), .B(n501), .Z(n290) );
  NOR2_X1 U328 ( .A1(n498), .A2(n531), .ZN(n461) );
  XNOR2_X1 U329 ( .A(n391), .B(KEYINPUT47), .ZN(n392) );
  XNOR2_X1 U330 ( .A(n352), .B(KEYINPUT32), .ZN(n353) );
  XNOR2_X1 U331 ( .A(n393), .B(n392), .ZN(n400) );
  XNOR2_X1 U332 ( .A(G92GAT), .B(G36GAT), .ZN(n406) );
  XNOR2_X1 U333 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n419) );
  XNOR2_X1 U334 ( .A(n361), .B(n360), .ZN(n362) );
  INV_X1 U335 ( .A(n436), .ZN(n410) );
  XNOR2_X1 U336 ( .A(n420), .B(n419), .ZN(n572) );
  XNOR2_X1 U337 ( .A(n363), .B(n362), .ZN(n397) );
  XNOR2_X1 U338 ( .A(n491), .B(n490), .ZN(n517) );
  NOR2_X1 U339 ( .A1(n531), .A2(n458), .ZN(n568) );
  XNOR2_X1 U340 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n459) );
  XNOR2_X1 U341 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n292) );
  XNOR2_X1 U343 ( .A(G43GAT), .B(G99GAT), .ZN(n291) );
  XNOR2_X1 U344 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U345 ( .A(G120GAT), .B(G71GAT), .Z(n348) );
  XOR2_X1 U346 ( .A(n293), .B(n348), .Z(n295) );
  XNOR2_X1 U347 ( .A(G169GAT), .B(G15GAT), .ZN(n294) );
  XNOR2_X1 U348 ( .A(n295), .B(n294), .ZN(n308) );
  XOR2_X1 U349 ( .A(KEYINPUT84), .B(G176GAT), .Z(n297) );
  NAND2_X1 U350 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U351 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U352 ( .A(n298), .B(KEYINPUT85), .Z(n306) );
  XOR2_X1 U353 ( .A(KEYINPUT17), .B(G190GAT), .Z(n300) );
  XNOR2_X1 U354 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U356 ( .A(KEYINPUT19), .B(n301), .Z(n416) );
  XOR2_X1 U357 ( .A(KEYINPUT0), .B(G134GAT), .Z(n303) );
  XNOR2_X1 U358 ( .A(KEYINPUT83), .B(G127GAT), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U360 ( .A(G113GAT), .B(n304), .Z(n450) );
  XNOR2_X1 U361 ( .A(n416), .B(n450), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U363 ( .A(KEYINPUT76), .B(G162GAT), .Z(n429) );
  XOR2_X1 U364 ( .A(G85GAT), .B(KEYINPUT74), .Z(n310) );
  XNOR2_X1 U365 ( .A(G99GAT), .B(G92GAT), .ZN(n309) );
  XNOR2_X1 U366 ( .A(n310), .B(n309), .ZN(n355) );
  XOR2_X1 U367 ( .A(n429), .B(n355), .Z(n312) );
  NAND2_X1 U368 ( .A1(G232GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U370 ( .A(KEYINPUT11), .B(G106GAT), .Z(n314) );
  XNOR2_X1 U371 ( .A(G190GAT), .B(G134GAT), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U373 ( .A(n316), .B(n315), .Z(n326) );
  XOR2_X1 U374 ( .A(G43GAT), .B(G29GAT), .Z(n318) );
  XNOR2_X1 U375 ( .A(KEYINPUT8), .B(G50GAT), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U377 ( .A(n319), .B(KEYINPUT69), .Z(n321) );
  XNOR2_X1 U378 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n338) );
  XOR2_X1 U380 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n323) );
  XNOR2_X1 U381 ( .A(G218GAT), .B(KEYINPUT77), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U383 ( .A(n338), .B(n324), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n326), .B(n325), .ZN(n556) );
  XOR2_X1 U385 ( .A(G113GAT), .B(G197GAT), .Z(n328) );
  XOR2_X1 U386 ( .A(G169GAT), .B(G8GAT), .Z(n403) );
  XOR2_X1 U387 ( .A(G15GAT), .B(G1GAT), .Z(n377) );
  XNOR2_X1 U388 ( .A(n403), .B(n377), .ZN(n327) );
  XNOR2_X1 U389 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U390 ( .A(G141GAT), .B(G22GAT), .Z(n430) );
  XOR2_X1 U391 ( .A(n329), .B(n430), .Z(n334) );
  XOR2_X1 U392 ( .A(KEYINPUT67), .B(KEYINPUT65), .Z(n331) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U395 ( .A(KEYINPUT66), .B(n332), .ZN(n333) );
  XNOR2_X1 U396 ( .A(n334), .B(n333), .ZN(n340) );
  XOR2_X1 U397 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n336) );
  XNOR2_X1 U398 ( .A(KEYINPUT70), .B(KEYINPUT68), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U400 ( .A(n338), .B(n337), .Z(n339) );
  XNOR2_X1 U401 ( .A(n340), .B(n339), .ZN(n575) );
  INV_X1 U402 ( .A(G148GAT), .ZN(n341) );
  NAND2_X1 U403 ( .A1(n341), .A2(G78GAT), .ZN(n344) );
  INV_X1 U404 ( .A(G78GAT), .ZN(n342) );
  NAND2_X1 U405 ( .A1(n342), .A2(G148GAT), .ZN(n343) );
  NAND2_X1 U406 ( .A1(n344), .A2(n343), .ZN(n346) );
  XNOR2_X1 U407 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n431) );
  INV_X1 U409 ( .A(n431), .ZN(n347) );
  NAND2_X1 U410 ( .A1(n347), .A2(n348), .ZN(n351) );
  INV_X1 U411 ( .A(n348), .ZN(n349) );
  NAND2_X1 U412 ( .A1(n431), .A2(n349), .ZN(n350) );
  NAND2_X1 U413 ( .A1(n351), .A2(n350), .ZN(n354) );
  NAND2_X1 U414 ( .A1(G230GAT), .A2(G233GAT), .ZN(n352) );
  XOR2_X1 U415 ( .A(n355), .B(KEYINPUT72), .Z(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n363) );
  XOR2_X1 U417 ( .A(KEYINPUT75), .B(KEYINPUT31), .Z(n359) );
  XNOR2_X1 U418 ( .A(G204GAT), .B(KEYINPUT33), .ZN(n358) );
  XOR2_X1 U419 ( .A(n359), .B(n358), .Z(n361) );
  XOR2_X1 U420 ( .A(G176GAT), .B(G64GAT), .Z(n402) );
  XOR2_X1 U421 ( .A(KEYINPUT13), .B(G57GAT), .Z(n373) );
  XNOR2_X1 U422 ( .A(n402), .B(n373), .ZN(n360) );
  XNOR2_X1 U423 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n397), .B(n364), .ZN(n505) );
  NAND2_X1 U425 ( .A1(n575), .A2(n505), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n365), .B(KEYINPUT46), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n366), .B(KEYINPUT107), .ZN(n388) );
  XOR2_X1 U428 ( .A(G78GAT), .B(G155GAT), .Z(n368) );
  XNOR2_X1 U429 ( .A(G22GAT), .B(G211GAT), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U431 ( .A(G64GAT), .B(G71GAT), .Z(n370) );
  XNOR2_X1 U432 ( .A(G183GAT), .B(G127GAT), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U434 ( .A(n372), .B(n371), .Z(n379) );
  XOR2_X1 U435 ( .A(n373), .B(KEYINPUT15), .Z(n375) );
  NAND2_X1 U436 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U439 ( .A(n379), .B(n378), .ZN(n387) );
  XOR2_X1 U440 ( .A(KEYINPUT81), .B(KEYINPUT12), .Z(n381) );
  XNOR2_X1 U441 ( .A(G8GAT), .B(KEYINPUT78), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U443 ( .A(KEYINPUT82), .B(KEYINPUT14), .Z(n383) );
  XNOR2_X1 U444 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U446 ( .A(n385), .B(n384), .Z(n386) );
  XNOR2_X1 U447 ( .A(n387), .B(n386), .ZN(n583) );
  NOR2_X1 U448 ( .A1(n388), .A2(n583), .ZN(n389) );
  XOR2_X1 U449 ( .A(KEYINPUT108), .B(n389), .Z(n390) );
  NOR2_X1 U450 ( .A1(n556), .A2(n390), .ZN(n393) );
  INV_X1 U451 ( .A(KEYINPUT109), .ZN(n391) );
  INV_X1 U452 ( .A(n575), .ZN(n506) );
  XNOR2_X1 U453 ( .A(n506), .B(KEYINPUT71), .ZN(n561) );
  XOR2_X1 U454 ( .A(KEYINPUT45), .B(KEYINPUT110), .Z(n395) );
  XNOR2_X1 U455 ( .A(n556), .B(KEYINPUT36), .ZN(n585) );
  NAND2_X1 U456 ( .A1(n585), .A2(n583), .ZN(n394) );
  XOR2_X1 U457 ( .A(n395), .B(n394), .Z(n396) );
  NOR2_X1 U458 ( .A1(n561), .A2(n396), .ZN(n398) );
  NAND2_X1 U459 ( .A1(n398), .A2(n397), .ZN(n399) );
  NAND2_X1 U460 ( .A1(n400), .A2(n399), .ZN(n401) );
  XNOR2_X1 U461 ( .A(KEYINPUT48), .B(n401), .ZN(n530) );
  XOR2_X1 U462 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n405) );
  XNOR2_X1 U463 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n407), .B(n406), .ZN(n411) );
  XNOR2_X1 U466 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n289), .B(n408), .ZN(n409) );
  XOR2_X1 U468 ( .A(G197GAT), .B(n409), .Z(n436) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U470 ( .A(KEYINPUT94), .B(KEYINPUT78), .Z(n413) );
  NAND2_X1 U471 ( .A1(G226GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U473 ( .A(n415), .B(n414), .Z(n418) );
  XNOR2_X1 U474 ( .A(n416), .B(KEYINPUT91), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n520) );
  NAND2_X1 U476 ( .A1(n530), .A2(n520), .ZN(n420) );
  XOR2_X1 U477 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n422) );
  XNOR2_X1 U478 ( .A(G50GAT), .B(KEYINPUT88), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n428) );
  XOR2_X1 U480 ( .A(G155GAT), .B(KEYINPUT2), .Z(n424) );
  XNOR2_X1 U481 ( .A(KEYINPUT3), .B(KEYINPUT87), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n443) );
  XOR2_X1 U483 ( .A(n443), .B(KEYINPUT24), .Z(n426) );
  NAND2_X1 U484 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U485 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n468) );
  XOR2_X1 U491 ( .A(KEYINPUT1), .B(KEYINPUT89), .Z(n438) );
  XNOR2_X1 U492 ( .A(G1GAT), .B(G57GAT), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U494 ( .A(G148GAT), .B(G162GAT), .Z(n440) );
  XNOR2_X1 U495 ( .A(G141GAT), .B(G120GAT), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n454) );
  XOR2_X1 U498 ( .A(G85GAT), .B(n443), .Z(n445) );
  NAND2_X1 U499 ( .A1(G225GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U501 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n447) );
  XNOR2_X1 U502 ( .A(KEYINPUT90), .B(KEYINPUT5), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U504 ( .A(n449), .B(n448), .Z(n452) );
  XNOR2_X1 U505 ( .A(G29GAT), .B(n450), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n571) );
  INV_X1 U508 ( .A(n571), .ZN(n518) );
  NOR2_X1 U509 ( .A1(n468), .A2(n518), .ZN(n455) );
  AND2_X1 U510 ( .A1(n572), .A2(n455), .ZN(n457) );
  XNOR2_X1 U511 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n457), .B(n456), .ZN(n458) );
  NAND2_X1 U513 ( .A1(n568), .A2(n556), .ZN(n460) );
  XOR2_X1 U514 ( .A(KEYINPUT34), .B(KEYINPUT97), .Z(n478) );
  INV_X1 U515 ( .A(n520), .ZN(n498) );
  NOR2_X1 U516 ( .A1(n461), .A2(n468), .ZN(n462) );
  XOR2_X1 U517 ( .A(KEYINPUT25), .B(n462), .Z(n466) );
  XOR2_X1 U518 ( .A(n520), .B(KEYINPUT27), .Z(n528) );
  XOR2_X1 U519 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n464) );
  NAND2_X1 U520 ( .A1(n531), .A2(n468), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n464), .B(n463), .ZN(n574) );
  NOR2_X1 U522 ( .A1(n528), .A2(n574), .ZN(n465) );
  NAND2_X1 U523 ( .A1(n571), .A2(n467), .ZN(n472) );
  XNOR2_X1 U524 ( .A(KEYINPUT28), .B(n468), .ZN(n534) );
  NOR2_X1 U525 ( .A1(n534), .A2(n528), .ZN(n469) );
  NAND2_X1 U526 ( .A1(n469), .A2(n531), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n518), .A2(n470), .ZN(n471) );
  INV_X1 U528 ( .A(n583), .ZN(n473) );
  NOR2_X1 U529 ( .A1(n556), .A2(n473), .ZN(n474) );
  XOR2_X1 U530 ( .A(KEYINPUT16), .B(n474), .Z(n475) );
  NOR2_X1 U531 ( .A1(n487), .A2(n475), .ZN(n476) );
  XOR2_X1 U532 ( .A(KEYINPUT96), .B(n476), .Z(n507) );
  NAND2_X1 U533 ( .A1(n397), .A2(n561), .ZN(n492) );
  NOR2_X1 U534 ( .A1(n507), .A2(n492), .ZN(n485) );
  NAND2_X1 U535 ( .A1(n485), .A2(n518), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U537 ( .A(G1GAT), .B(n479), .ZN(G1324GAT) );
  NAND2_X1 U538 ( .A1(n485), .A2(n520), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n480), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n482) );
  INV_X1 U541 ( .A(n531), .ZN(n522) );
  NAND2_X1 U542 ( .A1(n485), .A2(n522), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n482), .B(n481), .ZN(n484) );
  XOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT98), .Z(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  NAND2_X1 U546 ( .A1(n485), .A2(n534), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n486), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U548 ( .A1(n487), .A2(n583), .ZN(n488) );
  XNOR2_X1 U549 ( .A(KEYINPUT100), .B(n488), .ZN(n489) );
  NAND2_X1 U550 ( .A1(n489), .A2(n585), .ZN(n491) );
  NOR2_X1 U551 ( .A1(n517), .A2(n492), .ZN(n493) );
  XOR2_X1 U552 ( .A(KEYINPUT38), .B(n493), .Z(n494) );
  XNOR2_X1 U553 ( .A(KEYINPUT102), .B(n494), .ZN(n502) );
  NOR2_X1 U554 ( .A1(n571), .A2(n502), .ZN(n496) );
  XNOR2_X1 U555 ( .A(KEYINPUT39), .B(KEYINPUT103), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U557 ( .A(G29GAT), .B(n497), .Z(G1328GAT) );
  NOR2_X1 U558 ( .A1(n498), .A2(n502), .ZN(n499) );
  XOR2_X1 U559 ( .A(KEYINPUT104), .B(n499), .Z(n500) );
  XNOR2_X1 U560 ( .A(G36GAT), .B(n500), .ZN(G1329GAT) );
  NOR2_X1 U561 ( .A1(n531), .A2(n502), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(n290), .ZN(G1330GAT) );
  INV_X1 U563 ( .A(n534), .ZN(n503) );
  NOR2_X1 U564 ( .A1(n503), .A2(n502), .ZN(n504) );
  XOR2_X1 U565 ( .A(G50GAT), .B(n504), .Z(G1331GAT) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n509) );
  NAND2_X1 U567 ( .A1(n506), .A2(n505), .ZN(n516) );
  NOR2_X1 U568 ( .A1(n507), .A2(n516), .ZN(n512) );
  NAND2_X1 U569 ( .A1(n512), .A2(n518), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n509), .B(n508), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n512), .A2(n520), .ZN(n510) );
  XNOR2_X1 U572 ( .A(n510), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U573 ( .A1(n522), .A2(n512), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U576 ( .A1(n512), .A2(n534), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U578 ( .A(G78GAT), .B(n515), .Z(G1335GAT) );
  NOR2_X1 U579 ( .A1(n517), .A2(n516), .ZN(n525) );
  NAND2_X1 U580 ( .A1(n525), .A2(n518), .ZN(n519) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n519), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n525), .A2(n520), .ZN(n521) );
  XNOR2_X1 U583 ( .A(n521), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U584 ( .A1(n522), .A2(n525), .ZN(n523) );
  XNOR2_X1 U585 ( .A(n523), .B(KEYINPUT106), .ZN(n524) );
  XNOR2_X1 U586 ( .A(G99GAT), .B(n524), .ZN(G1338GAT) );
  NAND2_X1 U587 ( .A1(n525), .A2(n534), .ZN(n526) );
  XNOR2_X1 U588 ( .A(n526), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n571), .A2(n528), .ZN(n529) );
  NAND2_X1 U591 ( .A1(n530), .A2(n529), .ZN(n548) );
  NOR2_X1 U592 ( .A1(n531), .A2(n548), .ZN(n532) );
  XNOR2_X1 U593 ( .A(n532), .B(KEYINPUT111), .ZN(n533) );
  NOR2_X1 U594 ( .A1(n534), .A2(n533), .ZN(n544) );
  NAND2_X1 U595 ( .A1(n561), .A2(n544), .ZN(n537) );
  XOR2_X1 U596 ( .A(G113GAT), .B(KEYINPUT112), .Z(n535) );
  XNOR2_X1 U597 ( .A(KEYINPUT113), .B(n535), .ZN(n536) );
  XNOR2_X1 U598 ( .A(n537), .B(n536), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U600 ( .A1(n544), .A2(n505), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n543) );
  XOR2_X1 U603 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n541) );
  NAND2_X1 U604 ( .A1(n544), .A2(n583), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U608 ( .A1(n544), .A2(n556), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(n547), .ZN(G1343GAT) );
  NOR2_X1 U611 ( .A1(n574), .A2(n548), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n557), .A2(n575), .ZN(n549) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n551) );
  NAND2_X1 U615 ( .A1(n557), .A2(n505), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n552), .ZN(G1345GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n554) );
  NAND2_X1 U619 ( .A1(n557), .A2(n583), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n555), .ZN(G1346GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n559) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n568), .A2(n561), .ZN(n562) );
  XNOR2_X1 U627 ( .A(G169GAT), .B(n562), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n564) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(n565), .Z(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n505), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  XOR2_X1 U634 ( .A(G183GAT), .B(KEYINPUT125), .Z(n570) );
  NAND2_X1 U635 ( .A1(n568), .A2(n583), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1350GAT) );
  XNOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n579) );
  XOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT126), .Z(n577) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n586) );
  NAND2_X1 U641 ( .A1(n586), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  INV_X1 U645 ( .A(n397), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n586), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n586), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n588) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

