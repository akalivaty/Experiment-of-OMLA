//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G128), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n190), .B(new_n192), .C1(G119), .C2(new_n191), .ZN(new_n193));
  XNOR2_X1  g007(.A(G119), .B(G128), .ZN(new_n194));
  XOR2_X1   g008(.A(KEYINPUT24), .B(G110), .Z(new_n195));
  AOI22_X1  g009(.A1(new_n193), .A2(G110), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G125), .B(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT16), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G125), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n198), .A2(G146), .A3(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(G146), .B1(new_n198), .B2(new_n201), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n196), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  OAI22_X1  g018(.A1(new_n193), .A2(G110), .B1(new_n194), .B2(new_n195), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n198), .A2(G146), .A3(new_n201), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n197), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G953), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(G221), .A3(G234), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n212), .B(KEYINPUT73), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT22), .B(G137), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n213), .B(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n204), .A3(new_n209), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n187), .B1(new_n219), .B2(G902), .ZN(new_n220));
  INV_X1    g034(.A(G902), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n217), .A2(KEYINPUT25), .A3(new_n221), .A4(new_n218), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n220), .A2(KEYINPUT74), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G217), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(G234), .B2(new_n221), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(new_n220), .B2(KEYINPUT74), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(G902), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  OAI22_X1  g042(.A1(new_n223), .A2(new_n226), .B1(new_n219), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n231));
  XNOR2_X1  g045(.A(G134), .B(G137), .ZN(new_n232));
  INV_X1    g046(.A(G131), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n235));
  INV_X1    g049(.A(G134), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G137), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT11), .A3(G134), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(G137), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n237), .A2(new_n239), .A3(new_n233), .A4(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n236), .A2(G137), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n238), .A2(G134), .ZN(new_n243));
  OAI211_X1 g057(.A(KEYINPUT66), .B(G131), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n234), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT1), .B1(new_n247), .B2(G146), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G128), .ZN(new_n249));
  XNOR2_X1  g063(.A(G143), .B(G146), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n207), .A2(G143), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(G146), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n252), .B(new_n253), .C1(KEYINPUT1), .C2(new_n191), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n246), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(new_n253), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(G128), .A3(new_n248), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT69), .A3(new_n254), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n245), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT65), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT0), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(new_n191), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n257), .A2(new_n261), .A3(new_n262), .A4(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n250), .A2(KEYINPUT0), .A3(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n237), .A2(new_n240), .A3(new_n239), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G131), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n268), .B1(new_n241), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n230), .B1(new_n260), .B2(new_n271), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n234), .A2(new_n241), .A3(new_n244), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n258), .A2(KEYINPUT69), .A3(new_n254), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT69), .B1(new_n258), .B2(new_n254), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n270), .A2(new_n241), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n266), .A3(new_n267), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n276), .A2(KEYINPUT70), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(KEYINPUT2), .A2(G113), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT67), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OR2_X1    g098(.A1(KEYINPUT2), .A2(G113), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n189), .A2(G116), .ZN(new_n287));
  INV_X1    g101(.A(G116), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G119), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G116), .B(G119), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT68), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n286), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n284), .A2(new_n285), .A3(new_n293), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n272), .A2(new_n279), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT28), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n260), .A2(new_n271), .A3(new_n297), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n298), .B1(new_n276), .B2(new_n278), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT72), .B1(new_n305), .B2(new_n301), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n276), .A2(new_n278), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n297), .B1(new_n307), .B2(new_n230), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT28), .B1(new_n308), .B2(new_n279), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n302), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G237), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(new_n211), .A3(G210), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT27), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT26), .B(G101), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n315), .A2(KEYINPUT29), .ZN(new_n316));
  AOI21_X1  g130(.A(G902), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n276), .A2(KEYINPUT30), .A3(new_n278), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n319));
  NAND2_X1  g133(.A1(new_n258), .A2(new_n254), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n245), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n319), .B1(new_n271), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n318), .A2(new_n322), .A3(new_n297), .ZN(new_n323));
  INV_X1    g137(.A(new_n303), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n315), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT29), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n299), .A2(new_n301), .ZN(new_n328));
  INV_X1    g142(.A(new_n321), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n298), .B1(new_n329), .B2(new_n278), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT28), .B1(new_n303), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n331), .A3(new_n315), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT71), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n327), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n327), .A2(new_n332), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT71), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n317), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G472), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n323), .A2(new_n324), .A3(new_n315), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT31), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT31), .A4(new_n315), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n328), .A2(new_n331), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n326), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT32), .ZN(new_n347));
  INV_X1    g161(.A(G472), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .A4(new_n221), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n341), .A2(new_n342), .B1(new_n344), .B2(new_n326), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n221), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT32), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n229), .B1(new_n338), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT9), .B(G234), .ZN(new_n355));
  OAI21_X1  g169(.A(G221), .B1(new_n355), .B2(G902), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G469), .ZN(new_n358));
  OR2_X1    g172(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n359));
  INV_X1    g173(.A(G107), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G104), .ZN(new_n361));
  AND2_X1   g175(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT76), .B(G101), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n360), .A2(G104), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(G107), .ZN(new_n368));
  NOR2_X1   g182(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n363), .A2(new_n364), .A3(new_n366), .A4(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT77), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n365), .B1(new_n369), .B2(new_n368), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n374), .A2(KEYINPUT77), .A3(new_n364), .A4(new_n363), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n320), .ZN(new_n377));
  INV_X1    g191(.A(G101), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n378), .B1(new_n366), .B2(new_n361), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n376), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT10), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n378), .B1(new_n374), .B2(new_n363), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n376), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n268), .B1(new_n385), .B2(new_n384), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n277), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n382), .B1(new_n256), .B2(new_n259), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n379), .B1(new_n373), .B2(new_n375), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n383), .A2(new_n389), .A3(new_n390), .A4(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(G110), .B(G140), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n211), .A2(G227), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n395), .B(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n377), .B1(new_n376), .B2(new_n380), .ZN(new_n400));
  AOI211_X1 g214(.A(new_n379), .B(new_n320), .C1(new_n373), .C2(new_n375), .ZN(new_n401));
  OAI211_X1 g215(.A(KEYINPUT12), .B(new_n277), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n277), .B1(new_n400), .B2(new_n401), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT12), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n399), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n387), .A2(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n383), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n277), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n398), .B1(new_n409), .B2(new_n394), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n358), .B(new_n221), .C1(new_n406), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT78), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n376), .A2(new_n380), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n320), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n381), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT12), .B1(new_n415), .B2(new_n277), .ZN(new_n416));
  INV_X1    g230(.A(new_n402), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n394), .B(new_n398), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n394), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n390), .B1(new_n407), .B2(new_n383), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n397), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(G902), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT78), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n358), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n412), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n405), .A2(new_n402), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n398), .B1(new_n426), .B2(new_n394), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n399), .A2(new_n420), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G469), .B1(new_n429), .B2(G902), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n357), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(G214), .B1(G237), .B2(G902), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G110), .B(G122), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n384), .A2(new_n385), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n297), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(new_n376), .B2(new_n386), .ZN(new_n438));
  INV_X1    g252(.A(new_n296), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(new_n287), .ZN(new_n441));
  INV_X1    g255(.A(G113), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n290), .A2(new_n291), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n293), .A2(KEYINPUT68), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n440), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n439), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n447), .A2(new_n392), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n435), .B1(new_n438), .B2(new_n448), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n297), .A2(new_n436), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n450), .A2(new_n387), .B1(new_n392), .B2(new_n447), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n434), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n452), .A3(KEYINPUT6), .ZN(new_n453));
  OR3_X1    g267(.A1(new_n451), .A2(KEYINPUT6), .A3(new_n434), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n268), .A2(G125), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n455), .B1(G125), .B2(new_n377), .ZN(new_n456));
  INV_X1    g270(.A(G224), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(G953), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n456), .B(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n453), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT7), .B1(new_n457), .B2(G953), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n461), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n455), .B(new_n463), .C1(G125), .C2(new_n377), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n465), .B1(new_n434), .B2(new_n451), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n442), .B(new_n441), .C1(KEYINPUT5), .C2(new_n293), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n392), .B1(new_n467), .B2(new_n439), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n413), .A2(new_n447), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n434), .B(KEYINPUT8), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(G902), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n460), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G210), .B1(G237), .B2(G902), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n460), .A2(new_n474), .A3(new_n472), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n433), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n202), .A2(new_n203), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n311), .A2(new_n211), .A3(G214), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n247), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n311), .A2(new_n211), .A3(G143), .A4(G214), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(KEYINPUT17), .A3(G131), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(G131), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n479), .B(new_n484), .C1(new_n485), .C2(KEYINPUT17), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT80), .B1(new_n197), .B2(new_n207), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(new_n207), .B2(new_n197), .ZN(new_n488));
  INV_X1    g302(.A(new_n197), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(KEYINPUT80), .A3(G146), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n483), .A2(KEYINPUT18), .A3(G131), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n483), .ZN(new_n493));
  NAND2_X1  g307(.A1(KEYINPUT18), .A2(G131), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT81), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n493), .A2(KEYINPUT82), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n481), .A3(new_n482), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT82), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n492), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n486), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G113), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(new_n367), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(KEYINPUT84), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n221), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n503), .A2(new_n506), .ZN(new_n509));
  OAI21_X1  g323(.A(G475), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT83), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n197), .B(KEYINPUT19), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n202), .B1(new_n207), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n501), .A2(new_n492), .B1(new_n513), .B2(new_n485), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n511), .B1(new_n514), .B2(new_n505), .ZN(new_n515));
  INV_X1    g329(.A(new_n505), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n492), .A2(new_n501), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n512), .A2(new_n207), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n485), .A2(new_n206), .A3(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(KEYINPUT83), .B(new_n516), .C1(new_n517), .C2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n486), .A2(new_n502), .A3(new_n505), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n515), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT20), .ZN(new_n523));
  NOR2_X1   g337(.A1(G475), .A2(G902), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n523), .B1(new_n522), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n510), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT85), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n191), .A2(G143), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n528), .B1(new_n529), .B2(KEYINPUT13), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n247), .A2(G128), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT13), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(KEYINPUT85), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n191), .A2(G143), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n531), .B2(new_n532), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT86), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n539), .A3(G134), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n536), .B1(new_n530), .B2(new_n533), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT86), .B1(new_n541), .B2(new_n236), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n531), .A2(new_n535), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(KEYINPUT87), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT87), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n531), .B2(new_n535), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n236), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(G116), .B(G122), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(new_n360), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n545), .ZN(new_n553));
  INV_X1    g367(.A(new_n547), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(G134), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n548), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n288), .A2(G122), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n360), .B1(new_n557), .B2(KEYINPUT14), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(new_n549), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n355), .A2(new_n224), .A3(G953), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n552), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n552), .B2(new_n560), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n221), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G478), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT88), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(KEYINPUT15), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(KEYINPUT15), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n552), .A2(new_n560), .ZN(new_n572));
  INV_X1    g386(.A(new_n561), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n552), .A2(new_n560), .A3(new_n561), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n570), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n221), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n571), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(KEYINPUT89), .A2(G952), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(KEYINPUT89), .A2(G952), .ZN(new_n582));
  AOI21_X1  g396(.A(G953), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(G234), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(new_n311), .ZN(new_n585));
  AOI211_X1 g399(.A(new_n221), .B(new_n211), .C1(G234), .C2(G237), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT21), .B(G898), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n527), .A2(new_n579), .A3(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n354), .A2(new_n431), .A3(new_n478), .A4(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n591), .B(new_n364), .Z(G3));
  OAI21_X1  g406(.A(G472), .B1(new_n350), .B2(G902), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n350), .B2(new_n351), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(new_n229), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n431), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT33), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n573), .B2(KEYINPUT90), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n576), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n574), .A2(new_n575), .A3(new_n598), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n565), .A2(G902), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n564), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT91), .B(G478), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n527), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n589), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n460), .A2(new_n474), .A3(new_n472), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n474), .B1(new_n460), .B2(new_n472), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n432), .B(new_n608), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n596), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT34), .B(G104), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  INV_X1    g428(.A(KEYINPUT92), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n579), .B(new_n510), .C1(new_n525), .C2(new_n526), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n615), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n616), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n478), .A2(new_n618), .A3(KEYINPUT92), .A4(new_n608), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(new_n431), .A3(new_n595), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT35), .B(G107), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  INV_X1    g437(.A(KEYINPUT93), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n210), .B(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n216), .A2(KEYINPUT36), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n227), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n629), .B1(new_n223), .B2(new_n226), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT94), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT94), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n629), .B(new_n632), .C1(new_n223), .C2(new_n226), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n594), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n431), .A2(new_n635), .A3(new_n478), .A4(new_n590), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT37), .B(G110), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT96), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(KEYINPUT95), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n636), .B(new_n639), .ZN(G12));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n641));
  INV_X1    g455(.A(new_n585), .ZN(new_n642));
  INV_X1    g456(.A(G900), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n642), .B1(new_n643), .B2(new_n586), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n616), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n431), .A2(new_n478), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n634), .B1(new_n338), .B2(new_n353), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n641), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n418), .A2(new_n421), .ZN(new_n650));
  AND4_X1   g464(.A1(new_n423), .A2(new_n650), .A3(new_n358), .A4(new_n221), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n423), .B1(new_n422), .B2(new_n358), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n430), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n653), .A2(new_n356), .A3(new_n478), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n654), .A2(KEYINPUT97), .A3(new_n647), .A4(new_n645), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  NAND2_X1  g471(.A1(new_n476), .A2(new_n477), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n527), .A2(new_n579), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n432), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n644), .B(KEYINPUT39), .Z(new_n663));
  NAND2_X1  g477(.A1(new_n431), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n662), .B1(KEYINPUT40), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n305), .A2(new_n315), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT99), .ZN(new_n667));
  INV_X1    g481(.A(new_n339), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n221), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(G472), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n353), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n353), .A2(new_n670), .A3(KEYINPUT100), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n630), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n665), .B(new_n675), .C1(KEYINPUT40), .C2(new_n664), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  NOR2_X1   g491(.A1(new_n607), .A2(new_n644), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n654), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n648), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT101), .B(G146), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G48));
  OR2_X1    g496(.A1(new_n422), .A2(new_n358), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n425), .A2(new_n356), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n607), .ZN(new_n685));
  INV_X1    g499(.A(new_n611), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n684), .A2(new_n354), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT41), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G113), .ZN(G15));
  NAND3_X1  g503(.A1(new_n620), .A2(new_n354), .A3(new_n684), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G116), .ZN(G18));
  NAND4_X1  g505(.A1(new_n684), .A2(new_n647), .A3(new_n478), .A4(new_n590), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G119), .ZN(G21));
  AOI21_X1  g507(.A(new_n348), .B1(new_n346), .B2(new_n221), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n326), .B(new_n302), .C1(new_n306), .C2(new_n309), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n351), .B1(new_n695), .B2(new_n343), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n694), .A2(new_n229), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n684), .A2(new_n686), .A3(new_n661), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G122), .ZN(G24));
  NAND2_X1  g513(.A1(new_n684), .A2(new_n478), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n694), .A2(new_n696), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n678), .A2(new_n630), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G125), .ZN(G27));
  AND3_X1   g520(.A1(new_n425), .A2(KEYINPUT102), .A3(new_n430), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT102), .B1(new_n425), .B2(new_n430), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n658), .A2(new_n357), .A3(new_n433), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(new_n354), .A3(new_n678), .A4(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT104), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n653), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n425), .A2(KEYINPUT102), .A3(new_n430), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n715), .A2(new_n354), .A3(new_n710), .A4(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n678), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n720), .A3(KEYINPUT42), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n712), .B1(new_n717), .B2(new_n718), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT103), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n724), .B(new_n712), .C1(new_n717), .C2(new_n718), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n713), .A2(new_n721), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n233), .ZN(G33));
  NAND4_X1  g541(.A1(new_n709), .A2(new_n354), .A3(new_n645), .A4(new_n710), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G134), .ZN(G36));
  NAND2_X1  g543(.A1(new_n429), .A2(KEYINPUT45), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n427), .B2(new_n428), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(G469), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(G469), .A2(G902), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT46), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n412), .B2(new_n424), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n733), .A2(KEYINPUT46), .A3(new_n734), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n357), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n663), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT105), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n658), .A2(new_n433), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n604), .A2(new_n605), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n600), .A2(new_n601), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n743), .B1(new_n744), .B2(new_n602), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n527), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT43), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n594), .A3(new_n630), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n742), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n750), .B1(new_n749), .B2(new_n748), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n740), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G137), .ZN(G39));
  NAND2_X1  g567(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n738), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g569(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n756));
  OAI21_X1  g570(.A(new_n755), .B1(new_n738), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n338), .A2(new_n353), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n678), .A2(new_n741), .A3(new_n229), .ZN(new_n759));
  OR3_X1    g573(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G140), .ZN(G42));
  NOR2_X1   g575(.A1(G952), .A2(G953), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT116), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n425), .A2(new_n683), .ZN(new_n764));
  NOR4_X1   g578(.A1(new_n742), .A2(new_n764), .A3(new_n357), .A4(new_n585), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n747), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n702), .A2(new_n630), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n747), .A2(new_n642), .A3(new_n697), .ZN(new_n769));
  INV_X1    g583(.A(new_n660), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n433), .A3(new_n770), .A4(new_n684), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT113), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n673), .A2(new_n674), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n229), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(new_n765), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n527), .A2(new_n606), .ZN(new_n778));
  AOI211_X1 g592(.A(new_n768), .B(new_n774), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT51), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n764), .B(KEYINPUT107), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n757), .B1(new_n356), .B2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n769), .A2(new_n741), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n785), .B1(new_n782), .B2(new_n783), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n780), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n782), .A2(new_n741), .A3(new_n769), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT51), .B1(new_n779), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n765), .A2(new_n354), .A3(new_n747), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT48), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n769), .A2(new_n478), .A3(new_n684), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n583), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n795), .B1(new_n792), .B2(new_n793), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n777), .A2(new_n685), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n791), .A2(new_n794), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  OR3_X1    g612(.A1(new_n787), .A2(new_n789), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n800));
  OAI22_X1  g614(.A1(new_n679), .A2(new_n648), .B1(new_n700), .B2(new_n703), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n649), .B2(new_n655), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n661), .A2(new_n478), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n357), .A3(new_n644), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n675), .A2(new_n709), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT52), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n801), .ZN(new_n807));
  AND4_X1   g621(.A1(KEYINPUT52), .A2(new_n807), .A3(new_n656), .A4(new_n805), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n690), .A2(new_n692), .A3(new_n687), .A4(new_n698), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n654), .B(new_n590), .C1(new_n354), .C2(new_n635), .ZN(new_n811));
  INV_X1    g625(.A(new_n526), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT108), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n815), .A3(new_n579), .A4(new_n510), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n616), .A2(KEYINPUT108), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n817), .A3(new_n607), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n431), .A2(new_n595), .A3(new_n686), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n811), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT109), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT109), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n811), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n810), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n709), .A2(new_n704), .A3(new_n710), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n634), .A2(new_n579), .A3(new_n527), .A4(new_n644), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n758), .A3(new_n653), .A4(new_n710), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n728), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n713), .A2(new_n721), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n723), .A2(new_n725), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n809), .A2(KEYINPUT53), .A3(new_n824), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n806), .A2(new_n808), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n724), .B1(new_n711), .B2(new_n712), .ZN(new_n834));
  INV_X1    g648(.A(new_n725), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n720), .B1(new_n719), .B2(KEYINPUT42), .ZN(new_n836));
  NOR4_X1   g650(.A1(new_n717), .A2(KEYINPUT104), .A3(new_n712), .A4(new_n718), .ZN(new_n837));
  OAI22_X1  g651(.A1(new_n834), .A2(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n828), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n824), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT110), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT110), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n831), .A2(new_n842), .A3(new_n824), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n833), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  XOR2_X1   g658(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n800), .B(new_n832), .C1(new_n844), .C2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT112), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n842), .B1(new_n831), .B2(new_n824), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n687), .A2(new_n690), .A3(new_n692), .A4(new_n698), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n822), .B1(new_n811), .B2(new_n819), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n822), .A2(new_n591), .A3(new_n636), .A4(new_n819), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR4_X1   g668(.A1(new_n726), .A2(new_n854), .A3(KEYINPUT110), .A4(new_n828), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n809), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT53), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n844), .A2(new_n845), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT54), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n845), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n860), .A2(KEYINPUT112), .A3(new_n800), .A4(new_n832), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n849), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n763), .B1(new_n799), .B2(new_n862), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n781), .A2(KEYINPUT49), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n781), .A2(KEYINPUT49), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n356), .A2(new_n770), .A3(new_n432), .A4(new_n746), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n864), .A2(new_n776), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n863), .A2(new_n867), .ZN(G75));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n833), .A2(new_n869), .A3(new_n840), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n856), .B2(new_n845), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n871), .A2(new_n221), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(G210), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n453), .A2(new_n454), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(new_n459), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT55), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n873), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n877), .B1(new_n873), .B2(new_n874), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n211), .A2(G952), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G51));
  XOR2_X1   g695(.A(new_n734), .B(KEYINPUT57), .Z(new_n882));
  NOR2_X1   g696(.A1(new_n871), .A2(new_n800), .ZN(new_n883));
  INV_X1    g697(.A(new_n847), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT117), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n887), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n650), .A3(new_n888), .ZN(new_n889));
  OR3_X1    g703(.A1(new_n871), .A2(new_n221), .A3(new_n733), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n880), .B1(new_n889), .B2(new_n890), .ZN(G54));
  NAND3_X1  g705(.A1(new_n872), .A2(KEYINPUT58), .A3(G475), .ZN(new_n892));
  INV_X1    g706(.A(new_n522), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(new_n880), .ZN(G60));
  NAND2_X1  g710(.A1(new_n860), .A2(new_n832), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n847), .ZN(new_n899));
  XNOR2_X1  g713(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n900));
  NAND2_X1  g714(.A1(G478), .A2(G902), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n900), .B(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n744), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n880), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n744), .B1(new_n862), .B2(new_n902), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n904), .B1(new_n905), .B2(KEYINPUT119), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n907));
  AOI211_X1 g721(.A(new_n907), .B(new_n744), .C1(new_n862), .C2(new_n902), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n906), .A2(new_n908), .ZN(G63));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n910));
  XNOR2_X1  g724(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n224), .A2(new_n221), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n219), .B1(new_n871), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n880), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n627), .A2(new_n628), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n897), .A2(new_n918), .A3(new_n913), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT121), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n919), .A2(KEYINPUT121), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n910), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n917), .A2(KEYINPUT122), .A3(KEYINPUT61), .A4(new_n919), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n919), .A2(new_n915), .A3(KEYINPUT61), .A4(new_n916), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n923), .A2(new_n928), .ZN(G66));
  OAI21_X1  g743(.A(G953), .B1(new_n587), .B2(new_n457), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n824), .B2(G953), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n875), .B1(G898), .B2(new_n211), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(G69));
  AOI21_X1  g747(.A(new_n211), .B1(G227), .B2(G900), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n802), .A2(new_n676), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT62), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT123), .Z(new_n937));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n935), .A2(KEYINPUT62), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n354), .A2(new_n741), .A3(new_n818), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n940), .A2(new_n664), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n752), .A2(new_n939), .A3(new_n760), .A4(new_n941), .ZN(new_n942));
  OR3_X1    g756(.A1(new_n937), .A2(new_n938), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n938), .B1(new_n937), .B2(new_n942), .ZN(new_n944));
  AOI21_X1  g758(.A(G953), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n318), .A2(new_n322), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(new_n512), .Z(new_n947));
  NOR2_X1   g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n760), .A2(new_n728), .A3(new_n802), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n354), .A2(new_n478), .A3(new_n661), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n740), .B1(new_n751), .B2(new_n950), .ZN(new_n951));
  NOR4_X1   g765(.A1(new_n949), .A2(new_n951), .A3(G953), .A4(new_n726), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n947), .B1(new_n643), .B2(new_n211), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n934), .B1(new_n948), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n934), .ZN(new_n956));
  OAI221_X1 g770(.A(new_n956), .B1(new_n952), .B2(new_n953), .C1(new_n945), .C2(new_n947), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(G72));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n959));
  OR4_X1    g773(.A1(new_n726), .A2(new_n949), .A3(new_n854), .A4(new_n951), .ZN(new_n960));
  XOR2_X1   g774(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n961));
  NOR2_X1   g775(.A1(new_n348), .A2(new_n221), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n325), .B(KEYINPUT126), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n326), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n959), .B(new_n916), .C1(new_n964), .C2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n960), .B2(new_n963), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT127), .B1(new_n968), .B2(new_n880), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n943), .A2(new_n824), .A3(new_n944), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n963), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n965), .A2(new_n326), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n325), .A2(new_n326), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n339), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n857), .A2(new_n858), .A3(new_n963), .A4(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n970), .A2(new_n974), .A3(new_n977), .ZN(G57));
endmodule


