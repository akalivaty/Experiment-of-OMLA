//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1196, new_n1197, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1265, new_n1266, new_n1267, new_n1268;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G87), .A2(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n202), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n214), .C1(G116), .C2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G1), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n222), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NOR2_X1   g0029(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G20), .ZN(new_n233));
  OAI21_X1  g0033(.A(G50), .B1(G58), .B2(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT64), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n225), .B(new_n230), .C1(new_n233), .C2(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT66), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XOR2_X1   g0050(.A(G50), .B(G58), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  OR2_X1    g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G232), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n256), .B(new_n258), .C1(new_n213), .C2(new_n257), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n259), .B(new_n262), .C1(G107), .C2(new_n256), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n219), .B1(G41), .B2(G45), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n261), .A2(new_n264), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n263), .B(new_n267), .C1(new_n208), .C2(new_n268), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n269), .A2(G179), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n219), .A2(G13), .A3(G20), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G77), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G20), .A2(G77), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT15), .B(G87), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n220), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT8), .B(G58), .ZN(new_n278));
  OAI221_X1 g0078(.A(new_n273), .B1(new_n274), .B2(new_n275), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n231), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n272), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n281), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n219), .A2(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G77), .A3(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G169), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n269), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n270), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n256), .B1(G232), .B2(new_n257), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G226), .A2(G1698), .ZN(new_n293));
  INV_X1    g0093(.A(G33), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n292), .A2(new_n293), .B1(new_n294), .B2(new_n216), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n266), .B1(new_n295), .B2(new_n262), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT13), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n261), .A2(G238), .A3(new_n264), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n297), .B1(new_n296), .B2(new_n298), .ZN(new_n300));
  OAI21_X1  g0100(.A(G169), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT14), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n299), .A2(new_n300), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G179), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT14), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n305), .B(G169), .C1(new_n299), .C2(new_n300), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n302), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n283), .A2(new_n284), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT12), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n219), .A2(new_n212), .A3(G13), .A4(G20), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n308), .A2(new_n212), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n276), .A2(G50), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n312), .B1(new_n220), .B2(G68), .C1(new_n207), .C2(new_n275), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n281), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  XOR2_X1   g0115(.A(KEYINPUT72), .B(KEYINPUT11), .Z(new_n316));
  AOI21_X1  g0116(.A(new_n311), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n310), .A2(new_n309), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n317), .B(new_n318), .C1(new_n315), .C2(new_n316), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n319), .B(KEYINPUT73), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n307), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT73), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n319), .B(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n303), .A2(G190), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n323), .B(new_n324), .C1(new_n325), .C2(new_n303), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT74), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n291), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XOR2_X1   g0129(.A(KEYINPUT69), .B(G200), .Z(new_n330));
  NAND2_X1  g0130(.A1(new_n269), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n286), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT70), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G190), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n269), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT16), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n254), .A2(new_n220), .A3(new_n255), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT7), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n220), .A4(new_n255), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n212), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G58), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n212), .ZN(new_n346));
  OAI21_X1  g0146(.A(G20), .B1(new_n346), .B2(new_n201), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n276), .A2(G159), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n339), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(KEYINPUT3), .A2(G33), .ZN(new_n351));
  NOR2_X1   g0151(.A1(KEYINPUT3), .A2(G33), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT7), .B1(new_n353), .B2(new_n220), .ZN(new_n354));
  NOR4_X1   g0154(.A1(new_n351), .A2(new_n352), .A3(new_n341), .A4(G20), .ZN(new_n355));
  OAI21_X1  g0155(.A(G68), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n349), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(KEYINPUT16), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n350), .A2(new_n358), .A3(new_n281), .ZN(new_n359));
  INV_X1    g0159(.A(G223), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n257), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n211), .A2(G1698), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n361), .B(new_n362), .C1(new_n351), .C2(new_n352), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G87), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n262), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n261), .A2(G232), .A3(new_n264), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n366), .A2(new_n335), .A3(new_n368), .A4(new_n267), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n261), .B1(new_n363), .B2(new_n364), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n370), .A2(new_n367), .A3(new_n266), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n369), .B1(new_n371), .B2(G200), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT75), .ZN(new_n373));
  OR2_X1    g0173(.A1(KEYINPUT8), .A2(G58), .ZN(new_n374));
  NAND2_X1  g0174(.A1(KEYINPUT8), .A2(G58), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(KEYINPUT67), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n271), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT67), .B1(new_n374), .B2(new_n375), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT67), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n278), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(new_n376), .B1(new_n283), .B2(new_n284), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n373), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n308), .B1(new_n377), .B2(new_n379), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n271), .A3(new_n376), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(KEYINPUT75), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n389));
  AND4_X1   g0189(.A1(new_n359), .A2(new_n372), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n359), .A2(new_n372), .A3(new_n388), .ZN(new_n391));
  OR2_X1    g0191(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n359), .A2(new_n388), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n266), .B1(new_n365), .B2(new_n262), .ZN(new_n396));
  AOI21_X1  g0196(.A(G169), .B1(new_n396), .B2(new_n368), .ZN(new_n397));
  NOR4_X1   g0197(.A1(new_n370), .A2(G179), .A3(new_n367), .A4(new_n266), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT18), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n395), .A2(KEYINPUT18), .A3(new_n399), .ZN(new_n401));
  OAI221_X1 g0201(.A(new_n394), .B1(new_n400), .B2(new_n401), .C1(new_n327), .C2(new_n328), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n271), .A2(G50), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n284), .A2(KEYINPUT68), .A3(G50), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT68), .B1(new_n284), .B2(G50), .ZN(new_n406));
  NOR4_X1   g0206(.A1(new_n405), .A2(new_n406), .A3(new_n378), .A4(new_n281), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n203), .A2(G20), .ZN(new_n408));
  INV_X1    g0208(.A(G150), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n377), .A2(new_n379), .ZN(new_n410));
  OAI221_X1 g0210(.A(new_n408), .B1(new_n409), .B2(new_n277), .C1(new_n410), .C2(new_n275), .ZN(new_n411));
  AOI211_X1 g0211(.A(new_n403), .B(new_n407), .C1(new_n411), .C2(new_n281), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n412), .A2(KEYINPUT9), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n257), .A2(G222), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n256), .B(new_n414), .C1(new_n360), .C2(new_n257), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n415), .B(new_n262), .C1(G77), .C2(new_n256), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n416), .B(new_n267), .C1(new_n211), .C2(new_n268), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n417), .A2(new_n335), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n412), .A2(KEYINPUT9), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT71), .B1(new_n417), .B2(new_n330), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n413), .A2(new_n418), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT10), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n419), .A2(new_n420), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT10), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n423), .A2(new_n413), .A3(new_n424), .A4(new_n418), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n412), .B1(new_n288), .B2(new_n417), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(G179), .B2(new_n417), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n338), .A2(new_n402), .A3(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT5), .B(G41), .ZN(new_n431));
  INV_X1    g0231(.A(G45), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(G1), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n431), .A2(new_n433), .B1(new_n232), .B2(new_n260), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n434), .A2(G264), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n217), .A2(G1698), .ZN(new_n436));
  OAI221_X1 g0236(.A(new_n436), .B1(G250), .B2(G1698), .C1(new_n351), .C2(new_n352), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G294), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n261), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n219), .A2(G45), .ZN(new_n440));
  NOR2_X1   g0240(.A1(KEYINPUT5), .A2(G41), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G274), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n435), .A2(new_n439), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(G169), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G116), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(G20), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT81), .B1(new_n220), .B2(G107), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT23), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT23), .ZN(new_n453));
  OAI211_X1 g0253(.A(KEYINPUT81), .B(new_n453), .C1(new_n220), .C2(G107), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n450), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n220), .B(G87), .C1(new_n351), .C2(new_n352), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT80), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT22), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n457), .A2(new_n458), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n456), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n256), .A2(new_n220), .A3(G87), .A4(new_n460), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n455), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT24), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT24), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n455), .A2(new_n462), .A3(new_n466), .A4(new_n463), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n219), .A2(G33), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n283), .A2(new_n271), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n468), .A2(new_n281), .B1(G107), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G107), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n378), .B(new_n473), .C1(KEYINPUT82), .C2(KEYINPUT25), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n474), .B(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n448), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n437), .A2(new_n438), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n262), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n434), .A2(G264), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n445), .A3(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G179), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G303), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n261), .B1(new_n353), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n257), .A2(G257), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G264), .A2(G1698), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n488), .C1(new_n351), .C2(new_n352), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n486), .A2(new_n489), .B1(G274), .B2(new_n444), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT78), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n434), .B2(G270), .ZN(new_n492));
  INV_X1    g0292(.A(new_n443), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n433), .B1(new_n493), .B2(new_n441), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n494), .A2(new_n491), .A3(G270), .A4(new_n261), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n490), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G116), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n378), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n283), .A2(G116), .A3(new_n271), .A4(new_n469), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n280), .A2(new_n231), .B1(G20), .B2(new_n498), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G283), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n502), .B(new_n220), .C1(G33), .C2(new_n216), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n501), .A2(KEYINPUT20), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT20), .B1(new_n501), .B2(new_n503), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n499), .B(new_n500), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n497), .A2(G169), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT21), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n494), .A2(G270), .A3(new_n261), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT78), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n495), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n288), .B1(new_n512), .B2(new_n490), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(KEYINPUT21), .A3(new_n506), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n490), .B(G190), .C1(new_n492), .C2(new_n496), .ZN(new_n515));
  INV_X1    g0315(.A(new_n506), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n254), .A2(new_n485), .A3(new_n255), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n489), .A2(new_n262), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n445), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n511), .B2(new_n495), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n515), .B(new_n516), .C1(new_n520), .C2(new_n325), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(G179), .A3(new_n506), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n509), .A2(new_n514), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT79), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n523), .A2(new_n524), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n484), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n271), .A2(G97), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n470), .A2(new_n216), .ZN(new_n529));
  OAI21_X1  g0329(.A(G107), .B1(new_n354), .B2(new_n355), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT6), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n216), .A2(new_n473), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n473), .A2(KEYINPUT6), .A3(G97), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G20), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n276), .A2(G77), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n530), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI211_X1 g0339(.A(new_n528), .B(new_n529), .C1(new_n539), .C2(new_n281), .ZN(new_n540));
  OAI211_X1 g0340(.A(G244), .B(new_n257), .C1(new_n351), .C2(new_n352), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT77), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT4), .ZN(new_n544));
  OAI21_X1  g0344(.A(G250), .B1(new_n351), .B2(new_n352), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT4), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G1698), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n542), .B(new_n546), .C1(new_n353), .C2(new_n208), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n544), .A2(new_n549), .A3(new_n502), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n262), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n434), .A2(G257), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n552), .A2(G190), .A3(new_n445), .A4(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n553), .ZN(new_n555));
  AOI211_X1 g0355(.A(new_n446), .B(new_n555), .C1(new_n551), .C2(new_n262), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n540), .B(new_n554), .C1(new_n556), .C2(new_n325), .ZN(new_n557));
  INV_X1    g0357(.A(G179), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n552), .A2(new_n558), .A3(new_n445), .A4(new_n553), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n539), .A2(new_n281), .ZN(new_n560));
  INV_X1    g0360(.A(new_n528), .ZN(new_n561));
  INV_X1    g0361(.A(new_n529), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n559), .B(new_n563), .C1(new_n556), .C2(G169), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n208), .A2(G1698), .ZN(new_n565));
  OAI221_X1 g0365(.A(new_n565), .B1(G238), .B2(G1698), .C1(new_n351), .C2(new_n352), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n261), .B1(new_n566), .B2(new_n449), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n440), .A2(new_n265), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n261), .A2(G250), .A3(new_n440), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NOR4_X1   g0370(.A1(new_n567), .A2(new_n335), .A3(new_n568), .A4(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n568), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n566), .A2(new_n449), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n572), .B(new_n569), .C1(new_n573), .C2(new_n261), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n571), .B1(new_n574), .B2(new_n330), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n220), .B1(new_n294), .B2(new_n216), .ZN(new_n576));
  INV_X1    g0376(.A(G87), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n533), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n578), .A3(KEYINPUT19), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT19), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n275), .B2(new_n216), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n220), .B(G68), .C1(new_n351), .C2(new_n352), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(new_n281), .B1(new_n378), .B2(new_n274), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n471), .A2(G87), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n274), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n471), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n574), .A2(new_n288), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n558), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n575), .A2(new_n586), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n557), .A2(new_n564), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n479), .A2(new_n335), .A3(new_n445), .A4(new_n480), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n447), .B2(G200), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n468), .A2(new_n281), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n471), .A2(G107), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .A4(new_n476), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT83), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n472), .A2(KEYINPUT83), .A3(new_n476), .A4(new_n595), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n593), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n527), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n430), .A2(new_n604), .ZN(G372));
  AND3_X1   g0405(.A1(new_n509), .A2(new_n514), .A3(new_n522), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n484), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(new_n593), .A3(new_n602), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n589), .A2(new_n591), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n575), .A2(new_n586), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n609), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT26), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n612), .A2(new_n564), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n612), .B2(new_n564), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT84), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n617), .B(new_n613), .C1(new_n612), .C2(new_n564), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n614), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n610), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n430), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g0421(.A(new_n621), .B(KEYINPUT85), .Z(new_n622));
  NOR2_X1   g0422(.A1(new_n401), .A2(new_n400), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n326), .A2(new_n291), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n321), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n623), .B1(new_n625), .B2(new_n394), .ZN(new_n626));
  INV_X1    g0426(.A(new_n426), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n428), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT86), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n622), .A2(new_n630), .ZN(G369));
  INV_X1    g0431(.A(G13), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(G20), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n219), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n634), .A2(KEYINPUT27), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(KEYINPUT27), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(G213), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(G343), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n506), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n640), .B(KEYINPUT87), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n606), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n507), .A2(new_n508), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT21), .B1(new_n513), .B2(new_n506), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n645), .A2(KEYINPUT79), .A3(new_n522), .A4(new_n521), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n523), .A2(new_n524), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n642), .B1(new_n648), .B2(new_n641), .ZN(new_n649));
  INV_X1    g0449(.A(G330), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT88), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n484), .A2(new_n639), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n639), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n472), .B2(new_n476), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n600), .B2(new_n601), .ZN(new_n657));
  AOI211_X1 g0457(.A(new_n448), .B(new_n482), .C1(new_n472), .C2(new_n476), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n652), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n606), .A2(new_n639), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n654), .B(new_n661), .C1(new_n657), .C2(new_n658), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n654), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n660), .A2(new_n663), .ZN(G399));
  INV_X1    g0464(.A(new_n227), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G41), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n578), .A2(G116), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G1), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n234), .B2(new_n667), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  INV_X1    g0471(.A(new_n615), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n608), .B(new_n609), .C1(new_n614), .C2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n655), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT29), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n620), .A2(new_n655), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(KEYINPUT29), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n497), .A2(new_n481), .A3(new_n558), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n555), .B1(new_n551), .B2(new_n262), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n679), .A3(new_n590), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n497), .A2(new_n574), .A3(new_n558), .ZN(new_n683));
  OR3_X1    g0483(.A1(new_n556), .A2(new_n447), .A3(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n678), .A2(KEYINPUT30), .A3(new_n679), .A4(new_n590), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT31), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n686), .A2(new_n687), .A3(new_n639), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n687), .B1(new_n686), .B2(new_n639), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n658), .B1(new_n646), .B2(new_n647), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(new_n602), .A3(new_n593), .A4(new_n655), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT89), .ZN(new_n693));
  INV_X1    g0493(.A(new_n603), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT89), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(new_n691), .A4(new_n655), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n690), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(new_n650), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n677), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n671), .B1(new_n699), .B2(G1), .ZN(G364));
  AOI21_X1  g0500(.A(new_n231), .B1(G20), .B2(new_n288), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n330), .A2(new_n558), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT92), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G20), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G190), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n705), .A2(new_n335), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n709), .A2(KEYINPUT93), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(KEYINPUT93), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI221_X1 g0512(.A(new_n256), .B1(new_n473), .B2(new_n707), .C1(new_n712), .C2(new_n577), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT94), .ZN(new_n714));
  NOR2_X1   g0514(.A1(G190), .A2(G200), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(G20), .A3(new_n558), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G159), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT32), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n335), .A2(G200), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n558), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G97), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n220), .A2(new_n558), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n724), .A2(KEYINPUT91), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(KEYINPUT91), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(new_n715), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n725), .A2(new_n726), .A3(new_n720), .ZN(new_n728));
  OAI221_X1 g0528(.A(new_n723), .B1(new_n727), .B2(new_n207), .C1(new_n345), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n724), .A2(G200), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n335), .ZN(new_n731));
  AOI211_X1 g0531(.A(new_n719), .B(new_n729), .C1(G50), .C2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n730), .A2(G190), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n714), .B(new_n732), .C1(new_n212), .C2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n353), .B1(new_n712), .B2(new_n485), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n736), .A2(KEYINPUT95), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n731), .A2(G326), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n736), .A2(KEYINPUT95), .ZN(new_n739));
  INV_X1    g0539(.A(new_n727), .ZN(new_n740));
  INV_X1    g0540(.A(new_n728), .ZN(new_n741));
  AOI22_X1  g0541(.A1(G311), .A2(new_n740), .B1(new_n741), .B2(G322), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n722), .A2(G294), .B1(new_n717), .B2(G329), .ZN(new_n743));
  XOR2_X1   g0543(.A(KEYINPUT33), .B(G317), .Z(new_n744));
  OAI211_X1 g0544(.A(new_n742), .B(new_n743), .C1(new_n734), .C2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n706), .B2(G283), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n737), .A2(new_n738), .A3(new_n739), .A4(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n702), .B1(new_n735), .B2(new_n747), .ZN(new_n748));
  OR3_X1    g0548(.A1(KEYINPUT90), .A2(G13), .A3(G33), .ZN(new_n749));
  OAI21_X1  g0549(.A(KEYINPUT90), .B1(G13), .B2(G33), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n701), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n227), .A2(G355), .A3(new_n256), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n252), .A2(G45), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n665), .A2(new_n256), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(new_n235), .B2(G45), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n755), .B1(G116), .B2(new_n227), .C1(new_n756), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n748), .B1(new_n754), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n649), .A2(new_n753), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n219), .B1(new_n633), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n666), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n649), .B2(new_n650), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n762), .A2(new_n765), .B1(new_n652), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(G396));
  NOR2_X1   g0568(.A1(new_n290), .A2(new_n639), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n286), .A2(new_n655), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n334), .B2(new_n336), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n770), .B1(new_n772), .B2(new_n291), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n676), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n771), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n337), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n769), .B1(new_n776), .B2(new_n290), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n777), .B(new_n655), .C1(new_n610), .C2(new_n619), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(new_n698), .ZN(new_n780));
  INV_X1    g0580(.A(new_n765), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n722), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n741), .A2(G143), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n733), .A2(G150), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G137), .ZN(new_n787));
  INV_X1    g0587(.A(new_n731), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n786), .B1(new_n787), .B2(new_n788), .C1(new_n789), .C2(new_n727), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT34), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n256), .B1(new_n345), .B2(new_n783), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n707), .A2(new_n212), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n792), .B(new_n793), .C1(new_n791), .C2(new_n790), .ZN(new_n794));
  INV_X1    g0594(.A(G132), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n794), .B1(new_n202), .B2(new_n712), .C1(new_n795), .C2(new_n716), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n740), .A2(G116), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n256), .B1(new_n717), .B2(G311), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n733), .A2(G283), .B1(new_n731), .B2(G303), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n797), .A2(new_n723), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n706), .B2(G87), .ZN(new_n801));
  INV_X1    g0601(.A(G294), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n801), .B1(new_n802), .B2(new_n728), .C1(new_n712), .C2(new_n473), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n796), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n781), .B1(new_n804), .B2(new_n701), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n751), .A2(new_n701), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n805), .B1(G77), .B2(new_n807), .C1(new_n752), .C2(new_n777), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n782), .A2(new_n808), .ZN(G384));
  NAND4_X1  g0609(.A1(new_n366), .A2(new_n558), .A3(new_n368), .A4(new_n267), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n371), .B2(G169), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n359), .A2(new_n388), .B1(new_n811), .B2(new_n637), .ZN(new_n812));
  AND3_X1   g0612(.A1(new_n359), .A2(new_n372), .A3(new_n388), .ZN(new_n813));
  OAI21_X1  g0613(.A(KEYINPUT37), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND3_X1   g0614(.A1(new_n350), .A2(new_n358), .A3(new_n281), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n384), .A2(new_n387), .ZN(new_n816));
  INV_X1    g0616(.A(new_n637), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n815), .A2(new_n816), .B1(new_n399), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT37), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n818), .A2(new_n819), .A3(new_n391), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT96), .ZN(new_n821));
  AND3_X1   g0621(.A1(new_n814), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(new_n814), .B2(new_n820), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n637), .B1(new_n359), .B2(new_n388), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n623), .B2(new_n393), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n824), .A2(KEYINPUT97), .A3(KEYINPUT38), .A4(new_n826), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n812), .A2(new_n813), .A3(KEYINPUT37), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n819), .B1(new_n818), .B2(new_n391), .ZN(new_n829));
  OAI21_X1  g0629(.A(KEYINPUT96), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n814), .A2(new_n820), .A3(new_n821), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n826), .A2(new_n830), .A3(KEYINPUT38), .A4(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT97), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n826), .B1(new_n829), .B2(new_n828), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT38), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT39), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n827), .A2(new_n834), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT38), .B1(new_n824), .B2(new_n826), .ZN(new_n840));
  INV_X1    g0640(.A(new_n832), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT39), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT98), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n321), .A2(new_n639), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT98), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n839), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n844), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n623), .A2(new_n637), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n778), .A2(new_n770), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n840), .A2(new_n841), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n320), .A2(new_n639), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n321), .A2(new_n326), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n853), .B1(new_n321), .B2(new_n326), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n850), .A2(new_n852), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n848), .A2(new_n849), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n430), .A2(new_n677), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n630), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n859), .B(new_n861), .Z(new_n862));
  INV_X1    g0662(.A(new_n690), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n695), .B1(new_n604), .B2(new_n655), .ZN(new_n864));
  NOR4_X1   g0664(.A1(new_n527), .A2(new_n603), .A3(KEYINPUT89), .A4(new_n639), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n827), .A2(new_n834), .A3(new_n837), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n777), .B1(new_n854), .B2(new_n855), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n866), .A2(KEYINPUT40), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n693), .A2(new_n696), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n868), .B1(new_n872), .B2(new_n863), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT40), .B1(new_n873), .B2(new_n852), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n430), .A2(new_n866), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n875), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(G330), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n862), .B(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n219), .B2(new_n633), .ZN(new_n880));
  OAI211_X1 g0680(.A(G20), .B(new_n232), .C1(new_n536), .C2(KEYINPUT35), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n498), .B(new_n881), .C1(KEYINPUT35), .C2(new_n536), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT36), .Z(new_n883));
  OAI21_X1  g0683(.A(G77), .B1(new_n345), .B2(new_n212), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n884), .A2(new_n234), .B1(G50), .B2(new_n212), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(G1), .A3(new_n632), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n880), .A2(new_n883), .A3(new_n886), .ZN(G367));
  OR2_X1    g0687(.A1(new_n564), .A2(new_n655), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n557), .B(new_n564), .C1(new_n540), .C2(new_n655), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n660), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT42), .ZN(new_n892));
  INV_X1    g0692(.A(new_n890), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n662), .A2(new_n893), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n894), .A2(KEYINPUT101), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(KEYINPUT101), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n892), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT102), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n564), .B1(new_n889), .B2(new_n484), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT100), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(new_n639), .ZN(new_n901));
  OR3_X1    g0701(.A1(new_n897), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n898), .B1(new_n897), .B2(new_n901), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n895), .A2(new_n892), .A3(new_n896), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n586), .A2(new_n655), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n592), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n609), .B2(new_n906), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT99), .Z(new_n912));
  INV_X1    g0712(.A(KEYINPUT103), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n891), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n910), .A2(new_n891), .A3(new_n914), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n916), .B(new_n917), .C1(new_n913), .C2(new_n912), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n912), .A2(new_n913), .ZN(new_n919));
  INV_X1    g0719(.A(new_n917), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n919), .B1(new_n920), .B2(new_n915), .ZN(new_n921));
  INV_X1    g0721(.A(new_n699), .ZN(new_n922));
  INV_X1    g0722(.A(new_n660), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n652), .A2(new_n659), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n925), .A2(new_n661), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n661), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n663), .A2(new_n893), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT44), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n929), .B(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n663), .A2(new_n893), .ZN(new_n932));
  XNOR2_X1  g0732(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n923), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n923), .B1(new_n931), .B2(new_n934), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n922), .B1(new_n928), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n666), .B(KEYINPUT41), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n763), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n918), .A2(new_n921), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n712), .A2(new_n498), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(KEYINPUT46), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT106), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n707), .A2(new_n216), .ZN(new_n946));
  INV_X1    g0746(.A(G311), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n353), .B1(new_n788), .B2(new_n947), .C1(new_n802), .C2(new_n734), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(G303), .B2(new_n741), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n740), .A2(G283), .B1(G107), .B2(new_n722), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT105), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(KEYINPUT105), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n946), .B(new_n953), .C1(new_n943), .C2(KEYINPUT46), .ZN(new_n954));
  INV_X1    g0754(.A(G317), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n945), .B(new_n954), .C1(new_n955), .C2(new_n716), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n202), .A2(new_n727), .B1(new_n728), .B2(new_n409), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n353), .B(new_n957), .C1(G68), .C2(new_n722), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n733), .A2(G159), .B1(new_n731), .B2(G143), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n787), .B2(new_n716), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(new_n706), .B2(G77), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n958), .B(new_n961), .C1(new_n712), .C2(new_n345), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n956), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT47), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n701), .ZN(new_n965));
  INV_X1    g0765(.A(new_n757), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n754), .B1(new_n227), .B2(new_n274), .C1(new_n966), .C2(new_n244), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n907), .B(new_n753), .C1(new_n609), .C2(new_n906), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n965), .A2(new_n765), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n942), .A2(new_n969), .ZN(G387));
  OAI211_X1 g0770(.A(new_n668), .B(new_n432), .C1(new_n212), .C2(new_n207), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT107), .Z(new_n972));
  NOR2_X1   g0772(.A1(new_n278), .A2(G50), .ZN(new_n973));
  XOR2_X1   g0773(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n757), .B1(new_n241), .B2(new_n432), .C1(new_n972), .C2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n227), .A2(new_n256), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n976), .B1(G107), .B2(new_n227), .C1(new_n668), .C2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n754), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n733), .A2(G311), .B1(new_n731), .B2(G322), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT109), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n485), .B2(new_n727), .C1(new_n955), .C2(new_n728), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT48), .ZN(new_n983));
  INV_X1    g0783(.A(G283), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n983), .B1(new_n984), .B2(new_n783), .C1(new_n802), .C2(new_n712), .ZN(new_n985));
  XNOR2_X1  g0785(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n717), .A2(G326), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n985), .A2(new_n986), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n256), .B1(new_n706), .B2(G116), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n353), .B1(new_n717), .B2(G150), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n722), .A2(new_n587), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n788), .C2(new_n789), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n410), .A2(new_n734), .B1(new_n727), .B2(new_n212), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(G50), .C2(new_n741), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n216), .B2(new_n707), .C1(new_n712), .C2(new_n207), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n702), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n659), .A2(new_n753), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n998), .A2(new_n781), .A3(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n928), .A2(new_n764), .B1(new_n979), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n926), .A2(new_n922), .A3(new_n927), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n666), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n922), .B1(new_n926), .B2(new_n927), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(G393));
  OR3_X1    g0805(.A1(new_n1004), .A2(KEYINPUT112), .A3(new_n937), .ZN(new_n1006));
  OAI21_X1  g0806(.A(KEYINPUT112), .B1(new_n1004), .B2(new_n937), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n937), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n666), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n937), .A2(new_n764), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n947), .A2(new_n728), .B1(new_n788), .B2(new_n955), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT52), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n353), .B1(new_n734), .B2(new_n485), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G116), .B2(new_n722), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(new_n802), .C2(new_n727), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1013), .B(new_n1017), .C1(G107), .C2(new_n706), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n717), .A2(G322), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(new_n984), .C2(new_n712), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n783), .A2(new_n207), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n353), .B1(new_n717), .B2(G143), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n278), .A2(new_n727), .B1(new_n734), .B2(new_n202), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1022), .B1(new_n1023), .B2(KEYINPUT111), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1021), .B(new_n1024), .C1(KEYINPUT111), .C2(new_n1023), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n577), .B2(new_n707), .C1(new_n712), .C2(new_n212), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n741), .A2(G159), .B1(G150), .B2(new_n731), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT51), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1020), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n781), .B1(new_n1029), .B2(new_n701), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n754), .B1(new_n216), .B2(new_n227), .C1(new_n249), .C2(new_n966), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n893), .A2(new_n753), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1009), .A2(new_n1010), .A3(new_n1033), .ZN(G390));
  INV_X1    g0834(.A(new_n845), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n850), .A2(new_n857), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n844), .A2(new_n847), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n867), .A2(new_n1035), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n673), .B(new_n655), .C1(new_n291), .C2(new_n772), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n770), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1038), .B1(new_n1040), .B2(new_n857), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT113), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1036), .A2(new_n1035), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n846), .B1(new_n839), .B2(new_n842), .ZN(new_n1044));
  AND3_X1   g0844(.A1(new_n839), .A2(new_n842), .A3(new_n846), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT113), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1041), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n698), .A2(new_n869), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1042), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  OAI211_X1 g0852(.A(KEYINPUT113), .B(new_n1050), .C1(new_n1037), .C2(new_n1041), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n763), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n751), .B1(new_n1045), .B2(new_n1044), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n410), .A2(new_n806), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n712), .A2(new_n409), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT53), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n731), .A2(G128), .B1(G125), .B2(new_n717), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n787), .B2(new_n734), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(KEYINPUT54), .B(G143), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n795), .A2(new_n728), .B1(new_n727), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n353), .B1(new_n706), .B2(G50), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT114), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n1065), .B2(new_n1064), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1058), .B(new_n1067), .C1(new_n789), .C2(new_n783), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n734), .A2(new_n473), .B1(new_n788), .B2(new_n984), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n353), .B1(new_n716), .B2(new_n802), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1069), .A2(new_n1021), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n216), .B2(new_n727), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G116), .B2(new_n741), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n712), .B2(new_n577), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1068), .B1(new_n793), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n781), .B1(new_n1075), .B2(new_n701), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1055), .A2(new_n1056), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  OR3_X1    g0878(.A1(new_n1054), .A2(KEYINPUT115), .A3(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(KEYINPUT115), .B1(new_n1054), .B2(new_n1078), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n630), .B(new_n860), .C1(new_n650), .C2(new_n876), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n697), .A2(new_n650), .A3(new_n773), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1050), .B1(new_n1084), .B2(new_n857), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n850), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1040), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1050), .B(new_n1087), .C1(new_n857), .C2(new_n1084), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1083), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1081), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1090), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1092), .A2(new_n1093), .A3(new_n666), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1079), .A2(new_n1080), .A3(new_n1094), .ZN(G378));
  INV_X1    g0895(.A(KEYINPUT119), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n697), .A2(new_n851), .A3(new_n868), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n870), .B(G330), .C1(new_n1097), .C2(KEYINPUT40), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT118), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n852), .A2(new_n866), .A3(new_n869), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT40), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1103), .A2(KEYINPUT118), .A3(G330), .A4(new_n870), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n412), .A2(new_n637), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT55), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n426), .A2(new_n1106), .A3(new_n428), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1106), .B1(new_n426), .B2(new_n428), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1105), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1109), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1105), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1114), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1100), .A2(new_n1104), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1114), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n875), .A2(KEYINPUT118), .A3(new_n1123), .A4(G330), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1118), .A2(new_n859), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n859), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1096), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1117), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1124), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n859), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1118), .A2(new_n859), .A3(new_n1124), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(KEYINPUT119), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1127), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1092), .A2(new_n1083), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT57), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(KEYINPUT57), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1082), .B1(new_n1081), .B2(new_n1089), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n666), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n727), .A2(new_n787), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n731), .A2(G125), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n734), .B2(new_n795), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1143), .B(new_n1145), .C1(G128), .C2(new_n741), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n409), .B2(new_n783), .C1(new_n712), .C2(new_n1061), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT59), .Z(new_n1148));
  AOI21_X1  g0948(.A(G41), .B1(new_n706), .B2(G159), .ZN(new_n1149));
  AOI21_X1  g0949(.A(G33), .B1(new_n717), .B2(G124), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n706), .A2(G58), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT116), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n734), .A2(new_n216), .B1(new_n788), .B2(new_n498), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G68), .B2(new_n722), .ZN(new_n1155));
  AOI211_X1 g0955(.A(G41), .B(new_n256), .C1(new_n717), .C2(G283), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(new_n473), .C2(new_n728), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n587), .B2(new_n740), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1153), .B(new_n1158), .C1(new_n712), .C2(new_n207), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT58), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n202), .B1(new_n351), .B2(G41), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1151), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n765), .B1(new_n1162), .B2(new_n702), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1117), .A2(new_n752), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n202), .C2(new_n806), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n1135), .B2(new_n764), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1142), .A2(new_n1166), .ZN(G375));
  NAND2_X1  g0967(.A1(new_n740), .A2(G107), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n256), .B1(new_n717), .B2(G303), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n733), .A2(G116), .B1(new_n731), .B2(G294), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1168), .A2(new_n993), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n706), .B2(G77), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n984), .B2(new_n728), .C1(new_n712), .C2(new_n216), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT121), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n710), .A2(G159), .A3(new_n711), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n717), .A2(G128), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n787), .A2(new_n728), .B1(new_n727), .B2(new_n409), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n788), .A2(new_n795), .B1(new_n783), .B2(new_n202), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n256), .B1(new_n734), .B2(new_n1061), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1175), .A2(new_n1153), .A3(new_n1176), .A4(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n702), .B1(new_n1174), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n857), .A2(new_n752), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n807), .A2(G68), .ZN(new_n1184));
  NOR4_X1   g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n781), .A4(new_n1184), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n763), .B(KEYINPUT120), .Z(new_n1186));
  AOI21_X1  g0986(.A(new_n1185), .B1(new_n1089), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n939), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n1091), .B2(new_n1188), .ZN(G381));
  NOR2_X1   g0989(.A1(G375), .A2(G378), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1191), .A2(G384), .A3(G381), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(G387), .A2(G390), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(G393), .A2(G396), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(G407));
  NAND2_X1  g0995(.A1(new_n638), .A2(G213), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT122), .Z(new_n1197));
  OAI211_X1 g0997(.A(G407), .B(G213), .C1(new_n1191), .C2(new_n1197), .ZN(G409));
  NOR3_X1   g0998(.A1(new_n1125), .A2(new_n1126), .A3(new_n1096), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT119), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n939), .B(new_n1136), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1165), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1138), .A2(new_n1186), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(G378), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(G378), .B(new_n1166), .C1(new_n1137), .C2(new_n1141), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(KEYINPUT123), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n667), .B1(new_n1209), .B2(KEYINPUT60), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1210), .B(new_n1090), .C1(KEYINPUT60), .C2(new_n1209), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n1187), .ZN(new_n1212));
  INV_X1    g1012(.A(G384), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1211), .A2(G384), .A3(new_n1187), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1208), .A2(new_n1196), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT62), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1214), .A2(KEYINPUT62), .A3(new_n1215), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1208), .A2(new_n1197), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT126), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1208), .A2(new_n1221), .A3(KEYINPUT126), .A4(new_n1197), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1220), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n638), .A2(G213), .A3(G2897), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1214), .A2(new_n1215), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT124), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1214), .A2(KEYINPUT124), .A3(new_n1215), .A4(new_n1227), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1197), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1230), .A2(new_n1231), .B1(G2897), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1208), .A2(new_n1197), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT61), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1226), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT127), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G387), .A2(G390), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1009), .A2(new_n1010), .A3(new_n1033), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(new_n942), .A3(new_n969), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT125), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1238), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G393), .A2(G396), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n1242), .A2(new_n1243), .B1(new_n1194), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT125), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1245), .A2(new_n1194), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1238), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1246), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT127), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1226), .A2(new_n1253), .A3(new_n1235), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1237), .A2(new_n1252), .A3(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT63), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1234), .A2(new_n1256), .A3(new_n1216), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1252), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1218), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1208), .A2(new_n1196), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1256), .B1(new_n1233), .B2(new_n1261), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1258), .B(new_n1259), .C1(new_n1260), .C2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1255), .A2(new_n1263), .ZN(G405));
  AOI21_X1  g1064(.A(G378), .B1(new_n1142), .B2(new_n1166), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1207), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(new_n1216), .ZN(new_n1268));
  XOR2_X1   g1068(.A(new_n1268), .B(new_n1252), .Z(G402));
endmodule


