//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G235), .A3(G237), .A4(G238), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT66), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n472), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n461), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n469), .A2(G136), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n461), .B1(new_n467), .B2(new_n468), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI211_X1 g059(.A(G138), .B(new_n461), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n472), .A2(KEYINPUT67), .A3(G138), .A4(new_n461), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n483), .C2(new_n484), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  AND4_X1   g072(.A1(KEYINPUT68), .A2(new_n489), .A3(new_n491), .A4(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(KEYINPUT67), .B1(new_n469), .B2(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n496), .B1(new_n499), .B2(new_n490), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT68), .B1(new_n500), .B2(new_n489), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n498), .A2(new_n501), .ZN(G164));
  OR2_X1    g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n510), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(KEYINPUT69), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(new_n512), .B2(G50), .ZN(new_n516));
  OAI221_X1 g091(.A(new_n508), .B1(new_n509), .B2(new_n511), .C1(new_n514), .C2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  XOR2_X1   g093(.A(KEYINPUT70), .B(G89), .Z(new_n519));
  NAND2_X1  g094(.A1(new_n510), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n511), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n522), .A2(new_n526), .ZN(G168));
  INV_X1    g102(.A(G64), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n528), .B1(new_n503), .B2(new_n504), .ZN(new_n529));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  OR3_X1    g106(.A1(new_n529), .A2(KEYINPUT71), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT71), .B1(new_n529), .B2(new_n531), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n532), .A2(G651), .A3(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n505), .A2(new_n510), .ZN(new_n535));
  AOI22_X1  g110(.A1(G90), .A2(new_n535), .B1(new_n512), .B2(G52), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n503), .A2(new_n504), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G651), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n505), .A2(new_n510), .A3(G81), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n510), .A2(G43), .A3(G543), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT72), .ZN(new_n546));
  AOI21_X1  g121(.A(KEYINPUT72), .B1(new_n544), .B2(new_n545), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n543), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND4_X1  g129(.A1(new_n510), .A2(KEYINPUT73), .A3(G53), .A4(G543), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n507), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n535), .A2(G91), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(G299));
  INV_X1    g135(.A(G168), .ZN(G286));
  NAND2_X1  g136(.A1(new_n535), .A2(G87), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n512), .A2(G49), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(G288));
  AOI22_X1  g140(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G48), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n566), .A2(new_n507), .B1(new_n567), .B2(new_n520), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  AND3_X1   g144(.A1(new_n505), .A2(new_n510), .A3(G86), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n570), .A2(KEYINPUT74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(KEYINPUT74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(G305));
  AOI22_X1  g148(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n507), .ZN(new_n575));
  INV_X1    g150(.A(G85), .ZN(new_n576));
  INV_X1    g151(.A(G47), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n511), .A2(new_n576), .B1(new_n520), .B2(new_n577), .ZN(new_n578));
  OR3_X1    g153(.A1(new_n575), .A2(new_n578), .A3(KEYINPUT75), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT75), .B1(new_n575), .B2(new_n578), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G79), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G66), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n540), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(G651), .B1(new_n512), .B2(G54), .ZN(new_n585));
  XNOR2_X1  g160(.A(KEYINPUT77), .B(KEYINPUT10), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n588), .A2(new_n535), .A3(G92), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n586), .B(new_n587), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n505), .A2(new_n510), .A3(G92), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND3_X1   g168(.A1(new_n585), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT76), .B1(new_n594), .B2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  MUX2_X1   g171(.A(KEYINPUT76), .B(new_n595), .S(new_n596), .Z(G284));
  MUX2_X1   g172(.A(KEYINPUT76), .B(new_n595), .S(new_n596), .Z(G321));
  NAND2_X1  g173(.A1(G286), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n558), .A2(new_n559), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT9), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n555), .B(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n599), .B1(new_n603), .B2(G868), .ZN(G297));
  OAI21_X1  g179(.A(new_n599), .B1(new_n603), .B2(G868), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n594), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n594), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n463), .A2(new_n472), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT12), .Z(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT13), .Z(new_n614));
  XOR2_X1   g189(.A(KEYINPUT79), .B(G2100), .Z(new_n615));
  OR2_X1    g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n469), .A2(G135), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n477), .A2(G123), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n461), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(G2096), .Z(new_n623));
  NAND3_X1  g198(.A1(new_n616), .A2(new_n617), .A3(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n628), .A2(KEYINPUT14), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2443), .B(G2446), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n630), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G2451), .B(G2454), .Z(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n634), .A2(new_n637), .ZN(new_n639));
  AND3_X1   g214(.A1(new_n638), .A2(G14), .A3(new_n639), .ZN(G401));
  XOR2_X1   g215(.A(G2072), .B(G2078), .Z(new_n641));
  AND2_X1   g216(.A1(new_n641), .A2(KEYINPUT82), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  NOR3_X1   g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(KEYINPUT82), .B2(new_n641), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n641), .A2(KEYINPUT17), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n641), .A2(KEYINPUT17), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n647), .B(new_n648), .C1(new_n643), .C2(new_n644), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n643), .A2(new_n644), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n641), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT81), .B(KEYINPUT18), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2096), .B(G2100), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(G227));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  AND2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT20), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n659), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n659), .B2(new_n665), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G229));
  INV_X1    g249(.A(KEYINPUT98), .ZN(new_n675));
  INV_X1    g250(.A(G1986), .ZN(new_n676));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n677), .A2(G24), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(G290), .B2(G16), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n676), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n685), .A2(G1986), .A3(new_n681), .ZN(new_n686));
  NOR2_X1   g261(.A1(G25), .A2(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n469), .A2(G131), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n477), .A2(G119), .ZN(new_n689));
  OR2_X1    g264(.A1(G95), .A2(G2105), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n690), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n687), .B1(new_n693), .B2(G29), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT35), .B(G1991), .Z(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT83), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n694), .B(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n684), .A2(new_n686), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G1971), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n677), .A2(G22), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G303), .B2(G16), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT87), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n701), .A2(new_n702), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n699), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n701), .A2(new_n702), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n707), .A2(G1971), .A3(new_n703), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n677), .A2(G23), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n711));
  NAND2_X1  g286(.A1(G288), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT85), .A4(new_n564), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n710), .B1(new_n714), .B2(new_n677), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT33), .B(G1976), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT86), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(new_n717), .ZN(new_n719));
  MUX2_X1   g294(.A(G6), .B(G305), .S(G16), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT32), .B(G1981), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n718), .A2(new_n719), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n709), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT34), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n698), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT88), .ZN(new_n728));
  AND3_X1   g303(.A1(new_n718), .A2(new_n723), .A3(new_n722), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n729), .A2(new_n719), .A3(new_n708), .A4(new_n706), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n728), .B1(new_n730), .B2(KEYINPUT34), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n728), .B(KEYINPUT34), .C1(new_n709), .C2(new_n724), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n727), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(KEYINPUT36), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT36), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n727), .B(new_n736), .C1(new_n731), .C2(new_n733), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NOR2_X1   g314(.A1(G164), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G27), .B2(new_n739), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT97), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n743), .A2(G2078), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n594), .A2(G16), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G4), .B2(G16), .ZN(new_n747));
  INV_X1    g322(.A(G1348), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n739), .A2(G32), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT26), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n469), .A2(G141), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G105), .B2(new_n463), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n477), .A2(G129), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT93), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n751), .B1(new_n760), .B2(new_n739), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT27), .B(G1996), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n749), .A2(new_n750), .A3(new_n764), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n677), .A2(G21), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G286), .B2(G16), .ZN(new_n767));
  INV_X1    g342(.A(G1966), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT95), .ZN(new_n770));
  AND3_X1   g345(.A1(new_n739), .A2(KEYINPUT28), .A3(G26), .ZN(new_n771));
  AOI21_X1  g346(.A(KEYINPUT28), .B1(new_n739), .B2(G26), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n469), .A2(G140), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n477), .A2(G128), .ZN(new_n774));
  OR2_X1    g349(.A1(G104), .A2(G2105), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n775), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n771), .B(new_n772), .C1(new_n777), .C2(G29), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n767), .A2(new_n768), .B1(G2067), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT30), .B(G28), .ZN(new_n781));
  OR2_X1    g356(.A1(KEYINPUT31), .A2(G11), .ZN(new_n782));
  NAND2_X1  g357(.A1(KEYINPUT31), .A2(G11), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n781), .A2(new_n739), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n622), .B2(new_n739), .ZN(new_n785));
  INV_X1    g360(.A(G2067), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n785), .B1(new_n778), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n780), .A2(new_n787), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n765), .A2(new_n770), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n677), .A2(G20), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT23), .Z(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G299), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1956), .ZN(new_n793));
  INV_X1    g368(.A(G34), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n794), .A2(KEYINPUT24), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(KEYINPUT24), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n739), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G160), .B2(new_n739), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT92), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n793), .B1(new_n799), .B2(G2084), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n739), .A2(G35), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G162), .B2(new_n739), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT29), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2090), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G5), .A2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT96), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G301), .B2(new_n677), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(G1961), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n677), .A2(G19), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT89), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n549), .B2(new_n677), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1341), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  AND4_X1   g389(.A1(new_n745), .A2(new_n789), .A3(new_n805), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n743), .A2(new_n744), .ZN(new_n816));
  INV_X1    g391(.A(G2078), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT25), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n469), .A2(G139), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n472), .A2(G127), .ZN(new_n824));
  NAND2_X1  g399(.A1(G115), .A2(G2104), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n461), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT90), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT90), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n739), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n739), .A2(G33), .ZN(new_n833));
  OR3_X1    g408(.A1(new_n832), .A2(KEYINPUT91), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(KEYINPUT91), .B1(new_n832), .B2(new_n833), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G2072), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n834), .A2(G2072), .A3(new_n835), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n761), .A2(new_n763), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G2084), .B2(new_n799), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT94), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n815), .B(new_n818), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n675), .B1(new_n738), .B2(new_n847), .ZN(new_n848));
  AOI211_X1 g423(.A(KEYINPUT98), .B(new_n846), .C1(new_n735), .C2(new_n737), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(G311));
  NAND2_X1  g425(.A1(new_n738), .A2(new_n847), .ZN(G150));
  NAND3_X1  g426(.A1(new_n585), .A2(new_n593), .A3(new_n590), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(new_n606), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(new_n507), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT100), .B(G93), .ZN(new_n858));
  INV_X1    g433(.A(G55), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n511), .A2(new_n858), .B1(new_n520), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n548), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n857), .A2(new_n860), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n862), .B(new_n543), .C1(new_n547), .C2(new_n546), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n855), .B(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n867));
  INV_X1    g442(.A(G860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n862), .A2(new_n868), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT37), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(G145));
  XNOR2_X1  g448(.A(G160), .B(new_n622), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(G162), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n489), .A2(new_n491), .A3(new_n497), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n777), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n877), .A2(new_n759), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n759), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n828), .A2(KEYINPUT101), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n828), .A2(KEYINPUT90), .A3(KEYINPUT101), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n878), .A2(new_n831), .A3(new_n879), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n477), .A2(G130), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT102), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n889));
  INV_X1    g464(.A(G118), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n889), .B1(new_n890), .B2(G2105), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(G142), .B2(new_n469), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n883), .A2(new_n885), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n894), .B1(new_n883), .B2(new_n885), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n613), .B(new_n693), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n885), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n881), .B1(new_n878), .B2(new_n879), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n893), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n898), .B1(new_n903), .B2(new_n895), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n875), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n899), .B1(new_n896), .B2(new_n897), .ZN(new_n907));
  INV_X1    g482(.A(new_n875), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n903), .A2(new_n898), .A3(new_n895), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n907), .A2(new_n909), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n914), .B2(new_n875), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(KEYINPUT103), .A3(new_n910), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n913), .A2(KEYINPUT40), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT40), .B1(new_n913), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(G395));
  INV_X1    g494(.A(G290), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(G303), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n714), .A2(G305), .ZN(new_n922));
  NAND2_X1  g497(.A1(G166), .A2(G290), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n714), .A2(G305), .ZN(new_n924));
  AND4_X1   g499(.A1(new_n921), .A2(new_n922), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  AOI22_X1  g500(.A1(new_n924), .A2(new_n922), .B1(new_n921), .B2(new_n923), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT42), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n864), .B(new_n608), .Z(new_n929));
  OAI21_X1  g504(.A(KEYINPUT104), .B1(new_n594), .B2(G299), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n603), .A2(new_n931), .A3(new_n852), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n594), .A2(G299), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT41), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n930), .A2(new_n932), .A3(KEYINPUT41), .A4(new_n933), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n936), .B1(new_n929), .B2(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n928), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n928), .A2(new_n941), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(G868), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n862), .A2(G868), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G868), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n942), .B2(new_n943), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT105), .B1(new_n951), .B2(new_n947), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(G295));
  NAND2_X1  g528(.A1(new_n945), .A2(new_n948), .ZN(G331));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n925), .A2(new_n926), .ZN(new_n957));
  NAND2_X1  g532(.A1(G301), .A2(G286), .ZN(new_n958));
  NAND3_X1  g533(.A1(G168), .A2(new_n534), .A3(new_n536), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n864), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n861), .A2(new_n958), .A3(new_n863), .A4(new_n959), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n934), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n934), .A2(new_n961), .A3(KEYINPUT107), .A4(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n968));
  AND4_X1   g543(.A1(new_n861), .A2(new_n958), .A3(new_n863), .A4(new_n959), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n863), .A2(new_n861), .B1(new_n958), .B2(new_n959), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n962), .A2(KEYINPUT106), .ZN(new_n972));
  AOI22_X1  g547(.A1(new_n971), .A2(new_n972), .B1(new_n938), .B2(new_n939), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n957), .B1(new_n967), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n975), .A3(new_n906), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n965), .A2(new_n966), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n971), .A2(new_n972), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n940), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n927), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n975), .B1(new_n974), .B2(new_n906), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT43), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n980), .A2(new_n906), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n935), .A2(KEYINPUT110), .A3(KEYINPUT41), .ZN(new_n985));
  OAI221_X1 g560(.A(new_n985), .B1(new_n969), .B2(new_n970), .C1(new_n940), .C2(KEYINPUT110), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n971), .A2(new_n934), .A3(new_n972), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n927), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OR3_X1    g563(.A1(new_n984), .A2(new_n988), .A3(KEYINPUT43), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n956), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n982), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(new_n980), .A3(new_n976), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT109), .B1(new_n992), .B2(KEYINPUT43), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n955), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n984), .A2(new_n988), .A3(new_n995), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT44), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n994), .A2(new_n998), .ZN(G397));
  INV_X1    g574(.A(G1384), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n876), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n473), .A2(new_n461), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1004), .A2(G40), .A3(new_n464), .A4(new_n470), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1007), .A2(new_n676), .A3(new_n920), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1007), .A2(G1986), .A3(G290), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT111), .ZN(new_n1011));
  INV_X1    g586(.A(G1996), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n760), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n777), .B(new_n786), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n759), .A2(G1996), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n692), .B(new_n695), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1007), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1011), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1384), .B1(new_n500), .B2(new_n489), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1005), .B1(new_n1021), .B2(KEYINPUT45), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT68), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n876), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n500), .A2(KEYINPUT68), .A3(new_n489), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1384), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1022), .B1(new_n1026), .B2(KEYINPUT45), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(KEYINPUT112), .B(new_n1022), .C1(new_n1026), .C2(KEYINPUT45), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(new_n699), .A3(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(KEYINPUT50), .B(new_n1000), .C1(new_n498), .C2(new_n501), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1021), .A2(KEYINPUT50), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1005), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G2090), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1031), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G303), .A2(G8), .ZN(new_n1039));
  NAND2_X1  g614(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1038), .A2(G8), .A3(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1045));
  INV_X1    g620(.A(G8), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1981), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n569), .A2(new_n571), .A3(new_n1048), .A4(new_n572), .ZN(new_n1049));
  OAI21_X1  g624(.A(G1981), .B1(new_n568), .B2(new_n570), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(KEYINPUT49), .A3(new_n1050), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1047), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n712), .A2(G1976), .A3(new_n713), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1056), .B(G8), .C1(new_n1005), .C2(new_n1001), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT52), .ZN(new_n1058));
  XOR2_X1   g633(.A(KEYINPUT114), .B(G1976), .Z(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(G288), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1047), .A2(new_n1056), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1055), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1055), .A2(new_n1058), .A3(new_n1061), .A4(KEYINPUT116), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n876), .B2(new_n1000), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1069), .B2(new_n1005), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1068), .B(new_n1000), .C1(new_n498), .C2(new_n501), .ZN(new_n1071));
  INV_X1    g646(.A(G40), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n471), .A2(new_n1072), .A3(new_n474), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(KEYINPUT115), .C1(new_n1021), .C2(new_n1068), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1070), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1075), .A2(G2090), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1046), .B1(new_n1031), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1044), .B(new_n1066), .C1(new_n1043), .C2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G2084), .ZN(new_n1079));
  AOI211_X1 g654(.A(new_n1068), .B(G1384), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1079), .B(new_n1073), .C1(new_n1080), .C2(new_n1033), .ZN(new_n1081));
  AOI211_X1 g656(.A(new_n1002), .B(G1384), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1003), .A2(new_n1073), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n768), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(G168), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1085), .A2(new_n1086), .A3(G8), .ZN(new_n1087));
  AOI211_X1 g662(.A(G2084), .B(new_n1005), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1026), .A2(KEYINPUT45), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1005), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1090));
  AOI21_X1  g665(.A(G1966), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(G286), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(G8), .A3(new_n1085), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1087), .B1(KEYINPUT51), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1078), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1035), .A2(G1961), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1000), .B1(new_n498), .B2(new_n501), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1002), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT112), .B1(new_n1099), .B2(new_n1022), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1030), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n817), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1097), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1089), .A2(KEYINPUT53), .A3(new_n817), .A4(new_n1090), .ZN(new_n1105));
  AOI21_X1  g680(.A(G301), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1097), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT53), .B1(new_n1108), .B2(G2078), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n1108), .B2(G2078), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1090), .B(new_n1110), .C1(new_n1002), .C2(new_n1001), .ZN(new_n1111));
  AOI21_X1  g686(.A(G2078), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1107), .B(new_n1111), .C1(new_n1112), .C2(KEYINPUT53), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(G171), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1096), .B1(new_n1106), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1104), .A2(G301), .A3(new_n1105), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1113), .A2(G171), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(KEYINPUT54), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1095), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(G2072), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1099), .A2(new_n1022), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(G1956), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1075), .A2(KEYINPUT117), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT117), .B1(new_n1075), .B2(new_n1123), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1122), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n602), .A2(KEYINPUT118), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n602), .A2(KEYINPUT118), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1127), .A2(new_n1128), .A3(new_n600), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n1130));
  OR3_X1    g705(.A1(new_n1129), .A2(new_n1130), .A3(KEYINPUT57), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1129), .B2(KEYINPUT57), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n603), .A2(KEYINPUT57), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1126), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1134), .B(new_n1122), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(KEYINPUT61), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1045), .A2(new_n786), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1035), .B2(G1348), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n594), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n852), .B(new_n1139), .C1(new_n1035), .C2(G1348), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1140), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n852), .A2(KEYINPUT60), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1143), .A2(KEYINPUT60), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1138), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1136), .A2(new_n1148), .A3(new_n1137), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1126), .A2(KEYINPUT124), .A3(new_n1135), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1012), .B(new_n1022), .C1(new_n1026), .C2(KEYINPUT45), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n1156));
  XOR2_X1   g731(.A(KEYINPUT58), .B(G1341), .Z(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1155), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1156), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n549), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(KEYINPUT59), .B(new_n549), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1147), .A2(new_n1152), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1141), .B(KEYINPUT121), .Z(new_n1166));
  INV_X1    g741(.A(new_n1136), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1137), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1119), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1078), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1094), .A2(new_n1171), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1085), .A2(G8), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1086), .B1(new_n1173), .B2(new_n1092), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT62), .B1(new_n1174), .B2(new_n1087), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1170), .A2(new_n1172), .A3(new_n1175), .A4(new_n1106), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n1177));
  OAI211_X1 g752(.A(G8), .B(G168), .C1(new_n1088), .C2(new_n1091), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n1078), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1046), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1180), .A2(new_n1043), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1178), .A2(new_n1177), .A3(new_n1062), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1181), .A2(new_n1044), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1044), .A2(new_n1062), .ZN(new_n1185));
  NOR2_X1   g760(.A1(G288), .A2(G1976), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1055), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n1049), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1185), .B1(new_n1047), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1176), .A2(new_n1184), .A3(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1020), .B1(new_n1169), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT46), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1192), .B1(new_n1007), .B2(G1996), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g770(.A(new_n760), .B(new_n1014), .C1(new_n1192), .C2(G1996), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1006), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT47), .ZN(new_n1200));
  OR2_X1    g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1019), .B1(new_n1009), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1204), .B1(new_n1009), .B2(new_n1203), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n693), .A2(new_n695), .ZN(new_n1207));
  OAI22_X1  g782(.A1(new_n1016), .A2(new_n1207), .B1(G2067), .B2(new_n777), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(new_n1006), .ZN(new_n1209));
  AND4_X1   g784(.A1(new_n1201), .A2(new_n1205), .A3(new_n1206), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1191), .A2(new_n1210), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g786(.A1(new_n990), .A2(new_n993), .ZN(new_n1213));
  NOR4_X1   g787(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1214));
  AOI21_X1  g788(.A(KEYINPUT103), .B1(new_n915), .B2(new_n910), .ZN(new_n1215));
  AND4_X1   g789(.A1(KEYINPUT103), .A2(new_n905), .A3(new_n906), .A4(new_n910), .ZN(new_n1216));
  OAI21_X1  g790(.A(new_n1214), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g791(.A1(new_n1213), .A2(new_n1217), .ZN(G308));
  OAI221_X1 g792(.A(new_n1214), .B1(new_n1215), .B2(new_n1216), .C1(new_n990), .C2(new_n993), .ZN(G225));
endmodule


