//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1299, new_n1300, new_n1301, new_n1302, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G97), .A2(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n211), .B(new_n217), .C1(G116), .C2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n205), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n208), .B(new_n228), .C1(new_n231), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT64), .B(G250), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G257), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT65), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT75), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n253), .B(G274), .C1(G41), .C2(G45), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT72), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n254), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT72), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n256), .A2(new_n258), .B1(new_n263), .B2(G238), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT71), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n220), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n225), .A2(G1698), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n267), .B(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G97), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n265), .B1(new_n273), .B2(new_n259), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  OAI211_X1 g0075(.A(G1), .B(G13), .C1(new_n275), .C2(new_n260), .ZN(new_n276));
  AOI211_X1 g0076(.A(KEYINPUT71), .B(new_n276), .C1(new_n271), .C2(new_n272), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n264), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT13), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT13), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n280), .B(new_n264), .C1(new_n274), .C2(new_n277), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(KEYINPUT74), .A3(new_n281), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n274), .A2(new_n277), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT74), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n283), .A2(new_n284), .A3(new_n280), .A4(new_n264), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n252), .B1(new_n286), .B2(G179), .ZN(new_n287));
  INV_X1    g0087(.A(G179), .ZN(new_n288));
  AOI211_X1 g0088(.A(KEYINPUT75), .B(new_n288), .C1(new_n282), .C2(new_n285), .ZN(new_n289));
  INV_X1    g0089(.A(G169), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(new_n279), .B2(new_n281), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(KEYINPUT14), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT14), .ZN(new_n293));
  AOI211_X1 g0093(.A(new_n293), .B(new_n290), .C1(new_n279), .C2(new_n281), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n287), .A2(new_n289), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n229), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n230), .A2(G33), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n298), .A2(new_n221), .B1(new_n230), .B2(G68), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n230), .A2(new_n275), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(new_n219), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n297), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  XOR2_X1   g0102(.A(new_n302), .B(KEYINPUT11), .Z(new_n303));
  NAND3_X1  g0103(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT68), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT68), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n306), .A2(new_n253), .A3(G13), .A4(G20), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n253), .A2(G20), .ZN(new_n309));
  INV_X1    g0109(.A(new_n297), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n213), .B1(new_n311), .B2(KEYINPUT12), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n305), .A2(new_n307), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n313), .A2(KEYINPUT12), .A3(new_n213), .ZN(new_n314));
  INV_X1    g0114(.A(new_n304), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(KEYINPUT12), .ZN(new_n316));
  NOR4_X1   g0116(.A1(new_n303), .A2(new_n312), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n295), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n279), .B2(new_n281), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n321), .B(KEYINPUT73), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n318), .B1(G190), .B2(new_n286), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n263), .A2(G244), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n275), .ZN(new_n327));
  NAND2_X1  g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n266), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n330), .A2(new_n225), .B1(new_n209), .B2(new_n329), .ZN(new_n331));
  OAI21_X1  g0131(.A(G1698), .B1(new_n269), .B2(new_n270), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT67), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT67), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n329), .A2(new_n334), .A3(G1698), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n331), .B1(new_n336), .B2(G238), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n254), .B(new_n325), .C1(new_n337), .C2(new_n276), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n290), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n313), .A2(new_n221), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT8), .B(G58), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n300), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n342), .A2(new_n343), .B1(G20), .B2(G77), .ZN(new_n344));
  XOR2_X1   g0144(.A(KEYINPUT15), .B(G87), .Z(new_n345));
  INV_X1    g0145(.A(new_n298), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n340), .B1(new_n311), .B2(new_n221), .C1(new_n348), .C2(new_n310), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n339), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT69), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n338), .A2(G179), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT69), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n339), .A2(new_n353), .A3(new_n349), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n338), .A2(G200), .ZN(new_n356));
  INV_X1    g0156(.A(G190), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n357), .B2(new_n338), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n358), .A2(new_n349), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n319), .A2(new_n324), .A3(new_n355), .A4(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n269), .A2(new_n270), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT7), .B1(new_n361), .B2(new_n230), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT7), .ZN(new_n363));
  NOR4_X1   g0163(.A1(new_n269), .A2(new_n270), .A3(new_n363), .A4(G20), .ZN(new_n364));
  OAI21_X1  g0164(.A(G68), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n224), .A2(new_n213), .ZN(new_n366));
  NOR2_X1   g0166(.A1(G58), .A2(G68), .ZN(new_n367));
  OAI21_X1  g0167(.A(G20), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n343), .A2(G159), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n310), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT76), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n327), .A2(new_n230), .A3(new_n328), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n363), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n361), .A2(KEYINPUT7), .A3(new_n230), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n370), .B1(new_n379), .B2(G68), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n375), .B1(new_n380), .B2(KEYINPUT16), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n213), .B1(new_n377), .B2(new_n378), .ZN(new_n382));
  NOR4_X1   g0182(.A1(new_n382), .A2(KEYINPUT76), .A3(new_n373), .A4(new_n370), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n374), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n220), .A2(G1698), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n385), .B1(G223), .B2(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n257), .B1(new_n388), .B2(new_n259), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n263), .A2(G232), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(G190), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n390), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G200), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n342), .A2(new_n309), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT77), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n315), .A2(new_n297), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT77), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n342), .A2(new_n397), .A3(new_n309), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n341), .A2(new_n315), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n384), .A2(new_n391), .A3(new_n393), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT17), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n365), .A2(KEYINPUT16), .A3(new_n371), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT76), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n365), .A2(new_n375), .A3(new_n371), .A4(KEYINPUT16), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n401), .B1(new_n409), .B2(new_n374), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n410), .A2(KEYINPUT17), .A3(new_n393), .A4(new_n391), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n392), .A2(new_n288), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n290), .B1(new_n389), .B2(new_n390), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT78), .ZN(new_n416));
  AOI211_X1 g0216(.A(new_n416), .B(new_n401), .C1(new_n409), .C2(new_n374), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT78), .B1(new_n384), .B2(new_n402), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n297), .B1(new_n380), .B2(KEYINPUT16), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n408), .B2(new_n407), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n416), .B1(new_n423), .B2(new_n401), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n384), .A2(KEYINPUT78), .A3(new_n402), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(KEYINPUT18), .A3(new_n415), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n412), .B1(new_n421), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n263), .A2(G226), .ZN(new_n429));
  INV_X1    g0229(.A(G222), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT66), .B1(new_n330), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT66), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n329), .A2(new_n432), .A3(G222), .A4(new_n266), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G223), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n333), .B2(new_n335), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n329), .A2(new_n221), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n254), .B(new_n429), .C1(new_n438), .C2(new_n276), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n290), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n341), .A2(new_n298), .ZN(new_n441));
  NOR3_X1   g0241(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n442));
  INV_X1    g0242(.A(G150), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n442), .A2(new_n230), .B1(new_n300), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n297), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n396), .A2(G50), .A3(new_n309), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n315), .A2(new_n219), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  OR2_X1    g0248(.A1(new_n436), .A2(new_n437), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n259), .B1(new_n449), .B2(new_n434), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n450), .A2(new_n288), .A3(new_n254), .A4(new_n429), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n440), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT9), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n448), .A2(KEYINPUT70), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n448), .A2(KEYINPUT70), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n448), .A2(KEYINPUT70), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(new_n455), .A3(KEYINPUT9), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n450), .A2(G190), .A3(new_n254), .A4(new_n429), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n439), .A2(G200), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT10), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT10), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n461), .A2(new_n463), .A3(new_n466), .A4(new_n462), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n453), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n428), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n360), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n261), .A2(G1), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(G274), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G250), .B(new_n266), .C1(new_n269), .C2(new_n270), .ZN(new_n476));
  OAI211_X1 g0276(.A(G257), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G294), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n259), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n259), .B1(new_n472), .B2(new_n473), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G264), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT89), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n475), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n259), .A2(new_n479), .B1(new_n481), .B2(G264), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT89), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(G179), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(G169), .B1(new_n483), .B2(new_n475), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n275), .A2(G1), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n315), .A2(new_n297), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(new_n209), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n304), .A2(G107), .ZN(new_n496));
  XNOR2_X1  g0296(.A(new_n496), .B(KEYINPUT25), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n230), .B(G87), .C1(new_n269), .C2(new_n270), .ZN(new_n498));
  AND2_X1   g0298(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n499));
  NOR2_X1   g0299(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n329), .A2(new_n230), .A3(G87), .A4(new_n499), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n209), .A2(G20), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT23), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n504), .B(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n346), .A2(G116), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n502), .A2(new_n503), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  XNOR2_X1  g0309(.A(new_n508), .B(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n495), .B(new_n497), .C1(new_n510), .C2(new_n310), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n490), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT85), .B1(new_n332), .B2(new_n210), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n329), .A2(G257), .A3(new_n266), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT85), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n329), .A2(new_n515), .A3(G264), .A4(G1698), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n361), .A2(G303), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n513), .A2(new_n514), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n259), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n481), .A2(G270), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n474), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G283), .ZN(new_n523));
  INV_X1    g0323(.A(G97), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n523), .B(new_n230), .C1(G33), .C2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(G116), .ZN(new_n526));
  AOI221_X4 g0326(.A(KEYINPUT87), .B1(new_n526), .B2(G20), .C1(new_n296), .C2(new_n229), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT87), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(G20), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n528), .B1(new_n297), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n525), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT20), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(KEYINPUT20), .B(new_n525), .C1(new_n527), .C2(new_n530), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(G116), .B1(new_n275), .B2(G1), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n313), .A2(new_n297), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT86), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n308), .B2(G116), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n313), .A2(KEYINPUT86), .A3(new_n526), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n522), .A2(G179), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT21), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n290), .B1(new_n535), .B2(new_n541), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(new_n521), .ZN(new_n546));
  AND4_X1   g0346(.A1(new_n544), .A2(new_n542), .A3(G169), .A4(new_n521), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n512), .B(new_n543), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n329), .A2(new_n230), .A3(G68), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n272), .A2(new_n230), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n550), .B(KEYINPUT19), .C1(new_n203), .C2(G87), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n272), .A2(G20), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n549), .B(new_n551), .C1(KEYINPUT19), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n297), .ZN(new_n554));
  INV_X1    g0354(.A(new_n345), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n313), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n492), .A2(G87), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(G244), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT84), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n329), .A2(KEYINPUT84), .A3(G244), .A4(G1698), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G33), .A2(G116), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n330), .B2(new_n214), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n259), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT82), .B1(new_n261), .B2(G1), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT82), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n253), .A3(G45), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n276), .A2(G250), .A3(new_n568), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT83), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n216), .B1(new_n473), .B2(new_n569), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT83), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n573), .A2(new_n574), .A3(new_n276), .A4(new_n568), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n572), .A2(new_n575), .B1(G274), .B2(new_n473), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n567), .A2(G190), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n320), .B1(new_n567), .B2(new_n576), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n567), .A2(new_n288), .A3(new_n576), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n492), .A2(new_n345), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n554), .A2(new_n581), .A3(new_n556), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n567), .A2(new_n576), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n290), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n559), .A2(new_n579), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT79), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT4), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n587), .B(new_n588), .C1(new_n361), .C2(new_n222), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n329), .A2(G250), .B1(new_n587), .B2(new_n588), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n523), .C1(new_n590), .C2(new_n266), .ZN(new_n591));
  OAI211_X1 g0391(.A(G244), .B(new_n266), .C1(new_n269), .C2(new_n270), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n588), .B1(new_n592), .B2(new_n587), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n259), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n481), .A2(G257), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n474), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(G179), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(G250), .B1(new_n269), .B2(new_n270), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n587), .A2(new_n588), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n266), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n523), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n593), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(new_n589), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n596), .B1(new_n605), .B2(new_n259), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n598), .B1(new_n290), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n493), .A2(new_n524), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n379), .A2(G107), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n300), .A2(new_n221), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT6), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n524), .A2(new_n209), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n612), .B1(new_n613), .B2(new_n202), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n209), .A2(KEYINPUT6), .A3(G97), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n230), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n609), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n608), .B1(new_n618), .B2(new_n297), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT81), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n304), .A2(G97), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n608), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n209), .B1(new_n377), .B2(new_n378), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n625), .A2(new_n610), .A3(new_n616), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n622), .B(new_n624), .C1(new_n626), .C2(new_n310), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT81), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n607), .A2(new_n623), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT80), .B1(new_n606), .B2(new_n320), .ZN(new_n630));
  INV_X1    g0430(.A(new_n627), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n606), .A2(G190), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT80), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n600), .B1(new_n329), .B2(G244), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n601), .A2(new_n634), .A3(new_n602), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n276), .B1(new_n635), .B2(new_n604), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n633), .B(G200), .C1(new_n636), .C2(new_n596), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n630), .A2(new_n631), .A3(new_n632), .A4(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n503), .A2(new_n506), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n639), .A2(new_n509), .A3(new_n507), .A4(new_n502), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n508), .A2(KEYINPUT24), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n494), .B1(new_n642), .B2(new_n297), .ZN(new_n643));
  AOI21_X1  g0443(.A(G200), .B1(new_n485), .B2(new_n487), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n480), .A2(new_n482), .A3(new_n357), .A4(new_n474), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT90), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n486), .A2(KEYINPUT90), .A3(new_n357), .A4(new_n474), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n643), .B(new_n497), .C1(new_n644), .C2(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n586), .A2(new_n629), .A3(new_n638), .A4(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n542), .B1(G200), .B2(new_n521), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n522), .A2(G190), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR4_X1   g0455(.A1(new_n471), .A2(new_n548), .A3(new_n651), .A4(new_n655), .ZN(G372));
  XNOR2_X1  g0456(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n384), .A2(new_n402), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n657), .B1(new_n658), .B2(new_n415), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n658), .A2(new_n415), .A3(new_n657), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n355), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n318), .A2(new_n295), .B1(new_n663), .B2(new_n324), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n662), .B1(new_n664), .B2(new_n412), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n465), .A2(new_n467), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n453), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n585), .A2(new_n580), .A3(new_n582), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n543), .B1(new_n547), .B2(new_n546), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n490), .A2(new_n511), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n668), .B1(new_n671), .B2(new_n651), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n594), .A2(new_n597), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G169), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n631), .B1(new_n675), .B2(new_n598), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n586), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n584), .A2(G200), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n567), .A2(G190), .A3(new_n576), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n559), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n668), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n629), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n677), .B1(new_n682), .B2(new_n673), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n672), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n470), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n667), .A2(new_n685), .ZN(G369));
  INV_X1    g0486(.A(G13), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G20), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n253), .ZN(new_n689));
  XNOR2_X1  g0489(.A(KEYINPUT92), .B(KEYINPUT27), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n542), .A2(new_n695), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n669), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n696), .B1(new_n669), .B2(new_n655), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n670), .A2(new_n695), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n511), .B1(new_n490), .B2(new_n695), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(KEYINPUT93), .A3(new_n650), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT93), .B1(new_n703), .B2(new_n650), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n702), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT93), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n511), .A2(new_n695), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n512), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n650), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n709), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n695), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n669), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n713), .A2(new_n715), .A3(new_n704), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n670), .A2(new_n714), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n708), .A2(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n206), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G41), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G1), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n202), .A2(new_n215), .A3(new_n526), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n724), .A2(new_n725), .B1(new_n232), .B2(new_n723), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n586), .A2(new_n676), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT26), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n682), .A2(new_n673), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n714), .B1(new_n672), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT29), .ZN(new_n733));
  INV_X1    g0533(.A(new_n488), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n518), .A2(new_n259), .B1(G270), .B2(new_n481), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(new_n567), .A3(new_n576), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n734), .A2(KEYINPUT30), .A3(new_n606), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n584), .A2(KEYINPUT94), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT94), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n567), .A2(new_n740), .A3(new_n576), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n485), .A2(new_n487), .B1(new_n735), .B2(new_n474), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n742), .A2(new_n743), .A3(new_n288), .A4(new_n674), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n606), .A2(new_n485), .A3(G179), .A4(new_n487), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n745), .B1(new_n746), .B2(new_n736), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n738), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n695), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT31), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR4_X1   g0553(.A1(new_n651), .A2(new_n548), .A3(new_n655), .A4(new_n695), .ZN(new_n754));
  OAI21_X1  g0554(.A(G330), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT29), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n756), .B(new_n714), .C1(new_n672), .C2(new_n683), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n733), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n727), .B1(new_n758), .B2(G1), .ZN(G364));
  INV_X1    g0559(.A(new_n701), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n724), .B1(G45), .B2(new_n688), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n699), .A2(new_n700), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n760), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n762), .B1(new_n699), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n230), .A2(new_n288), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(G190), .A3(new_n320), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT95), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n769), .A2(KEYINPUT95), .A3(G190), .A4(new_n320), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT96), .Z(new_n775));
  NOR2_X1   g0575(.A1(new_n320), .A2(G190), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n769), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n775), .A2(G58), .B1(G68), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n357), .A2(new_n320), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n769), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n329), .B1(new_n781), .B2(new_n219), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n357), .A2(G179), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n230), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n769), .A2(new_n785), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n784), .A2(new_n524), .B1(new_n786), .B2(new_n221), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n230), .A2(G179), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n776), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n782), .B(new_n787), .C1(G107), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n780), .A2(new_n788), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n779), .B(new_n791), .C1(new_n215), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n788), .A2(new_n785), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G159), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT32), .ZN(new_n797));
  INV_X1    g0597(.A(G326), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n781), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n792), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G303), .A2(new_n800), .B1(new_n795), .B2(G329), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n801), .B(new_n361), .C1(new_n802), .C2(new_n786), .ZN(new_n803));
  INV_X1    g0603(.A(new_n784), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(G294), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n790), .A2(G283), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n774), .A2(G322), .ZN(new_n807));
  INV_X1    g0607(.A(G317), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(KEYINPUT33), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n808), .A2(KEYINPUT33), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n778), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n805), .A2(new_n806), .A3(new_n807), .A4(new_n811), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n793), .A2(new_n797), .B1(new_n799), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n229), .B1(G20), .B2(new_n290), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(G355), .A2(new_n329), .A3(new_n206), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n247), .A2(new_n261), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n721), .A2(new_n329), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(G45), .B2(new_n232), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n816), .B1(G116), .B2(new_n206), .C1(new_n817), .C2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n767), .A2(new_n814), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n768), .A2(new_n815), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n764), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT97), .ZN(G396));
  NAND2_X1  g0625(.A1(new_n349), .A2(new_n695), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT102), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n355), .A2(new_n359), .A3(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n829), .B(new_n714), .C1(new_n672), .C2(new_n683), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n684), .A2(new_n714), .ZN(new_n831));
  INV_X1    g0631(.A(new_n826), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n351), .A2(new_n352), .A3(new_n354), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n830), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n835), .A2(new_n755), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n755), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n836), .A2(new_n762), .A3(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n775), .A2(G143), .B1(G150), .B2(new_n778), .ZN(new_n839));
  INV_X1    g0639(.A(G137), .ZN(new_n840));
  INV_X1    g0640(.A(G159), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n839), .B1(new_n840), .B2(new_n781), .C1(new_n841), .C2(new_n786), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT34), .Z(new_n843));
  OAI22_X1  g0643(.A1(new_n792), .A2(new_n219), .B1(new_n789), .B2(new_n213), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n361), .B(new_n844), .C1(G58), .C2(new_n804), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n845), .B1(new_n846), .B2(new_n794), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT101), .Z(new_n848));
  NOR2_X1   g0648(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(G283), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n526), .A2(new_n786), .B1(new_n777), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT98), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n852), .B1(new_n524), .B2(new_n784), .C1(new_n209), .C2(new_n792), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(G294), .B2(new_n774), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n789), .A2(new_n215), .B1(new_n794), .B2(new_n802), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT99), .ZN(new_n856));
  INV_X1    g0656(.A(new_n781), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n329), .B1(new_n857), .B2(G303), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n854), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT100), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n814), .B1(new_n849), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n834), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n765), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n814), .A2(new_n765), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n221), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n861), .A2(new_n863), .A3(new_n761), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n838), .A2(new_n866), .ZN(G384));
  NOR2_X1   g0667(.A1(new_n317), .A2(new_n714), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n292), .A2(new_n294), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n286), .A2(G179), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT75), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n286), .A2(new_n252), .A3(G179), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n324), .B(new_n869), .C1(new_n874), .C2(new_n317), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n295), .A2(new_n868), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n651), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n878), .A2(new_n671), .A3(new_n654), .A4(new_n714), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n752), .A3(new_n751), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n877), .A2(new_n880), .A3(new_n834), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n693), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n417), .A2(new_n418), .B1(new_n415), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n403), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n403), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n413), .A2(new_n414), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT103), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n890), .B(new_n297), .C1(new_n380), .C2(KEYINPUT16), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT16), .B1(new_n365), .B2(new_n371), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT103), .B1(new_n892), .B2(new_n310), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n409), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n889), .B1(new_n894), .B2(new_n402), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n693), .B1(new_n894), .B2(new_n402), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n888), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n887), .B1(new_n897), .B2(new_n885), .ZN(new_n898));
  INV_X1    g0698(.A(new_n896), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n898), .B1(new_n428), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n898), .B(KEYINPUT38), .C1(new_n428), .C2(new_n899), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT40), .B1(new_n882), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n693), .B1(new_n424), .B2(new_n425), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n658), .A2(new_n415), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n403), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n887), .ZN(new_n911));
  INV_X1    g0711(.A(new_n657), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n410), .A2(new_n889), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n913), .A2(new_n659), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n907), .B1(new_n914), .B2(new_n412), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n412), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT18), .B1(new_n426), .B2(new_n415), .ZN(new_n918));
  AOI211_X1 g0718(.A(new_n420), .B(new_n889), .C1(new_n424), .C2(new_n425), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n899), .A2(new_n403), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT37), .B1(new_n921), .B2(new_n895), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n920), .A2(new_n896), .B1(new_n922), .B2(new_n887), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n916), .B1(new_n923), .B2(KEYINPUT38), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n924), .A2(new_n881), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n906), .A2(new_n927), .A3(new_n470), .A4(new_n880), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n905), .A2(new_n926), .A3(new_n700), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n748), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT31), .B1(new_n748), .B2(new_n695), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n700), .B1(new_n932), .B2(new_n879), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n470), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n928), .B1(new_n929), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n883), .B1(new_n417), .B2(new_n418), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(new_n403), .A3(new_n908), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n938), .A2(KEYINPUT37), .B1(new_n886), .B2(new_n884), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n937), .B1(new_n662), .B2(new_n917), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n901), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n903), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT39), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n902), .A2(KEYINPUT39), .A3(new_n903), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n319), .A2(new_n695), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n662), .A2(new_n883), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n663), .A2(new_n714), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n830), .A2(new_n949), .B1(new_n875), .B2(new_n876), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n948), .B1(new_n904), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n936), .B(new_n952), .Z(new_n953));
  INV_X1    g0753(.A(new_n757), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n629), .A2(new_n681), .A3(KEYINPUT26), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n673), .B1(new_n586), .B2(new_n676), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n629), .A2(new_n638), .ZN(new_n958));
  INV_X1    g0758(.A(new_n511), .ZN(new_n959));
  INV_X1    g0759(.A(new_n644), .ZN(new_n960));
  INV_X1    g0760(.A(new_n649), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n681), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n548), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n957), .A2(new_n964), .A3(new_n668), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n756), .B1(new_n965), .B2(new_n714), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n470), .B1(new_n954), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n667), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n953), .B(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n253), .B2(new_n688), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n614), .A2(new_n615), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n526), .B1(new_n971), .B2(KEYINPUT35), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n972), .B(new_n231), .C1(KEYINPUT35), .C2(new_n971), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT36), .ZN(new_n974));
  OAI21_X1  g0774(.A(G77), .B1(new_n224), .B2(new_n213), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n975), .A2(new_n232), .B1(G50), .B2(new_n213), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(G1), .A3(new_n687), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n970), .A2(new_n974), .A3(new_n977), .ZN(G367));
  NAND2_X1  g0778(.A1(new_n558), .A2(new_n695), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n668), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT104), .Z(new_n981));
  NAND3_X1  g0781(.A1(new_n586), .A2(KEYINPUT105), .A3(new_n979), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT105), .ZN(new_n983));
  INV_X1    g0783(.A(new_n979), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n983), .B1(new_n681), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n981), .A2(new_n982), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n767), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n786), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n804), .A2(G107), .B1(new_n989), .B2(G283), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n802), .B2(new_n781), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n329), .B(new_n991), .C1(G294), .C2(new_n778), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n775), .A2(G303), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G97), .A2(new_n790), .B1(new_n795), .B2(G317), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n800), .A2(G116), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT46), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n992), .A2(new_n993), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n784), .A2(new_n213), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G159), .B2(new_n778), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n840), .B2(new_n794), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n361), .B(new_n1000), .C1(G50), .C2(new_n989), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n857), .A2(G143), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G58), .A2(new_n800), .B1(new_n790), .B2(G77), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n774), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1005), .A2(new_n443), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n997), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT47), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n814), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n818), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n821), .B1(new_n206), .B2(new_n555), .C1(new_n242), .C2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n988), .A2(new_n761), .A3(new_n1009), .A4(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n253), .B1(new_n688), .B2(G45), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n676), .A2(new_n695), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n629), .A2(new_n638), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n631), .A2(new_n714), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n716), .A2(new_n717), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT45), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(KEYINPUT44), .B1(new_n719), .B2(new_n1018), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT44), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1018), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n718), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1021), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1026), .A2(new_n701), .A3(new_n707), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1021), .A2(new_n708), .A3(new_n1022), .A4(new_n1025), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n716), .A2(KEYINPUT108), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT108), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n713), .A2(new_n715), .A3(new_n1030), .A4(new_n704), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n669), .A2(new_n714), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n702), .B(new_n1032), .C1(new_n705), .C2(new_n706), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1029), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n701), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n760), .A2(new_n1029), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AND3_X1   g0837(.A1(new_n1037), .A2(new_n758), .A3(KEYINPUT109), .ZN(new_n1038));
  AOI21_X1  g0838(.A(KEYINPUT109), .B1(new_n1037), .B2(new_n758), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1027), .B(new_n1028), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n758), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n722), .B(KEYINPUT41), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1014), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT42), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n713), .A2(new_n715), .A3(new_n1045), .A4(new_n704), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(KEYINPUT106), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1046), .A2(KEYINPUT106), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1044), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1046), .A2(KEYINPUT106), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1051), .A2(KEYINPUT42), .A3(new_n1047), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n629), .B1(new_n1024), .B2(new_n512), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n714), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1050), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1050), .A2(new_n1052), .A3(new_n1056), .A4(new_n1054), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT107), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1059), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n708), .A2(new_n1024), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1065), .B(new_n1059), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1012), .B1(new_n1043), .B2(new_n1069), .ZN(G387));
  NOR2_X1   g0870(.A1(new_n792), .A2(new_n221), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n213), .A2(new_n786), .B1(new_n777), .B2(new_n341), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT110), .Z(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n219), .B2(new_n1005), .C1(new_n443), .C2(new_n794), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1071), .B(new_n1074), .C1(new_n345), .C2(new_n804), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n790), .A2(G97), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n857), .A2(G159), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1075), .A2(new_n329), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n775), .A2(G317), .B1(G311), .B2(new_n778), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n989), .A2(G303), .ZN(new_n1080));
  INV_X1    g0880(.A(G322), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1079), .B(new_n1080), .C1(new_n1081), .C2(new_n781), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1082), .A2(KEYINPUT48), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1082), .A2(KEYINPUT48), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT49), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n804), .A2(G283), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n800), .A2(G294), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1087), .B(new_n1088), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT49), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n361), .B1(new_n794), .B2(new_n798), .C1(new_n526), .C2(new_n789), .ZN(new_n1093));
  OAI211_X1 g0893(.A(KEYINPUT111), .B(new_n1078), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT111), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1093), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1078), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1094), .A2(new_n814), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n342), .A2(new_n219), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT50), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n213), .A2(new_n221), .ZN(new_n1102));
  NOR4_X1   g0902(.A1(new_n1101), .A2(G45), .A3(new_n1102), .A4(new_n725), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n818), .B1(new_n238), .B2(new_n261), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n329), .A2(new_n725), .A3(new_n206), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n206), .A2(G107), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n821), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1099), .A2(new_n761), .A3(new_n1108), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n707), .A2(new_n987), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1109), .A2(new_n1110), .B1(new_n1014), .B2(new_n1037), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n733), .A2(new_n755), .A3(new_n757), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n723), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1113), .B2(new_n1112), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1111), .A2(new_n1115), .ZN(G393));
  NOR2_X1   g0916(.A1(new_n792), .A2(new_n213), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n774), .A2(G159), .B1(G150), .B2(new_n857), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT51), .Z(new_n1119));
  NAND2_X1  g0919(.A1(new_n795), .A2(G143), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n361), .B1(new_n804), .B2(G77), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n989), .A2(new_n342), .B1(new_n790), .B2(G87), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1117), .B(new_n1123), .C1(G50), .C2(new_n778), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n774), .A2(G311), .B1(G317), .B2(new_n857), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT52), .Z(new_n1126));
  NAND2_X1  g0926(.A1(new_n778), .A2(G303), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n804), .A2(G116), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1126), .A2(new_n361), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n794), .A2(new_n1081), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n989), .A2(G294), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n792), .A2(new_n850), .B1(new_n789), .B2(new_n209), .ZN(new_n1132));
  NOR4_X1   g0932(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n814), .B1(new_n1124), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1024), .A2(new_n767), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n821), .B1(new_n524), .B2(new_n206), .C1(new_n250), .C2(new_n1010), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1134), .A2(new_n1135), .A3(new_n761), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n1013), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1139), .B1(new_n1144), .B2(new_n722), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(G390));
  AND3_X1   g0946(.A1(new_n902), .A2(KEYINPUT39), .A3(new_n903), .ZN(new_n1147));
  AOI21_X1  g0947(.A(KEYINPUT39), .B1(new_n941), .B2(new_n903), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1147), .A2(new_n1148), .B1(new_n946), .B2(new_n950), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n834), .B(new_n714), .C1(new_n672), .C2(new_n731), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n949), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n877), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n946), .B1(new_n941), .B2(new_n903), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n933), .A2(new_n834), .A3(new_n877), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1149), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AND4_X1   g0956(.A1(G330), .A2(new_n877), .A3(new_n880), .A4(new_n834), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n830), .A2(new_n949), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n877), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n946), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n944), .A2(new_n945), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1157), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n967), .A2(new_n667), .A3(new_n934), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n877), .B1(new_n933), .B2(new_n834), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1158), .B1(new_n1157), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1151), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n755), .A2(new_n862), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1167), .B(new_n1155), .C1(new_n1168), .C2(new_n877), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1164), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1156), .A2(new_n1163), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n722), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT112), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1156), .A2(new_n1163), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1170), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1171), .A2(KEYINPUT112), .A3(new_n722), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1174), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1156), .A2(new_n1163), .A3(new_n1014), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n765), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n762), .B1(new_n341), .B2(new_n864), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT113), .Z(new_n1183));
  AOI22_X1  g0983(.A1(new_n774), .A2(G116), .B1(G77), .B2(new_n804), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT114), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n795), .A2(G294), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n786), .A2(new_n524), .ZN(new_n1187));
  NOR4_X1   g0987(.A1(new_n1185), .A2(new_n329), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G87), .A2(new_n800), .B1(new_n790), .B2(G68), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n850), .C2(new_n781), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n777), .A2(new_n209), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n792), .A2(KEYINPUT53), .A3(new_n443), .ZN(new_n1192));
  OAI21_X1  g0992(.A(KEYINPUT53), .B1(new_n792), .B2(new_n443), .ZN(new_n1193));
  INV_X1    g0993(.A(G128), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(KEYINPUT54), .B(G143), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1193), .B1(new_n1194), .B2(new_n781), .C1(new_n786), .C2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G137), .B2(new_n778), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n361), .B1(new_n795), .B2(G125), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n841), .B2(new_n784), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G132), .B2(new_n774), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1197), .B(new_n1200), .C1(new_n219), .C2(new_n789), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n1190), .A2(new_n1191), .B1(new_n1192), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1183), .B1(new_n1202), .B2(new_n814), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT115), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1181), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1179), .A2(new_n1180), .A3(new_n1205), .ZN(G378));
  NAND3_X1  g1006(.A1(new_n906), .A2(new_n927), .A3(G330), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n456), .A2(new_n457), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n883), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT55), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n468), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n468), .A2(new_n1212), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1211), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n468), .A2(new_n1212), .ZN(new_n1216));
  AOI211_X1 g1016(.A(KEYINPUT55), .B(new_n453), .C1(new_n465), .C2(new_n467), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1211), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1209), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1213), .A2(new_n1214), .A3(new_n1211), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1218), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n1222), .A3(new_n1208), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n947), .A2(new_n1224), .A3(new_n951), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1224), .B1(new_n947), .B2(new_n951), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1207), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1224), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n952), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n947), .A2(new_n1224), .A3(new_n951), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n929), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1227), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1164), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1171), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT57), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1232), .A2(new_n1234), .A3(KEYINPUT57), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n722), .A3(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n789), .A2(new_n224), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT116), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n209), .B2(new_n1005), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1242), .A2(new_n329), .A3(new_n1071), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n345), .A2(new_n989), .B1(new_n795), .B2(G283), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n526), .B2(new_n781), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1245), .A2(G41), .A3(new_n998), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1243), .B(new_n1246), .C1(new_n524), .C2(new_n777), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT58), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n219), .B1(new_n269), .B2(G41), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n846), .A2(new_n777), .B1(new_n786), .B2(new_n840), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT117), .Z(new_n1251));
  OAI221_X1 g1051(.A(new_n1251), .B1(new_n443), .B2(new_n784), .C1(new_n792), .C2(new_n1195), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(G125), .B2(new_n857), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1194), .B2(new_n1005), .ZN(new_n1254));
  AOI21_X1  g1054(.A(G41), .B1(new_n1254), .B2(KEYINPUT59), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G33), .B1(new_n795), .B2(G124), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1255), .B(new_n1256), .C1(new_n841), .C2(new_n789), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1254), .A2(KEYINPUT59), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1248), .B(new_n1249), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT118), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n814), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n864), .A2(new_n219), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1220), .A2(new_n765), .A3(new_n1223), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1261), .A2(new_n761), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(KEYINPUT120), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1232), .A2(new_n1014), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1239), .A2(new_n1267), .ZN(G375));
  OAI22_X1  g1068(.A1(new_n555), .A2(new_n784), .B1(new_n526), .B2(new_n777), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n361), .B1(new_n1005), .B2(new_n850), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1269), .B(new_n1270), .C1(G107), .C2(new_n989), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n800), .A2(G97), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n857), .A2(G294), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(G77), .A2(new_n790), .B1(new_n795), .B2(G303), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1241), .B1(new_n1194), .B2(new_n794), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(new_n361), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n784), .A2(new_n219), .B1(new_n786), .B2(new_n443), .ZN(new_n1278));
  XOR2_X1   g1078(.A(new_n1278), .B(KEYINPUT121), .Z(new_n1279));
  OAI211_X1 g1079(.A(new_n1277), .B(new_n1279), .C1(new_n841), .C2(new_n792), .ZN(new_n1280));
  XOR2_X1   g1080(.A(new_n1280), .B(KEYINPUT122), .Z(new_n1281));
  NAND2_X1  g1081(.A1(new_n775), .A2(G137), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1281), .B(new_n1282), .C1(new_n846), .C2(new_n781), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n777), .A2(new_n1195), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1275), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n814), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1286), .B(new_n761), .C1(new_n766), .C2(new_n877), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n213), .B2(new_n864), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1288), .B1(new_n1289), .B2(new_n1014), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1042), .B1(new_n1289), .B2(new_n1233), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1290), .B1(new_n1291), .B2(new_n1170), .ZN(G381));
  NOR2_X1   g1092(.A1(G375), .A2(G378), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(G381), .A2(G384), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1145), .B(new_n1012), .C1(new_n1043), .C2(new_n1069), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(G393), .A2(G396), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1293), .A2(new_n1294), .A3(new_n1296), .A4(new_n1297), .ZN(G407));
  NAND2_X1  g1098(.A1(new_n694), .A2(G213), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(G375), .A2(G378), .A3(new_n1299), .ZN(new_n1300));
  OR2_X1    g1100(.A1(new_n1300), .A2(KEYINPUT123), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(KEYINPUT123), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1301), .A2(G213), .A3(G407), .A4(new_n1302), .ZN(G409));
  INV_X1    g1103(.A(new_n1299), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT124), .B1(new_n1289), .B2(new_n1233), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(KEYINPUT60), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT60), .ZN(new_n1307));
  OAI211_X1 g1107(.A(KEYINPUT124), .B(new_n1307), .C1(new_n1289), .C2(new_n1233), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1306), .A2(new_n722), .A3(new_n1176), .A4(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(G384), .B1(new_n1309), .B2(new_n1290), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1309), .A2(G384), .A3(new_n1290), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(G378), .A2(new_n1239), .A3(new_n1267), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1042), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1266), .B(new_n1264), .C1(new_n1235), .C2(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1316), .A2(new_n1180), .A3(new_n1179), .A4(new_n1205), .ZN(new_n1317));
  AOI211_X1 g1117(.A(new_n1304), .B(new_n1313), .C1(new_n1314), .C2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(KEYINPUT63), .B1(new_n1318), .B2(KEYINPUT125), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT61), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G387), .A2(G390), .ZN(new_n1321));
  INV_X1    g1121(.A(G396), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1322), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1297), .A2(new_n1323), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1321), .A2(new_n1324), .A3(new_n1295), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1324), .B1(new_n1321), .B2(new_n1295), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1320), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1312), .ZN(new_n1328));
  OAI211_X1 g1128(.A(G2897), .B(new_n1304), .C1(new_n1328), .C2(new_n1310), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1304), .A2(G2897), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1311), .A2(new_n1312), .A3(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1314), .A2(new_n1317), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1299), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1327), .B1(new_n1333), .B2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT125), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT63), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n1337), .B(new_n1338), .C1(new_n1335), .C2(new_n1313), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1319), .A2(new_n1336), .A3(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1304), .B1(new_n1314), .B2(new_n1317), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT62), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1313), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1341), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  XOR2_X1   g1144(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1345));
  OAI21_X1  g1145(.A(new_n1345), .B1(new_n1341), .B2(new_n1332), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1342), .B1(new_n1341), .B2(new_n1343), .ZN(new_n1347));
  NOR3_X1   g1147(.A1(new_n1344), .A2(new_n1346), .A3(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1326), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1321), .A2(new_n1295), .A3(new_n1324), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1340), .B1(new_n1348), .B2(new_n1351), .ZN(G405));
  INV_X1    g1152(.A(G375), .ZN(new_n1353));
  OR2_X1    g1153(.A1(new_n1353), .A2(G378), .ZN(new_n1354));
  OAI211_X1 g1154(.A(new_n1354), .B(new_n1314), .C1(KEYINPUT127), .C2(new_n1313), .ZN(new_n1355));
  OAI211_X1 g1155(.A(KEYINPUT127), .B(new_n1313), .C1(new_n1325), .C2(new_n1326), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1313), .A2(KEYINPUT127), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1349), .A2(new_n1350), .A3(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1356), .A2(new_n1358), .ZN(new_n1359));
  XNOR2_X1  g1159(.A(new_n1355), .B(new_n1359), .ZN(G402));
endmodule


