//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n590, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT66), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT68), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n459), .A2(G2105), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n463), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n464), .A2(G136), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n475), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  AND2_X1   g055(.A1(new_n460), .A2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n473), .ZN(new_n482));
  INV_X1    g057(.A(G138), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT4), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n464), .A2(new_n485), .A3(G138), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G114), .C2(new_n473), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n474), .A2(G126), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(G164));
  NAND2_X1  g066(.A1(G75), .A2(G543), .ZN(new_n492));
  INV_X1    g067(.A(G543), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT5), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G62), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n492), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G651), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  XNOR2_X1  g076(.A(new_n500), .B(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n494), .A2(new_n496), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G88), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n504), .A2(new_n506), .A3(G543), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n512), .B(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n502), .A2(new_n509), .A3(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  INV_X1    g091(.A(G51), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n510), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT5), .B(G543), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n520), .A2(new_n522), .A3(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT7), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n526), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n523), .A2(KEYINPUT71), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(KEYINPUT71), .B1(new_n523), .B2(new_n528), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n519), .B(new_n521), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(G168));
  XNOR2_X1  g107(.A(KEYINPUT73), .B(G52), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n510), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n520), .A2(new_n522), .A3(G90), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n520), .B2(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(KEYINPUT72), .B1(new_n538), .B2(new_n503), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n494), .A2(new_n496), .A3(G64), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(new_n536), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n541), .A2(new_n542), .A3(G651), .ZN(new_n543));
  AOI211_X1 g118(.A(new_n534), .B(new_n535), .C1(new_n539), .C2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n508), .A2(G81), .B1(new_n511), .B2(G43), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OAI21_X1  g121(.A(KEYINPUT74), .B1(new_n546), .B2(new_n503), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n497), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n550), .A2(new_n551), .A3(G651), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n545), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G860), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n553), .A2(new_n554), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  NAND4_X1  g135(.A1(new_n504), .A2(new_n506), .A3(G53), .A4(G543), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n562), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT9), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n565), .A2(new_n566), .B1(G91), .B2(new_n508), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n495), .A2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n493), .A2(KEYINPUT5), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT76), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n494), .A2(new_n496), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(G65), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  AND3_X1   g149(.A1(new_n573), .A2(KEYINPUT77), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(KEYINPUT77), .B1(new_n573), .B2(new_n574), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(KEYINPUT78), .B1(new_n577), .B2(G651), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n494), .A2(new_n496), .A3(new_n571), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n571), .B1(new_n494), .B2(new_n496), .ZN(new_n581));
  INV_X1    g156(.A(G65), .ZN(new_n582));
  NOR3_X1   g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n574), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n579), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n573), .A2(KEYINPUT77), .A3(new_n574), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT78), .A4(G651), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n567), .B1(new_n578), .B2(new_n588), .ZN(G299));
  AOI21_X1  g164(.A(new_n535), .B1(new_n539), .B2(new_n543), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(new_n510), .B2(new_n533), .ZN(G301));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n531), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G89), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n528), .B1(new_n507), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT71), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n523), .A2(KEYINPUT71), .A3(new_n528), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n599), .A2(KEYINPUT79), .A3(new_n519), .A4(new_n521), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n593), .A2(new_n600), .ZN(G286));
  NAND2_X1  g176(.A1(new_n508), .A2(G87), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n511), .A2(G49), .ZN(new_n603));
  OAI21_X1  g178(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(G288));
  AOI22_X1  g180(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(new_n503), .ZN(new_n607));
  INV_X1    g182(.A(G86), .ZN(new_n608));
  INV_X1    g183(.A(G48), .ZN(new_n609));
  OAI22_X1  g184(.A1(new_n507), .A2(new_n608), .B1(new_n510), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(G305));
  AOI22_X1  g187(.A1(new_n508), .A2(G85), .B1(new_n511), .B2(G47), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n503), .B2(new_n614), .ZN(G290));
  NAND2_X1  g190(.A1(G301), .A2(G868), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n507), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n520), .A2(new_n522), .A3(KEYINPUT10), .A4(G92), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n570), .A2(G66), .A3(new_n572), .ZN(new_n622));
  NAND2_X1  g197(.A1(G79), .A2(G543), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n503), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n510), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n522), .A2(KEYINPUT80), .A3(G543), .ZN(new_n627));
  AND3_X1   g202(.A1(new_n626), .A2(new_n627), .A3(G54), .ZN(new_n628));
  NOR3_X1   g203(.A1(new_n621), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n616), .B1(G868), .B2(new_n629), .ZN(G284));
  OAI21_X1  g205(.A(new_n616), .B1(G868), .B2(new_n629), .ZN(G321));
  NAND2_X1  g206(.A1(G286), .A2(G868), .ZN(new_n632));
  INV_X1    g207(.A(new_n567), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n585), .A2(G651), .A3(new_n586), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT78), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n633), .B1(new_n636), .B2(new_n587), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n632), .B1(new_n637), .B2(G868), .ZN(G297));
  OAI21_X1  g213(.A(new_n632), .B1(new_n637), .B2(G868), .ZN(G280));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n629), .B1(new_n640), .B2(G860), .ZN(G148));
  INV_X1    g216(.A(G868), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n553), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n629), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n644), .A2(G559), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n643), .B1(new_n645), .B2(new_n642), .ZN(G323));
  XNOR2_X1  g221(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g222(.A1(new_n481), .A2(new_n465), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT13), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G2100), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT81), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n474), .A2(G123), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT83), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n473), .A2(G111), .ZN(new_n659));
  AOI22_X1  g234(.A1(new_n464), .A2(G135), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n474), .A2(KEYINPUT83), .A3(G123), .ZN(new_n661));
  AND3_X1   g236(.A1(new_n656), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2096), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n651), .A2(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT82), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n653), .A2(new_n663), .A3(new_n665), .ZN(G156));
  XNOR2_X1  g241(.A(G2427), .B(G2438), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2430), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT15), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n669), .A2(G2435), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(G2435), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(KEYINPUT14), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2451), .B(G2454), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT16), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2443), .B(G2446), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1341), .B(G1348), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT84), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n681), .B(G14), .C1(new_n679), .C2(new_n677), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G401));
  XOR2_X1   g258(.A(G2084), .B(G2090), .Z(new_n684));
  XNOR2_X1  g259(.A(G2072), .B(G2078), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT85), .Z(new_n686));
  XOR2_X1   g261(.A(G2067), .B(G2678), .Z(new_n687));
  AOI21_X1  g262(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n685), .B(KEYINPUT17), .Z(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n687), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(new_n685), .A3(new_n684), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT18), .Z(new_n693));
  NAND3_X1  g268(.A1(new_n689), .A2(new_n687), .A3(new_n684), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n690), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G2096), .B(G2100), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G227));
  XNOR2_X1  g272(.A(G1971), .B(G1976), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n698), .B(new_n699), .Z(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1956), .B(G2474), .Z(new_n702));
  XOR2_X1   g277(.A(G1961), .B(G1966), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT20), .Z(new_n706));
  NOR2_X1   g281(.A1(new_n702), .A2(new_n703), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n700), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT87), .Z(new_n709));
  INV_X1    g284(.A(new_n707), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n701), .A2(new_n710), .A3(new_n704), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n706), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT88), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n714));
  XNOR2_X1  g289(.A(G1981), .B(G1986), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n713), .B(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(G1991), .B(G1996), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(G229));
  NAND2_X1  g294(.A1(new_n474), .A2(G119), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n464), .A2(G131), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n473), .A2(G107), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n720), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT89), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT90), .ZN(new_n726));
  MUX2_X1   g301(.A(G25), .B(new_n726), .S(G29), .Z(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT91), .Z(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT35), .B(G1991), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  MUX2_X1   g306(.A(G24), .B(G290), .S(G16), .Z(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(G1986), .Z(new_n733));
  NAND3_X1  g308(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G22), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G166), .B2(new_n735), .ZN(new_n737));
  INV_X1    g312(.A(G1971), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G16), .A2(G23), .ZN(new_n740));
  INV_X1    g315(.A(G288), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT33), .B(G1976), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(G6), .A2(G16), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n611), .B2(G16), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT32), .B(G1981), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n739), .A2(new_n744), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT34), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n734), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT92), .B(KEYINPUT36), .Z(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n752), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n734), .A2(new_n750), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT28), .ZN(new_n757));
  INV_X1    g332(.A(G26), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(G29), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(G29), .ZN(new_n760));
  OAI21_X1  g335(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n761));
  INV_X1    g336(.A(G116), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(G2105), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT93), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n474), .A2(G128), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n464), .A2(G140), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n760), .B1(new_n767), .B2(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n759), .B1(new_n768), .B2(new_n757), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(G2067), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n662), .A2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT97), .ZN(new_n772));
  NOR2_X1   g347(.A1(G27), .A2(G29), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G164), .B2(G29), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G2078), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n769), .A2(G2067), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n770), .A2(new_n772), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G29), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G33), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT25), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n464), .A2(G139), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n481), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n781), .B(new_n782), .C1(new_n783), .C2(new_n473), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT94), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n779), .B1(new_n786), .B2(new_n778), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n787), .A2(G2072), .ZN(new_n788));
  OR2_X1    g363(.A1(G29), .A2(G32), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n464), .A2(G141), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n474), .A2(G129), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n465), .A2(G105), .ZN(new_n792));
  NAND3_X1  g367(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT26), .Z(new_n794));
  NAND4_X1  g369(.A1(new_n790), .A2(new_n791), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n789), .B1(new_n795), .B2(new_n778), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT27), .B(G1996), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT95), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT30), .B(G28), .Z(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(G29), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n774), .A2(G2078), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n777), .A2(new_n788), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(G168), .A2(new_n735), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n735), .B2(G21), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT96), .B(G1966), .Z(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OAI22_X1  g382(.A1(new_n787), .A2(G2072), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n807), .B2(new_n805), .ZN(new_n809));
  NAND2_X1  g384(.A1(G171), .A2(G16), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G5), .B2(G16), .ZN(new_n811));
  INV_X1    g386(.A(G1961), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n735), .A2(KEYINPUT23), .A3(G20), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT23), .ZN(new_n815));
  INV_X1    g390(.A(G20), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(G16), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n814), .B(new_n817), .C1(new_n637), .C2(new_n735), .ZN(new_n818));
  INV_X1    g393(.A(G1956), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n803), .A2(new_n809), .A3(new_n813), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n778), .A2(G35), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G162), .B2(new_n778), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT29), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(G2090), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n735), .A2(G4), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n629), .B2(new_n735), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(G1348), .Z(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT31), .B(G11), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n824), .A2(G2090), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT99), .Z(new_n832));
  MUX2_X1   g407(.A(G19), .B(new_n553), .S(G16), .Z(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(G1341), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR4_X1   g410(.A1(new_n821), .A2(new_n825), .A3(new_n830), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n811), .A2(new_n812), .ZN(new_n837));
  OR2_X1    g412(.A1(KEYINPUT24), .A2(G34), .ZN(new_n838));
  NAND2_X1  g413(.A1(KEYINPUT24), .A2(G34), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n838), .A2(new_n778), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G160), .B2(new_n778), .ZN(new_n841));
  OAI221_X1 g416(.A(new_n837), .B1(G2084), .B2(new_n841), .C1(new_n796), .C2(new_n797), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT98), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(G2084), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n836), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT100), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n756), .A2(new_n846), .ZN(G311));
  NAND2_X1  g422(.A1(new_n756), .A2(new_n846), .ZN(G150));
  AOI22_X1  g423(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n849), .A2(new_n503), .ZN(new_n850));
  INV_X1    g425(.A(G93), .ZN(new_n851));
  XNOR2_X1  g426(.A(KEYINPUT101), .B(G55), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n507), .A2(new_n851), .B1(new_n510), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n854), .A2(new_n554), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n629), .A2(G559), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT38), .Z(new_n858));
  OR2_X1    g433(.A1(new_n510), .A2(new_n852), .ZN(new_n859));
  OAI221_X1 g434(.A(new_n859), .B1(new_n851), .B2(new_n507), .C1(new_n503), .C2(new_n849), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n860), .A2(new_n545), .A3(new_n547), .A4(new_n552), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n553), .A2(new_n854), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n858), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT102), .Z(new_n867));
  OAI21_X1  g442(.A(new_n554), .B1(new_n865), .B2(KEYINPUT39), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n856), .B1(new_n867), .B2(new_n868), .ZN(G145));
  AOI22_X1  g444(.A1(new_n484), .A2(new_n486), .B1(G126), .B2(new_n474), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n489), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n795), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n767), .ZN(new_n873));
  MUX2_X1   g448(.A(new_n786), .B(new_n784), .S(new_n873), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n464), .A2(G142), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n473), .A2(G118), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(G130), .B2(new_n474), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(new_n649), .Z(new_n880));
  XNOR2_X1  g455(.A(new_n874), .B(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(G162), .B(new_n471), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n662), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n725), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n881), .A2(new_n884), .ZN(new_n886));
  NOR3_X1   g461(.A1(new_n885), .A2(new_n886), .A3(G37), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(G395));
  NAND2_X1  g464(.A1(new_n860), .A2(new_n642), .ZN(new_n890));
  NAND2_X1  g465(.A1(G299), .A2(new_n629), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n637), .A2(new_n644), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n636), .A2(new_n587), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n644), .B1(new_n895), .B2(new_n567), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT103), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n645), .B(new_n863), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI211_X1 g475(.A(new_n633), .B(new_n629), .C1(new_n636), .C2(new_n587), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n896), .A2(new_n901), .A3(KEYINPUT41), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n637), .A2(new_n892), .A3(new_n644), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n896), .A2(new_n901), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n904), .B2(new_n892), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n902), .B1(new_n905), .B2(KEYINPUT41), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n900), .B1(new_n906), .B2(new_n899), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT42), .ZN(new_n908));
  XNOR2_X1  g483(.A(G303), .B(new_n611), .ZN(new_n909));
  XNOR2_X1  g484(.A(G290), .B(G288), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n908), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n890), .B1(new_n912), .B2(new_n642), .ZN(G295));
  OAI21_X1  g488(.A(new_n890), .B1(new_n912), .B2(new_n642), .ZN(G331));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n915));
  INV_X1    g490(.A(new_n911), .ZN(new_n916));
  INV_X1    g491(.A(new_n863), .ZN(new_n917));
  NOR2_X1   g492(.A1(G171), .A2(new_n531), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n919));
  AOI22_X1  g494(.A1(G286), .A2(G171), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT105), .B1(G171), .B2(new_n531), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(G301), .B1(new_n593), .B2(new_n600), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n919), .B1(G301), .B2(G168), .ZN(new_n924));
  NOR3_X1   g499(.A1(G171), .A2(new_n531), .A3(KEYINPUT105), .ZN(new_n925));
  NOR4_X1   g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .A4(new_n863), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n894), .A2(KEYINPUT41), .A3(new_n897), .ZN(new_n928));
  INV_X1    g503(.A(new_n902), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(G286), .A2(G171), .ZN(new_n931));
  INV_X1    g506(.A(new_n925), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n921), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n863), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n920), .A2(new_n917), .A3(new_n921), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n905), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n916), .B1(new_n930), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G37), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n936), .B(KEYINPUT41), .C1(new_n896), .C2(new_n901), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n936), .A2(KEYINPUT41), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n940), .B(new_n911), .C1(new_n941), .C2(new_n905), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n938), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n930), .A2(new_n937), .A3(new_n916), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT106), .B1(new_n944), .B2(G37), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n927), .A2(new_n898), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n911), .B(new_n946), .C1(new_n906), .C2(new_n927), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(new_n948), .A3(new_n939), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n938), .A3(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n951));
  OAI221_X1 g526(.A(KEYINPUT44), .B1(new_n915), .B2(new_n943), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n951), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n938), .A2(new_n942), .A3(new_n939), .A4(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT107), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n950), .A2(new_n951), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT108), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n960));
  AOI211_X1 g535(.A(new_n960), .B(KEYINPUT44), .C1(new_n955), .C2(new_n956), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n952), .B1(new_n959), .B2(new_n961), .ZN(G397));
  INV_X1    g537(.A(KEYINPUT117), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n964));
  NOR3_X1   g539(.A1(G164), .A2(new_n964), .A3(G1384), .ZN(new_n965));
  AOI21_X1  g540(.A(G1384), .B1(new_n870), .B2(new_n489), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(KEYINPUT45), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT110), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n466), .A2(G40), .A3(new_n470), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n964), .B1(G164), .B2(G1384), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT56), .B(G2072), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n968), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n966), .ZN(new_n976));
  XNOR2_X1  g551(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n966), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n969), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n975), .B1(G1956), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(G299), .B(KEYINPUT57), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n963), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n969), .B1(new_n967), .B2(KEYINPUT110), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n966), .A2(KEYINPUT45), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n972), .B1(new_n971), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n989), .A2(new_n974), .B1(new_n819), .B2(new_n981), .ZN(new_n990));
  INV_X1    g565(.A(new_n984), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(KEYINPUT117), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n983), .A2(new_n984), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n985), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT61), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n989), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n871), .A2(new_n999), .A3(new_n969), .ZN(new_n1000));
  XOR2_X1   g575(.A(KEYINPUT58), .B(G1341), .Z(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n553), .B1(new_n998), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT59), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1000), .A2(G2067), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n977), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n871), .A2(new_n999), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n969), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n966), .A2(new_n979), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1006), .B(new_n1008), .C1(new_n1013), .C2(G1348), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n970), .B1(new_n966), .B2(new_n1009), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1348), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT118), .B1(new_n1017), .B2(new_n1007), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n644), .B1(new_n1019), .B2(KEYINPUT60), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT60), .ZN(new_n1021));
  AOI211_X1 g596(.A(new_n1021), .B(new_n629), .C1(new_n1014), .C2(new_n1018), .ZN(new_n1022));
  OAI22_X1  g597(.A1(new_n1020), .A2(new_n1022), .B1(KEYINPUT60), .B2(new_n1019), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n990), .A2(new_n991), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(new_n993), .A3(KEYINPUT61), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n996), .A2(new_n1005), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n993), .B1(new_n644), .B2(new_n1019), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(new_n985), .A3(new_n992), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n971), .A2(new_n987), .A3(new_n969), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n807), .ZN(new_n1032));
  INV_X1    g607(.A(G2084), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1015), .A2(new_n1016), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1030), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n531), .A2(G8), .ZN(new_n1036));
  XOR2_X1   g611(.A(new_n1036), .B(KEYINPUT119), .Z(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT120), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1013), .A2(new_n1033), .B1(new_n1031), .B2(new_n807), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1040), .B(new_n1037), .C1(new_n1041), .C2(new_n1030), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1042), .A3(KEYINPUT51), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1041), .A2(new_n1037), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT120), .B(new_n1045), .C1(new_n1035), .C2(new_n1038), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1961), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1048));
  INV_X1    g623(.A(G2078), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n968), .A2(new_n973), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(KEYINPUT53), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1031), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1052), .A2(new_n1053), .A3(G301), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n1060));
  AOI211_X1 g635(.A(new_n1048), .B(new_n1055), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(G301), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(KEYINPUT121), .A3(G171), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT122), .B1(new_n1063), .B2(G171), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1059), .A2(new_n1062), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1063), .A2(G171), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1061), .A2(G301), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT54), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1047), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G305), .A2(G1981), .ZN(new_n1071));
  OR3_X1    g646(.A1(new_n607), .A2(new_n610), .A3(G1981), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(KEYINPUT114), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n1074));
  NAND3_X1  g649(.A1(G305), .A2(new_n1074), .A3(G1981), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1076), .B1(new_n1077), .B2(KEYINPUT49), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1000), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(new_n1030), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1077), .A2(KEYINPUT49), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1073), .A2(new_n1081), .A3(new_n1075), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1078), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT113), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n741), .A2(G1976), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1000), .A2(new_n1085), .A3(G8), .A4(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1976), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1000), .A2(G8), .A3(new_n1088), .A4(G288), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1087), .B1(new_n1090), .B2(new_n1089), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1083), .B(new_n1084), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1087), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1091), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1084), .B1(new_n1099), .B2(new_n1083), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT112), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1104), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT112), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n1107), .A3(new_n1102), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1971), .B1(new_n968), .B2(new_n973), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1011), .A2(G2090), .A3(new_n1012), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1109), .B(G8), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n981), .A2(G2090), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n738), .B1(new_n986), .B2(new_n988), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1030), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1106), .A2(new_n1102), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1112), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1101), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1029), .A2(new_n1070), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1043), .A2(new_n1120), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1118), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT123), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n1047), .A2(new_n1120), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1118), .A2(new_n1121), .A3(new_n1122), .A4(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1112), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1099), .A2(new_n1083), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  OAI221_X1 g707(.A(new_n1112), .B1(new_n1115), .B2(new_n1116), .C1(new_n1095), .C2(new_n1100), .ZN(new_n1133));
  INV_X1    g708(.A(G286), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1035), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1132), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(G8), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1116), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1132), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1135), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1139), .A2(new_n1112), .A3(new_n1130), .A4(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1083), .A2(new_n1088), .A3(new_n741), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1072), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1136), .A2(new_n1141), .B1(new_n1080), .B2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1119), .A2(new_n1128), .A3(new_n1131), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(G2067), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n767), .B(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(G1996), .B2(new_n795), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n971), .A2(new_n970), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n725), .B(new_n729), .Z(new_n1153));
  NAND2_X1  g728(.A1(new_n1150), .A2(new_n997), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT109), .ZN(new_n1155));
  OAI221_X1 g730(.A(new_n1152), .B1(new_n1151), .B2(new_n1153), .C1(new_n1155), .C2(new_n795), .ZN(new_n1156));
  XNOR2_X1  g731(.A(G290), .B(G1986), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1156), .B1(new_n1150), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1145), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1152), .B1(new_n1155), .B2(new_n795), .ZN(new_n1160));
  OR3_X1    g735(.A1(new_n1160), .A2(new_n729), .A3(new_n726), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n767), .A2(G2067), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1151), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1150), .B1(new_n795), .B2(new_n1148), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1155), .A2(KEYINPUT46), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1155), .A2(KEYINPUT46), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(KEYINPUT124), .B(KEYINPUT47), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1167), .B(new_n1168), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1151), .A2(G1986), .A3(G290), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT127), .ZN(new_n1171));
  XOR2_X1   g746(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1172));
  XNOR2_X1  g747(.A(new_n1171), .B(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1156), .B(KEYINPUT125), .Z(new_n1174));
  AOI211_X1 g749(.A(new_n1163), .B(new_n1169), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1159), .A2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g751(.A(G229), .ZN(new_n1178));
  NAND2_X1  g752(.A1(new_n957), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g753(.A(G319), .ZN(new_n1180));
  NOR2_X1   g754(.A1(G227), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g755(.A1(new_n682), .A2(new_n1181), .ZN(new_n1182));
  NOR3_X1   g756(.A1(new_n1179), .A2(new_n887), .A3(new_n1182), .ZN(G308));
  NOR2_X1   g757(.A1(new_n887), .A2(new_n1182), .ZN(new_n1184));
  NAND3_X1  g758(.A1(new_n1184), .A2(new_n1178), .A3(new_n957), .ZN(G225));
endmodule


