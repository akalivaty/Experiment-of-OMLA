//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT31), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT2), .B(G113), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G116), .B(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  XOR2_X1   g006(.A(G116), .B(G119), .Z(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(new_n189), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT1), .B1(new_n196), .B2(G146), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(G146), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  OAI211_X1 g014(.A(G128), .B(new_n197), .C1(new_n198), .C2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n196), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n202), .B(new_n203), .C1(KEYINPUT1), .C2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G134), .ZN(new_n209));
  OAI21_X1  g023(.A(G131), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n201), .A2(new_n205), .A3(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(KEYINPUT11), .A3(G134), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n206), .A2(G137), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT11), .B1(new_n208), .B2(G134), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT11), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(new_n206), .B2(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT67), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT68), .B(G131), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n214), .A2(new_n217), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n211), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n212), .B(new_n213), .C1(new_n215), .C2(new_n216), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n219), .A2(KEYINPUT67), .ZN(new_n225));
  OAI21_X1  g039(.A(G131), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n226), .A2(new_n222), .ZN(new_n227));
  XNOR2_X1  g041(.A(G143), .B(G146), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT0), .A3(G128), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT0), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n202), .A2(new_n203), .B1(new_n230), .B2(new_n204), .ZN(new_n231));
  AND3_X1   g045(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n231), .A2(KEYINPUT66), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT66), .B1(new_n231), .B2(new_n234), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n229), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n223), .B1(new_n227), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT30), .B1(new_n238), .B2(KEYINPUT64), .ZN(new_n239));
  INV_X1    g053(.A(new_n229), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n230), .A2(new_n204), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n198), .B2(new_n200), .ZN(new_n243));
  INV_X1    g057(.A(new_n233), .ZN(new_n244));
  NAND3_X1  g058(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n241), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n231), .A2(KEYINPUT66), .A3(new_n234), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n240), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n226), .A2(new_n222), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n249), .A2(new_n250), .B1(new_n222), .B2(new_n211), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT64), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT30), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(KEYINPUT69), .B(new_n195), .C1(new_n239), .C2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n195), .B(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n195), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n253), .B1(new_n251), .B2(new_n252), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n238), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(KEYINPUT69), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G101), .ZN(new_n266));
  INV_X1    g080(.A(G237), .ZN(new_n267));
  INV_X1    g081(.A(G953), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(G210), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n266), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n270), .B(new_n271), .Z(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n188), .B1(new_n265), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n195), .B(KEYINPUT70), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n238), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(new_n263), .B2(KEYINPUT69), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n195), .B1(new_n239), .B2(new_n254), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n277), .A2(new_n280), .A3(new_n188), .A4(new_n273), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n276), .A2(KEYINPUT28), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n238), .A2(new_n195), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT28), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n258), .A2(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  OR2_X1    g100(.A1(new_n286), .A2(new_n273), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT32), .B(new_n187), .C1(new_n274), .C2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT75), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n187), .B1(new_n274), .B2(new_n288), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n277), .A2(new_n273), .A3(new_n280), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT31), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(new_n287), .A3(new_n281), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(KEYINPUT75), .A3(KEYINPUT32), .A4(new_n187), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n272), .B1(new_n259), .B2(new_n264), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT29), .B1(new_n286), .B2(new_n273), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n238), .A2(new_n275), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(new_n258), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n251), .A2(KEYINPUT73), .A3(new_n257), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(KEYINPUT28), .A3(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n273), .A2(KEYINPUT29), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n285), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G902), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT74), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n308), .A2(new_n312), .A3(new_n309), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n301), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G472), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n291), .A2(new_n294), .A3(new_n298), .A4(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G217), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(G234), .B2(new_n309), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT23), .ZN(new_n319));
  INV_X1    g133(.A(G119), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n319), .B1(new_n320), .B2(G128), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n321), .B(new_n322), .C1(G119), .C2(new_n204), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G110), .ZN(new_n324));
  XOR2_X1   g138(.A(KEYINPUT24), .B(G110), .Z(new_n325));
  XNOR2_X1  g139(.A(G119), .B(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n329), .A2(KEYINPUT16), .A3(G140), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n330), .A2(KEYINPUT76), .ZN(new_n331));
  XNOR2_X1  g145(.A(G125), .B(G140), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n330), .B1(new_n332), .B2(KEYINPUT16), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n199), .ZN(new_n336));
  OAI211_X1 g150(.A(G146), .B(new_n331), .C1(new_n333), .C2(new_n334), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n328), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n268), .A2(G221), .A3(G234), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT77), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT22), .B(G137), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  OAI22_X1  g157(.A1(new_n323), .A2(G110), .B1(new_n326), .B2(new_n325), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n332), .A2(new_n199), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n337), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  OR3_X1    g160(.A1(new_n338), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n343), .B1(new_n338), .B2(new_n346), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT25), .B1(new_n349), .B2(new_n309), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT25), .ZN(new_n351));
  AOI211_X1 g165(.A(new_n351), .B(G902), .C1(new_n347), .C2(new_n348), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n318), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n318), .A2(G902), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n316), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(G214), .B1(G237), .B2(G902), .ZN(new_n359));
  XOR2_X1   g173(.A(new_n359), .B(KEYINPUT84), .Z(new_n360));
  NAND2_X1  g174(.A1(new_n249), .A2(G125), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n201), .A2(new_n205), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n329), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G224), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(G953), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n364), .B(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(G110), .B(G122), .ZN(new_n369));
  INV_X1    g183(.A(G104), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT3), .B1(new_n370), .B2(G107), .ZN(new_n371));
  AOI21_X1  g185(.A(G101), .B1(new_n370), .B2(G107), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n373));
  INV_X1    g187(.A(G107), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(G104), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT79), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n371), .A2(new_n372), .A3(new_n375), .A4(KEYINPUT79), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n370), .A2(G107), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n371), .A2(new_n375), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G101), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n382), .A2(KEYINPUT78), .A3(G101), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n380), .A2(new_n385), .A3(KEYINPUT4), .A4(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n382), .A2(new_n388), .A3(G101), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n195), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G113), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G116), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(G119), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n392), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n191), .A2(new_n393), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n397), .A2(new_n398), .B1(new_n191), .B2(new_n190), .ZN(new_n399));
  INV_X1    g213(.A(G101), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n370), .A2(G107), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n402), .B2(new_n381), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n378), .B2(new_n379), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n391), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n369), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n387), .A2(new_n390), .B1(new_n404), .B2(new_n399), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT86), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(KEYINPUT6), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n369), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n408), .A2(new_n410), .B1(KEYINPUT6), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n368), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(G210), .B1(G237), .B2(G902), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT7), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n417), .B1(new_n366), .B2(KEYINPUT88), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n364), .B(new_n418), .C1(KEYINPUT88), .C2(new_n366), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n361), .B(new_n363), .C1(new_n417), .C2(new_n366), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT5), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n397), .B1(new_n421), .B2(new_n193), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n192), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n404), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n378), .A2(new_n379), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n399), .B1(new_n425), .B2(new_n403), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT87), .B(KEYINPUT8), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n369), .B(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n424), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n419), .A2(new_n420), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n413), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n309), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n415), .A2(new_n416), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n416), .ZN(new_n435));
  INV_X1    g249(.A(new_n368), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n413), .A2(KEYINPUT6), .ZN(new_n437));
  INV_X1    g251(.A(new_n410), .ZN(new_n438));
  INV_X1    g252(.A(new_n369), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(new_n409), .B2(KEYINPUT86), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n437), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n436), .B1(new_n441), .B2(new_n411), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n435), .B1(new_n442), .B2(new_n432), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n360), .B1(new_n434), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(G475), .A2(G902), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n267), .A2(new_n268), .A3(G214), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(KEYINPUT89), .B2(new_n196), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT89), .B(G143), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n447), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n221), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT17), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n447), .B(new_n221), .C1(new_n446), .C2(new_n448), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n449), .A2(KEYINPUT17), .A3(new_n450), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n454), .A2(new_n336), .A3(new_n337), .A4(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G113), .B(G122), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT90), .B(G104), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n457), .B(new_n458), .Z(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(KEYINPUT18), .A2(G131), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n449), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n332), .B(new_n199), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n449), .A2(new_n461), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n456), .A2(new_n460), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n451), .A2(new_n453), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n332), .B(KEYINPUT19), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n199), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n337), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n460), .B1(new_n470), .B2(new_n465), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n445), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT20), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n460), .B1(new_n456), .B2(new_n465), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n309), .B1(new_n466), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G122), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT91), .B1(new_n479), .B2(G116), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT91), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n395), .A3(G122), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT14), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT93), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n395), .A2(G122), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT14), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(new_n480), .B2(new_n482), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT93), .B1(new_n490), .B2(new_n486), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n480), .A2(new_n482), .A3(new_n489), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G107), .ZN(new_n494));
  XNOR2_X1  g308(.A(G128), .B(G143), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(new_n206), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n483), .A2(new_n374), .A3(new_n487), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT92), .ZN(new_n501));
  AOI211_X1 g315(.A(G107), .B(new_n486), .C1(new_n480), .C2(new_n482), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n374), .B1(new_n483), .B2(new_n487), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n481), .B1(new_n395), .B2(G122), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n479), .A2(KEYINPUT91), .A3(G116), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n487), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G107), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n497), .A3(KEYINPUT92), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n495), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT13), .B1(new_n204), .B2(G143), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(new_n206), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n511), .B(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT9), .B(G234), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n517), .A2(new_n317), .A3(G953), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n500), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n518), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n498), .B1(new_n493), .B2(G107), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n514), .B1(new_n504), .B2(new_n509), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n519), .A2(KEYINPUT94), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT94), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n525), .B(new_n520), .C1(new_n521), .C2(new_n522), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n309), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G478), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n527), .A2(new_n532), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n478), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(G234), .A2(G237), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(G952), .A3(new_n268), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(G902), .A3(G953), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT21), .B(G898), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n537), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G469), .ZN(new_n546));
  XNOR2_X1  g360(.A(G110), .B(G140), .ZN(new_n547));
  INV_X1    g361(.A(G227), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(G953), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n547), .B(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT80), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n229), .B(new_n389), .C1(new_n235), .C2(new_n236), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n374), .A2(G104), .ZN(new_n555));
  OAI21_X1  g369(.A(G101), .B1(new_n401), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n201), .A2(new_n205), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT10), .B1(new_n425), .B2(new_n557), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n201), .A2(new_n205), .A3(new_n556), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT10), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n380), .A3(new_n560), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n387), .A2(new_n554), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n552), .B1(new_n562), .B2(new_n227), .ZN(new_n563));
  AND4_X1   g377(.A1(KEYINPUT4), .A2(new_n380), .A3(new_n385), .A4(new_n386), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n559), .A2(new_n380), .A3(new_n560), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n560), .B1(new_n559), .B2(new_n380), .ZN(new_n566));
  OAI22_X1  g380(.A1(new_n564), .A2(new_n553), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(KEYINPUT80), .A3(new_n250), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n558), .A2(new_n561), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n387), .A2(new_n249), .A3(new_n389), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n571), .A3(new_n227), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n551), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT82), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n551), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n380), .A2(new_n556), .B1(new_n205), .B2(new_n201), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n557), .B1(new_n378), .B2(new_n379), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n250), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT12), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT12), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n580), .B(new_n250), .C1(new_n576), .C2(new_n577), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n574), .B1(new_n575), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n550), .B1(new_n562), .B2(new_n227), .ZN(new_n584));
  INV_X1    g398(.A(new_n581), .ZN(new_n585));
  OAI22_X1  g399(.A1(new_n425), .A2(new_n557), .B1(new_n404), .B2(new_n362), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n580), .B1(new_n586), .B2(new_n250), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n584), .A2(KEYINPUT82), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n546), .B(new_n309), .C1(new_n573), .C2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n575), .B1(new_n563), .B2(new_n568), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n551), .B1(new_n588), .B2(new_n572), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT81), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI211_X1 g408(.A(new_n552), .B(new_n227), .C1(new_n570), .C2(new_n571), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT80), .B1(new_n567), .B2(new_n250), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n584), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT81), .ZN(new_n598));
  INV_X1    g412(.A(new_n572), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n550), .B1(new_n582), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n594), .A2(G469), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n546), .A2(new_n309), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n591), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT83), .ZN(new_n606));
  OAI21_X1  g420(.A(G221), .B1(new_n517), .B2(G902), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n606), .B1(new_n605), .B2(new_n607), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n444), .B(new_n545), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n358), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(new_n400), .ZN(G3));
  NAND2_X1  g426(.A1(new_n605), .A2(new_n607), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT83), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(G472), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n297), .B2(new_n309), .ZN(new_n618));
  INV_X1    g432(.A(new_n187), .ZN(new_n619));
  INV_X1    g433(.A(new_n288), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n619), .B1(new_n620), .B2(new_n296), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n616), .A2(new_n357), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n527), .A2(new_n528), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT99), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT99), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n527), .A2(new_n626), .A3(new_n528), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT96), .B(KEYINPUT33), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n524), .A2(new_n526), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT97), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n524), .A2(KEYINPUT97), .A3(new_n526), .A4(new_n629), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n523), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n523), .A2(new_n634), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n635), .A2(KEYINPUT33), .A3(new_n519), .A4(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n528), .A2(G902), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n632), .A2(new_n633), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n628), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT100), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n628), .A2(new_n642), .A3(new_n639), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n544), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n644), .A2(new_n444), .A3(new_n645), .A4(new_n477), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n623), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT34), .B(G104), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  NAND3_X1  g463(.A1(new_n475), .A2(KEYINPUT101), .A3(G475), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n473), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(new_n652), .B2(new_n476), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n535), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n544), .B(KEYINPUT102), .Z(new_n656));
  AND2_X1   g470(.A1(new_n444), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n623), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT35), .B(G107), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NOR2_X1   g476(.A1(new_n338), .A2(new_n346), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n342), .A2(KEYINPUT36), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n663), .B(new_n664), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n354), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n353), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n478), .A2(new_n536), .A3(new_n645), .A4(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n616), .A2(new_n444), .A3(new_n622), .A4(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  INV_X1    g486(.A(new_n444), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n614), .B2(new_n615), .ZN(new_n674));
  INV_X1    g488(.A(G900), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n540), .B1(new_n542), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n654), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n674), .A2(new_n316), .A3(new_n667), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  XOR2_X1   g493(.A(new_n676), .B(KEYINPUT39), .Z(new_n680));
  NAND2_X1  g494(.A1(new_n616), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n265), .A2(new_n272), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n304), .A2(new_n305), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n309), .B1(new_n684), .B2(new_n273), .ZN(new_n685));
  OAI21_X1  g499(.A(G472), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n291), .A2(new_n294), .A3(new_n298), .A4(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n434), .A2(new_n443), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n477), .A2(new_n535), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n690), .A2(new_n360), .A3(new_n667), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n682), .A2(new_n687), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  NAND4_X1  g509(.A1(new_n316), .A2(new_n616), .A3(new_n444), .A4(new_n667), .ZN(new_n696));
  INV_X1    g510(.A(new_n676), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n628), .A2(new_n642), .A3(new_n639), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n642), .B1(new_n628), .B2(new_n639), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n477), .B(new_n697), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n644), .A2(KEYINPUT104), .A3(new_n477), .A4(new_n697), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n696), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT105), .B(G146), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G48));
  INV_X1    g521(.A(new_n646), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n309), .B1(new_n573), .B2(new_n590), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G469), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n607), .ZN(new_n712));
  INV_X1    g526(.A(new_n591), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n708), .A2(new_n316), .A3(new_n357), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT41), .B(G113), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NAND4_X1  g531(.A1(new_n658), .A2(new_n316), .A3(new_n714), .A4(new_n357), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  AND4_X1   g533(.A1(new_n607), .A2(new_n444), .A3(new_n591), .A4(new_n710), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n316), .A2(new_n669), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  NAND3_X1  g536(.A1(new_n444), .A2(new_n535), .A3(new_n477), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n710), .A2(new_n607), .A3(new_n591), .A4(new_n656), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n306), .A2(new_n285), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n306), .A2(KEYINPUT106), .A3(new_n285), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n272), .A3(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n296), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n281), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n731), .B1(new_n730), .B2(new_n296), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n187), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n618), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n725), .A2(new_n735), .A3(new_n357), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  AND2_X1   g552(.A1(new_n702), .A2(new_n703), .ZN(new_n739));
  AND4_X1   g553(.A1(new_n736), .A2(new_n720), .A3(new_n735), .A4(new_n667), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  INV_X1    g557(.A(new_n360), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n434), .A2(new_n443), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n592), .A2(new_n593), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n603), .B1(new_n747), .B2(G469), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n591), .A2(new_n748), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n746), .A2(new_n607), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n316), .A2(new_n357), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n743), .B1(new_n751), .B2(new_n704), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n315), .A2(new_n289), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT32), .B1(new_n297), .B2(new_n187), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n753), .B(new_n357), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT32), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n292), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n289), .A3(new_n315), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n753), .B1(new_n760), .B2(new_n357), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT42), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n702), .A2(new_n703), .A3(new_n750), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n752), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  NAND4_X1  g579(.A1(new_n316), .A2(new_n357), .A3(new_n677), .A4(new_n750), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  NAND2_X1  g581(.A1(new_n644), .A2(new_n478), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT43), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n736), .A2(new_n292), .B1(new_n353), .B2(new_n666), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n644), .A2(new_n771), .A3(new_n478), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n769), .A2(new_n770), .A3(KEYINPUT44), .A4(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n746), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n594), .A2(new_n601), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n546), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT45), .B1(new_n594), .B2(new_n601), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT109), .B1(new_n780), .B2(new_n546), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n592), .A2(new_n593), .A3(new_n776), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n779), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT46), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n603), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT110), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n784), .A2(new_n789), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT46), .B1(new_n784), .B2(new_n604), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n713), .B1(new_n792), .B2(KEYINPUT111), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n782), .B1(new_n777), .B2(new_n778), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n603), .B1(new_n795), .B2(new_n781), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n794), .B1(new_n796), .B2(KEYINPUT46), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n791), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n680), .A2(new_n607), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n774), .A2(new_n798), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  AOI21_X1  g618(.A(new_n789), .B1(new_n784), .B2(new_n786), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n784), .A2(new_n789), .A3(new_n786), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n797), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n784), .A2(new_n604), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(KEYINPUT111), .A3(new_n785), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n591), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n607), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT47), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT47), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n813), .B(new_n607), .C1(new_n807), .C2(new_n810), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n704), .A2(new_n316), .A3(new_n357), .A4(new_n745), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  INV_X1    g631(.A(G952), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n268), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n769), .A2(new_n540), .A3(new_n772), .ZN(new_n820));
  INV_X1    g634(.A(new_n714), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n820), .A2(new_n821), .A3(new_n745), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n757), .B2(new_n761), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT48), .ZN(new_n824));
  INV_X1    g638(.A(new_n820), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n735), .A2(new_n357), .A3(new_n736), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n720), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n714), .A2(new_n357), .A3(new_n540), .A4(new_n746), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n687), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n478), .B1(new_n641), .B2(new_n643), .ZN(new_n831));
  AOI211_X1 g645(.A(new_n818), .B(G953), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n824), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n735), .A2(new_n736), .A3(new_n667), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n644), .A2(new_n477), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n822), .A2(new_n835), .B1(new_n830), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n769), .A2(new_n772), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n690), .A2(new_n360), .A3(new_n714), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n838), .A2(new_n540), .A3(new_n827), .A4(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT50), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT117), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n820), .A2(new_n839), .A3(new_n826), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT116), .B1(new_n844), .B2(KEYINPUT50), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n841), .A2(new_n846), .A3(new_n842), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n844), .A2(new_n848), .A3(KEYINPUT50), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n843), .A2(new_n845), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n711), .A2(new_n713), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n812), .A2(new_n814), .B1(new_n712), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n825), .A2(new_n827), .A3(new_n746), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n837), .B(new_n850), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n854), .A2(KEYINPUT115), .A3(KEYINPUT51), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT51), .B1(new_n854), .B2(KEYINPUT115), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n833), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n291), .A2(new_n294), .A3(new_n298), .A4(new_n315), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n444), .B(new_n667), .C1(new_n608), .C2(new_n609), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n677), .A2(new_n861), .B1(new_n739), .B2(new_n740), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n353), .A2(new_n666), .A3(new_n697), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n749), .A2(new_n863), .A3(new_n607), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT113), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n673), .A2(new_n691), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n749), .A2(new_n863), .A3(new_n867), .A4(new_n607), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n861), .A2(new_n739), .B1(new_n687), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n862), .A2(new_n870), .A3(KEYINPUT52), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n720), .A2(new_n735), .A3(new_n736), .A4(new_n667), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n678), .B1(new_n704), .B2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n687), .A2(new_n866), .A3(new_n865), .A4(new_n868), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n696), .B2(new_n704), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n872), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n715), .A2(new_n718), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n616), .A2(new_n357), .A3(new_n622), .A4(new_n657), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n537), .B1(new_n644), .B2(new_n478), .ZN(new_n881));
  OAI22_X1  g695(.A1(new_n880), .A2(new_n881), .B1(new_n358), .B2(new_n610), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n670), .A2(new_n721), .A3(new_n737), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n879), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n536), .A2(new_n653), .A3(new_n667), .A4(new_n697), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n316), .A2(new_n616), .A3(new_n746), .A4(new_n885), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n886), .B(new_n766), .C1(new_n763), .C2(new_n834), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n884), .A2(new_n764), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n858), .B1(new_n878), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n882), .A2(new_n883), .ZN(new_n891));
  INV_X1    g705(.A(new_n879), .ZN(new_n892));
  AND4_X1   g706(.A1(new_n764), .A2(new_n891), .A3(new_n892), .A4(new_n888), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT114), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n871), .A2(new_n877), .A3(new_n894), .ZN(new_n895));
  OAI211_X1 g709(.A(KEYINPUT114), .B(new_n872), .C1(new_n874), .C2(new_n876), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n893), .A2(new_n895), .A3(KEYINPUT53), .A4(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n890), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n878), .A2(new_n889), .A3(new_n858), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n858), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n899), .B1(new_n902), .B2(new_n898), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n819), .B1(new_n857), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n851), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(KEYINPUT49), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT112), .Z(new_n907));
  NOR3_X1   g721(.A1(new_n356), .A2(new_n712), .A3(new_n360), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT49), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n690), .B(new_n908), .C1(new_n909), .C2(new_n851), .ZN(new_n910));
  OR4_X1    g724(.A1(new_n687), .A2(new_n907), .A3(new_n768), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n904), .A2(new_n911), .ZN(G75));
  NOR2_X1   g726(.A1(new_n268), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n309), .B1(new_n890), .B2(new_n897), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT56), .B1(new_n915), .B2(G210), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n412), .A2(new_n414), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n436), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n415), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT55), .Z(new_n920));
  OAI21_X1  g734(.A(new_n914), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT56), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n915), .ZN(new_n925));
  INV_X1    g739(.A(G210), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT118), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT118), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n929), .B(new_n924), .C1(new_n925), .C2(new_n926), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n921), .B1(new_n928), .B2(new_n930), .ZN(G51));
  XNOR2_X1  g745(.A(new_n603), .B(KEYINPUT57), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n890), .A2(new_n897), .A3(new_n898), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n898), .B1(new_n890), .B2(new_n897), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n573), .B2(new_n590), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n784), .B(KEYINPUT119), .Z(new_n937));
  NAND2_X1  g751(.A1(new_n915), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n913), .B1(new_n936), .B2(new_n938), .ZN(G54));
  NAND2_X1  g753(.A1(new_n890), .A2(new_n897), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n466), .A2(new_n471), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(KEYINPUT58), .A2(G475), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n940), .A2(G902), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT120), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n915), .A2(new_n943), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n913), .B1(new_n948), .B2(new_n941), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(G60));
  NAND3_X1  g764(.A1(new_n632), .A2(new_n633), .A3(new_n637), .ZN(new_n951));
  NAND2_X1  g765(.A1(G478), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT59), .Z(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n933), .B2(new_n934), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n914), .ZN(new_n956));
  INV_X1    g770(.A(new_n953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n903), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n958), .B2(new_n951), .ZN(G63));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n960));
  NAND2_X1  g774(.A1(G217), .A2(G902), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT60), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n890), .B2(new_n897), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n665), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n914), .B1(new_n963), .B2(new_n349), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n960), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n963), .A2(new_n349), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n968), .A2(KEYINPUT61), .A3(new_n914), .A4(new_n964), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(G66));
  OAI21_X1  g784(.A(G953), .B1(new_n543), .B2(new_n365), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n884), .B2(G953), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n917), .B1(G898), .B2(new_n268), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT121), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n972), .B(new_n974), .ZN(G69));
  INV_X1    g789(.A(new_n761), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n723), .B1(new_n976), .B2(new_n756), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n798), .A2(new_n977), .A3(new_n802), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n978), .A2(new_n764), .A3(new_n766), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT122), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n874), .B2(new_n705), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n861), .A2(new_n739), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n982), .A2(new_n741), .A3(KEYINPUT122), .A4(new_n678), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n979), .A2(new_n816), .A3(new_n984), .A4(new_n803), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(KEYINPUT125), .ZN(new_n986));
  AND4_X1   g800(.A1(new_n764), .A2(new_n803), .A3(new_n766), .A4(new_n978), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT125), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n987), .A2(new_n988), .A3(new_n816), .A4(new_n984), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n986), .A2(new_n989), .A3(new_n268), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n261), .A2(new_n262), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(new_n468), .Z(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(G900), .B2(G953), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT123), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n981), .A2(new_n694), .A3(new_n983), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT62), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n981), .A2(KEYINPUT62), .A3(new_n983), .A4(new_n694), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OR4_X1    g814(.A1(new_n358), .A2(new_n681), .A3(new_n745), .A4(new_n881), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n801), .B(new_n802), .C1(new_n807), .C2(new_n810), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n773), .A2(new_n746), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n814), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n813), .B1(new_n798), .B2(new_n607), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1004), .B1(new_n1007), .B2(new_n815), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n1000), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n995), .B(new_n992), .C1(new_n1009), .C2(G953), .ZN(new_n1010));
  AOI21_X1  g824(.A(G953), .B1(new_n1000), .B2(new_n1008), .ZN(new_n1011));
  INV_X1    g825(.A(new_n992), .ZN(new_n1012));
  OAI21_X1  g826(.A(KEYINPUT123), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g827(.A(G953), .B1(new_n548), .B2(new_n675), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT124), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n994), .A2(new_n1010), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1017), .B1(new_n990), .B2(new_n993), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1016), .B1(new_n1014), .B2(new_n1018), .ZN(G72));
  NAND3_X1  g833(.A1(new_n1000), .A2(new_n1008), .A3(new_n884), .ZN(new_n1020));
  XNOR2_X1  g834(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n617), .A2(new_n309), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1021), .B(new_n1022), .Z(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(KEYINPUT127), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT127), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1020), .A2(new_n1027), .A3(new_n1024), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1026), .A2(new_n683), .A3(new_n1028), .ZN(new_n1029));
  NOR3_X1   g843(.A1(new_n259), .A2(new_n264), .A3(new_n273), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n986), .A2(new_n884), .A3(new_n989), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1030), .B1(new_n1031), .B2(new_n1023), .ZN(new_n1032));
  INV_X1    g846(.A(new_n902), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1023), .B1(new_n299), .B2(new_n295), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n913), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AND3_X1   g849(.A1(new_n1029), .A2(new_n1032), .A3(new_n1035), .ZN(G57));
endmodule


