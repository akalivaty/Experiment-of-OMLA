

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588;

  XNOR2_X1 U321 ( .A(n399), .B(KEYINPUT48), .ZN(n400) );
  XNOR2_X1 U322 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U323 ( .A(n401), .B(n400), .ZN(n536) );
  XNOR2_X1 U324 ( .A(n413), .B(n315), .ZN(n316) );
  XNOR2_X1 U325 ( .A(n435), .B(n316), .ZN(n317) );
  XNOR2_X1 U326 ( .A(n414), .B(n348), .ZN(n349) );
  XNOR2_X1 U327 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U328 ( .A(n325), .B(n324), .ZN(n334) );
  XNOR2_X1 U329 ( .A(n455), .B(KEYINPUT122), .ZN(n568) );
  XNOR2_X1 U330 ( .A(KEYINPUT95), .B(n477), .ZN(n523) );
  XNOR2_X1 U331 ( .A(n456), .B(KEYINPUT124), .ZN(n457) );
  XNOR2_X1 U332 ( .A(n458), .B(n457), .ZN(G1350GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT6), .B(KEYINPUT91), .Z(n290) );
  XNOR2_X1 U334 ( .A(G1GAT), .B(G162GAT), .ZN(n289) );
  XNOR2_X1 U335 ( .A(n290), .B(n289), .ZN(n294) );
  XOR2_X1 U336 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n292) );
  XNOR2_X1 U337 ( .A(KEYINPUT92), .B(KEYINPUT1), .ZN(n291) );
  XNOR2_X1 U338 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U339 ( .A(n294), .B(n293), .Z(n299) );
  XOR2_X1 U340 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n296) );
  NAND2_X1 U341 ( .A1(G225GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U343 ( .A(KEYINPUT94), .B(n297), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n304) );
  XNOR2_X1 U345 ( .A(G120GAT), .B(G148GAT), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n300), .B(G57GAT), .ZN(n344) );
  XOR2_X1 U347 ( .A(G29GAT), .B(KEYINPUT78), .Z(n319) );
  XOR2_X1 U348 ( .A(n344), .B(n319), .Z(n302) );
  XNOR2_X1 U349 ( .A(G134GAT), .B(G85GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U351 ( .A(n304), .B(n303), .Z(n310) );
  XOR2_X1 U352 ( .A(G127GAT), .B(KEYINPUT0), .Z(n306) );
  XNOR2_X1 U353 ( .A(G113GAT), .B(KEYINPUT84), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n444) );
  XOR2_X1 U355 ( .A(G155GAT), .B(KEYINPUT3), .Z(n308) );
  XNOR2_X1 U356 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n421) );
  XNOR2_X1 U358 ( .A(n444), .B(n421), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n477) );
  XOR2_X1 U360 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n312) );
  XNOR2_X1 U361 ( .A(KEYINPUT76), .B(KEYINPUT11), .ZN(n311) );
  XNOR2_X1 U362 ( .A(n312), .B(n311), .ZN(n318) );
  XOR2_X1 U363 ( .A(G162GAT), .B(KEYINPUT75), .Z(n314) );
  XNOR2_X1 U364 ( .A(G50GAT), .B(G218GAT), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n435) );
  XOR2_X1 U366 ( .A(G36GAT), .B(G190GAT), .Z(n413) );
  AND2_X1 U367 ( .A1(G232GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n325) );
  XOR2_X1 U369 ( .A(G43GAT), .B(G134GAT), .Z(n445) );
  XOR2_X1 U370 ( .A(n445), .B(n319), .Z(n323) );
  XOR2_X1 U371 ( .A(KEYINPUT65), .B(KEYINPUT79), .Z(n321) );
  XNOR2_X1 U372 ( .A(KEYINPUT77), .B(KEYINPUT66), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U374 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n326), .B(KEYINPUT7), .ZN(n355) );
  XNOR2_X1 U376 ( .A(G99GAT), .B(G106GAT), .ZN(n332) );
  INV_X1 U377 ( .A(G85GAT), .ZN(n327) );
  NAND2_X1 U378 ( .A1(n327), .A2(G92GAT), .ZN(n330) );
  INV_X1 U379 ( .A(G92GAT), .ZN(n328) );
  NAND2_X1 U380 ( .A1(n328), .A2(G85GAT), .ZN(n329) );
  NAND2_X1 U381 ( .A1(n330), .A2(n329), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n337) );
  XOR2_X1 U383 ( .A(n355), .B(n337), .Z(n333) );
  XNOR2_X1 U384 ( .A(n334), .B(n333), .ZN(n562) );
  XNOR2_X1 U385 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n371) );
  XOR2_X1 U386 ( .A(KEYINPUT73), .B(KEYINPUT13), .Z(n336) );
  XNOR2_X1 U387 ( .A(KEYINPUT72), .B(KEYINPUT32), .ZN(n335) );
  XNOR2_X1 U388 ( .A(n336), .B(n335), .ZN(n352) );
  XNOR2_X1 U389 ( .A(n337), .B(KEYINPUT33), .ZN(n341) );
  INV_X1 U390 ( .A(n341), .ZN(n339) );
  NAND2_X1 U391 ( .A1(G230GAT), .A2(G233GAT), .ZN(n340) );
  INV_X1 U392 ( .A(n340), .ZN(n338) );
  NAND2_X1 U393 ( .A1(n339), .A2(n338), .ZN(n343) );
  NAND2_X1 U394 ( .A1(n341), .A2(n340), .ZN(n342) );
  NAND2_X1 U395 ( .A1(n343), .A2(n342), .ZN(n345) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n347) );
  XOR2_X1 U397 ( .A(G176GAT), .B(G71GAT), .Z(n448) );
  XOR2_X1 U398 ( .A(KEYINPUT71), .B(G78GAT), .Z(n422) );
  XOR2_X1 U399 ( .A(n448), .B(n422), .Z(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n350) );
  XOR2_X1 U401 ( .A(G204GAT), .B(G64GAT), .Z(n414) );
  XNOR2_X1 U402 ( .A(KEYINPUT70), .B(KEYINPUT31), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n352), .B(n351), .ZN(n393) );
  XNOR2_X1 U404 ( .A(n393), .B(KEYINPUT41), .ZN(n506) );
  XOR2_X1 U405 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n358) );
  XOR2_X1 U406 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n354) );
  XNOR2_X1 U407 ( .A(G197GAT), .B(G141GAT), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n356) );
  XNOR2_X1 U409 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U410 ( .A(n358), .B(n357), .ZN(n364) );
  XOR2_X1 U411 ( .A(G1GAT), .B(G8GAT), .Z(n360) );
  XNOR2_X1 U412 ( .A(G15GAT), .B(G22GAT), .ZN(n359) );
  XNOR2_X1 U413 ( .A(n360), .B(n359), .ZN(n378) );
  XOR2_X1 U414 ( .A(G29GAT), .B(n378), .Z(n362) );
  NAND2_X1 U415 ( .A1(G229GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U417 ( .A(n364), .B(n363), .Z(n369) );
  XOR2_X1 U418 ( .A(G113GAT), .B(G50GAT), .Z(n366) );
  XNOR2_X1 U419 ( .A(G169GAT), .B(G43GAT), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U421 ( .A(n367), .B(G36GAT), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n369), .B(n368), .ZN(n574) );
  NOR2_X1 U423 ( .A1(n506), .A2(n574), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n371), .B(n370), .ZN(n389) );
  XOR2_X1 U425 ( .A(G211GAT), .B(G127GAT), .Z(n373) );
  XNOR2_X1 U426 ( .A(G183GAT), .B(G71GAT), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U428 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n375) );
  NAND2_X1 U429 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U431 ( .A(n377), .B(n376), .Z(n380) );
  XNOR2_X1 U432 ( .A(n378), .B(KEYINPUT82), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n380), .B(n379), .ZN(n388) );
  XOR2_X1 U434 ( .A(G64GAT), .B(G57GAT), .Z(n382) );
  XNOR2_X1 U435 ( .A(G155GAT), .B(G78GAT), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U437 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n384) );
  XNOR2_X1 U438 ( .A(KEYINPUT13), .B(KEYINPUT12), .ZN(n383) );
  XNOR2_X1 U439 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U440 ( .A(n386), .B(n385), .Z(n387) );
  XOR2_X1 U441 ( .A(n388), .B(n387), .Z(n558) );
  INV_X1 U442 ( .A(n558), .ZN(n584) );
  NOR2_X1 U443 ( .A1(n389), .A2(n584), .ZN(n390) );
  AND2_X1 U444 ( .A1(n562), .A2(n390), .ZN(n392) );
  INV_X1 U445 ( .A(KEYINPUT47), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n398) );
  XNOR2_X1 U447 ( .A(KEYINPUT80), .B(n562), .ZN(n459) );
  XNOR2_X1 U448 ( .A(KEYINPUT36), .B(n459), .ZN(n490) );
  NOR2_X1 U449 ( .A1(n490), .A2(n558), .ZN(n394) );
  XNOR2_X1 U450 ( .A(n394), .B(KEYINPUT45), .ZN(n395) );
  NAND2_X1 U451 ( .A1(n395), .A2(n574), .ZN(n396) );
  NOR2_X1 U452 ( .A1(n393), .A2(n396), .ZN(n397) );
  NOR2_X1 U453 ( .A1(n398), .A2(n397), .ZN(n401) );
  XOR2_X1 U454 ( .A(KEYINPUT64), .B(KEYINPUT115), .Z(n399) );
  XOR2_X1 U455 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n403) );
  XNOR2_X1 U456 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U458 ( .A(G169GAT), .B(n404), .Z(n443) );
  XOR2_X1 U459 ( .A(G211GAT), .B(KEYINPUT21), .Z(n406) );
  XNOR2_X1 U460 ( .A(G197GAT), .B(KEYINPUT89), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n434) );
  XOR2_X1 U462 ( .A(KEYINPUT96), .B(n434), .Z(n408) );
  NAND2_X1 U463 ( .A1(G226GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U465 ( .A(G92GAT), .B(G218GAT), .Z(n410) );
  XNOR2_X1 U466 ( .A(G8GAT), .B(G176GAT), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U468 ( .A(n412), .B(n411), .Z(n416) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U471 ( .A(n443), .B(n417), .Z(n526) );
  INV_X1 U472 ( .A(n526), .ZN(n466) );
  NOR2_X1 U473 ( .A1(n536), .A2(n466), .ZN(n419) );
  INV_X1 U474 ( .A(KEYINPUT54), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n420) );
  NOR2_X1 U476 ( .A1(n523), .A2(n420), .ZN(n573) );
  XOR2_X1 U477 ( .A(n422), .B(n421), .Z(n424) );
  XNOR2_X1 U478 ( .A(G106GAT), .B(KEYINPUT87), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U480 ( .A(G204GAT), .B(G148GAT), .Z(n426) );
  NAND2_X1 U481 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U483 ( .A(n428), .B(n427), .Z(n433) );
  XOR2_X1 U484 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n430) );
  XNOR2_X1 U485 ( .A(KEYINPUT88), .B(KEYINPUT23), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U487 ( .A(G22GAT), .B(n431), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U489 ( .A(n435), .B(n434), .Z(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n471) );
  NAND2_X1 U491 ( .A1(n573), .A2(n471), .ZN(n439) );
  XOR2_X1 U492 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n454) );
  XOR2_X1 U494 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n441) );
  XNOR2_X1 U495 ( .A(G15GAT), .B(G120GAT), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n453) );
  XOR2_X1 U498 ( .A(n445), .B(n444), .Z(n447) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n449) );
  XOR2_X1 U501 ( .A(n449), .B(n448), .Z(n451) );
  XNOR2_X1 U502 ( .A(G190GAT), .B(G99GAT), .ZN(n450) );
  XNOR2_X1 U503 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U504 ( .A(n453), .B(n452), .Z(n537) );
  INV_X1 U505 ( .A(n537), .ZN(n529) );
  NAND2_X1 U506 ( .A1(n454), .A2(n529), .ZN(n455) );
  NOR2_X1 U507 ( .A1(n568), .A2(n558), .ZN(n458) );
  INV_X1 U508 ( .A(G183GAT), .ZN(n456) );
  INV_X1 U509 ( .A(G190GAT), .ZN(n462) );
  NOR2_X1 U510 ( .A1(n568), .A2(n459), .ZN(n460) );
  XNOR2_X1 U511 ( .A(KEYINPUT58), .B(n460), .ZN(n461) );
  XNOR2_X1 U512 ( .A(n462), .B(n461), .ZN(G1351GAT) );
  NOR2_X1 U513 ( .A1(n393), .A2(n574), .ZN(n463) );
  XOR2_X1 U514 ( .A(n463), .B(KEYINPUT74), .Z(n494) );
  NAND2_X1 U515 ( .A1(n459), .A2(n584), .ZN(n464) );
  XOR2_X1 U516 ( .A(KEYINPUT16), .B(n464), .Z(n480) );
  XNOR2_X1 U517 ( .A(KEYINPUT27), .B(n526), .ZN(n473) );
  NAND2_X1 U518 ( .A1(n523), .A2(n473), .ZN(n551) );
  XOR2_X1 U519 ( .A(KEYINPUT28), .B(n471), .Z(n531) );
  NOR2_X1 U520 ( .A1(n551), .A2(n531), .ZN(n539) );
  XNOR2_X1 U521 ( .A(n537), .B(KEYINPUT86), .ZN(n465) );
  NAND2_X1 U522 ( .A1(n539), .A2(n465), .ZN(n479) );
  NOR2_X1 U523 ( .A1(n537), .A2(n466), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n467), .B(KEYINPUT97), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n468), .A2(n471), .ZN(n470) );
  XOR2_X1 U526 ( .A(KEYINPUT25), .B(KEYINPUT98), .Z(n469) );
  XNOR2_X1 U527 ( .A(n470), .B(n469), .ZN(n475) );
  NOR2_X1 U528 ( .A1(n471), .A2(n529), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n472), .B(KEYINPUT26), .ZN(n572) );
  NAND2_X1 U530 ( .A1(n572), .A2(n473), .ZN(n474) );
  NAND2_X1 U531 ( .A1(n475), .A2(n474), .ZN(n476) );
  NAND2_X1 U532 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U533 ( .A1(n479), .A2(n478), .ZN(n491) );
  NAND2_X1 U534 ( .A1(n480), .A2(n491), .ZN(n507) );
  NOR2_X1 U535 ( .A1(n494), .A2(n507), .ZN(n487) );
  NAND2_X1 U536 ( .A1(n487), .A2(n523), .ZN(n481) );
  XNOR2_X1 U537 ( .A(KEYINPUT34), .B(n481), .ZN(n482) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  XOR2_X1 U539 ( .A(G8GAT), .B(KEYINPUT99), .Z(n484) );
  NAND2_X1 U540 ( .A1(n487), .A2(n526), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U543 ( .A1(n487), .A2(n529), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NAND2_X1 U545 ( .A1(n531), .A2(n487), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n488), .B(KEYINPUT100), .ZN(n489) );
  XNOR2_X1 U547 ( .A(G22GAT), .B(n489), .ZN(G1327GAT) );
  XOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .Z(n498) );
  NAND2_X1 U549 ( .A1(n558), .A2(n491), .ZN(n492) );
  NOR2_X1 U550 ( .A1(n490), .A2(n492), .ZN(n493) );
  XNOR2_X1 U551 ( .A(KEYINPUT37), .B(n493), .ZN(n522) );
  OR2_X1 U552 ( .A1(n494), .A2(n522), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n495), .B(KEYINPUT101), .ZN(n496) );
  XNOR2_X1 U554 ( .A(KEYINPUT38), .B(n496), .ZN(n503) );
  NAND2_X1 U555 ( .A1(n503), .A2(n523), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(KEYINPUT102), .ZN(n500) );
  NAND2_X1 U558 ( .A1(n526), .A2(n503), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(G1329GAT) );
  NAND2_X1 U560 ( .A1(n503), .A2(n529), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n501), .B(KEYINPUT40), .ZN(n502) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  XOR2_X1 U563 ( .A(G50GAT), .B(KEYINPUT103), .Z(n505) );
  NAND2_X1 U564 ( .A1(n503), .A2(n531), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n505), .B(n504), .ZN(G1331GAT) );
  XNOR2_X1 U566 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n512) );
  XOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT107), .Z(n510) );
  XOR2_X1 U568 ( .A(n506), .B(KEYINPUT104), .Z(n541) );
  NAND2_X1 U569 ( .A1(n574), .A2(n541), .ZN(n521) );
  NOR2_X1 U570 ( .A1(n521), .A2(n507), .ZN(n508) );
  XOR2_X1 U571 ( .A(KEYINPUT105), .B(n508), .Z(n516) );
  NAND2_X1 U572 ( .A1(n516), .A2(n523), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n512), .B(n511), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n516), .A2(n526), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n513), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n516), .A2(n529), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n514), .B(KEYINPUT108), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(n515), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U581 ( .A1(n516), .A2(n531), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(n520) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT110), .Z(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  XOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT111), .Z(n525) );
  NOR2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n532) );
  NAND2_X1 U587 ( .A1(n532), .A2(n523), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U589 ( .A1(n532), .A2(n526), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n527), .B(KEYINPUT112), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G92GAT), .B(n528), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n532), .A2(n529), .ZN(n530) );
  XNOR2_X1 U593 ( .A(n530), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n534) );
  NAND2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U596 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n535), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n536), .A2(n537), .ZN(n538) );
  NAND2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n547) );
  NOR2_X1 U600 ( .A1(n574), .A2(n547), .ZN(n540) );
  XOR2_X1 U601 ( .A(G113GAT), .B(n540), .Z(G1340GAT) );
  INV_X1 U602 ( .A(n541), .ZN(n567) );
  NOR2_X1 U603 ( .A1(n567), .A2(n547), .ZN(n543) );
  XNOR2_X1 U604 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(n544), .ZN(G1341GAT) );
  NOR2_X1 U607 ( .A1(n558), .A2(n547), .ZN(n545) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(n545), .Z(n546) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  NOR2_X1 U610 ( .A1(n459), .A2(n547), .ZN(n549) );
  XNOR2_X1 U611 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n548) );
  XNOR2_X1 U612 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U613 ( .A(G134GAT), .B(n550), .Z(G1343GAT) );
  NOR2_X1 U614 ( .A1(n536), .A2(n551), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n552), .A2(n572), .ZN(n561) );
  NOR2_X1 U616 ( .A1(n574), .A2(n561), .ZN(n553) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n553), .Z(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n555) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(n557) );
  NOR2_X1 U621 ( .A1(n506), .A2(n561), .ZN(n556) );
  XOR2_X1 U622 ( .A(n557), .B(n556), .Z(G1345GAT) );
  NOR2_X1 U623 ( .A1(n558), .A2(n561), .ZN(n560) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1346GAT) );
  NOR2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U627 ( .A(KEYINPUT120), .B(n563), .Z(n564) );
  XNOR2_X1 U628 ( .A(G162GAT), .B(n564), .ZN(G1347GAT) );
  NOR2_X1 U629 ( .A1(n568), .A2(n574), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(G169GAT), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(KEYINPUT123), .ZN(G1348GAT) );
  NOR2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n570) );
  XNOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(n571), .ZN(G1349GAT) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n586) );
  NOR2_X1 U637 ( .A1(n574), .A2(n586), .ZN(n579) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n576) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(n577), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n581) );
  INV_X1 U644 ( .A(n586), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n583), .A2(n393), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(G204GAT), .B(n582), .Z(G1353GAT) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U650 ( .A1(n490), .A2(n586), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

