

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730;

  NOR2_X1 U370 ( .A1(n506), .A2(n505), .ZN(n508) );
  INV_X1 U371 ( .A(n663), .ZN(n498) );
  INV_X1 U372 ( .A(G472), .ZN(n355) );
  XNOR2_X1 U373 ( .A(n716), .B(G146), .ZN(n429) );
  XNOR2_X2 U374 ( .A(n391), .B(n371), .ZN(n408) );
  NOR2_X1 U375 ( .A1(n646), .A2(n650), .ZN(n687) );
  XNOR2_X1 U376 ( .A(n450), .B(n449), .ZN(n668) );
  OR2_X2 U377 ( .A1(n633), .A2(G902), .ZN(n431) );
  NOR2_X1 U378 ( .A1(G953), .A2(G237), .ZN(n409) );
  AND2_X1 U379 ( .A1(n727), .A2(n573), .ZN(n574) );
  NOR2_X2 U380 ( .A1(n568), .A2(n567), .ZN(n651) );
  INV_X1 U381 ( .A(KEYINPUT47), .ZN(n349) );
  INV_X1 U382 ( .A(n581), .ZN(n351) );
  OR2_X1 U383 ( .A1(n548), .A2(n547), .ZN(n568) );
  XNOR2_X1 U384 ( .A(n369), .B(n368), .ZN(n486) );
  XNOR2_X1 U385 ( .A(n404), .B(n403), .ZN(n464) );
  XNOR2_X1 U386 ( .A(n349), .B(n651), .ZN(n570) );
  INV_X1 U387 ( .A(n510), .ZN(n350) );
  INV_X1 U388 ( .A(n497), .ZN(n499) );
  AND2_X1 U389 ( .A1(n658), .A2(n352), .ZN(n353) );
  INV_X1 U390 ( .A(n580), .ZN(n352) );
  AND2_X1 U391 ( .A1(n351), .A2(n352), .ZN(n589) );
  INV_X1 U392 ( .A(n519), .ZN(n354) );
  XNOR2_X1 U393 ( .A(n508), .B(n507), .ZN(n620) );
  XNOR2_X2 U394 ( .A(n356), .B(n355), .ZN(n545) );
  NOR2_X1 U395 ( .A1(n606), .A2(G902), .ZN(n356) );
  NOR2_X1 U396 ( .A1(n620), .A2(KEYINPUT44), .ZN(n509) );
  XNOR2_X2 U397 ( .A(n408), .B(n407), .ZN(n716) );
  NOR2_X1 U398 ( .A1(n515), .A2(n728), .ZN(n520) );
  INV_X1 U399 ( .A(KEYINPUT88), .ZN(n516) );
  XNOR2_X1 U400 ( .A(G119), .B(G116), .ZN(n383) );
  INV_X1 U401 ( .A(KEYINPUT33), .ZN(n501) );
  NOR2_X1 U402 ( .A1(n500), .A2(n664), .ZN(n502) );
  XNOR2_X1 U403 ( .A(n545), .B(KEYINPUT6), .ZN(n497) );
  INV_X1 U404 ( .A(G134), .ZN(n371) );
  BUF_X1 U405 ( .A(n503), .Z(n528) );
  BUF_X1 U406 ( .A(n532), .Z(n653) );
  NAND2_X1 U407 ( .A1(n586), .A2(n585), .ZN(n659) );
  XNOR2_X2 U408 ( .A(n390), .B(n357), .ZN(n717) );
  BUF_X1 U409 ( .A(n621), .Z(n631) );
  XOR2_X2 U410 ( .A(n381), .B(G478), .Z(n487) );
  NOR2_X2 U411 ( .A1(n627), .A2(G902), .ZN(n381) );
  BUF_X1 U412 ( .A(n497), .Z(n510) );
  INV_X1 U413 ( .A(KEYINPUT70), .ZN(n577) );
  XNOR2_X1 U414 ( .A(n520), .B(n516), .ZN(n517) );
  XNOR2_X1 U415 ( .A(n577), .B(KEYINPUT48), .ZN(n578) );
  NAND2_X1 U416 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U417 ( .A(n429), .B(n415), .ZN(n606) );
  BUF_X1 U418 ( .A(n545), .Z(n672) );
  XNOR2_X1 U419 ( .A(n472), .B(n471), .ZN(n503) );
  BUF_X1 U420 ( .A(n464), .Z(n541) );
  INV_X1 U421 ( .A(KEYINPUT109), .ZN(n561) );
  XNOR2_X1 U422 ( .A(n562), .B(n561), .ZN(n727) );
  INV_X1 U423 ( .A(G475), .ZN(n369) );
  XNOR2_X2 U424 ( .A(G146), .B(G125), .ZN(n390) );
  XNOR2_X1 U425 ( .A(G140), .B(KEYINPUT10), .ZN(n357) );
  INV_X1 U426 ( .A(G113), .ZN(n358) );
  XNOR2_X1 U427 ( .A(n358), .B(G104), .ZN(n387) );
  NAND2_X1 U428 ( .A1(n409), .A2(G214), .ZN(n359) );
  XNOR2_X1 U429 ( .A(n387), .B(n359), .ZN(n360) );
  XNOR2_X1 U430 ( .A(n717), .B(n360), .ZN(n365) );
  XOR2_X1 U431 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n362) );
  XNOR2_X1 U432 ( .A(G143), .B(G122), .ZN(n361) );
  XNOR2_X1 U433 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U434 ( .A(KEYINPUT69), .B(G131), .ZN(n406) );
  XNOR2_X1 U435 ( .A(n363), .B(n406), .ZN(n364) );
  XNOR2_X1 U436 ( .A(n365), .B(n364), .ZN(n614) );
  NOR2_X1 U437 ( .A1(G902), .A2(n614), .ZN(n367) );
  XNOR2_X1 U438 ( .A(KEYINPUT13), .B(KEYINPUT101), .ZN(n366) );
  XNOR2_X1 U439 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X2 U440 ( .A(G143), .B(KEYINPUT82), .ZN(n370) );
  XNOR2_X2 U441 ( .A(n370), .B(G128), .ZN(n391) );
  XOR2_X1 U442 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n373) );
  INV_X2 U443 ( .A(G953), .ZN(n722) );
  NAND2_X1 U444 ( .A1(G234), .A2(n722), .ZN(n372) );
  XNOR2_X1 U445 ( .A(n373), .B(n372), .ZN(n438) );
  NAND2_X1 U446 ( .A1(G217), .A2(n438), .ZN(n377) );
  XOR2_X1 U447 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n375) );
  XNOR2_X1 U448 ( .A(G116), .B(KEYINPUT103), .ZN(n374) );
  XNOR2_X1 U449 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U450 ( .A(n377), .B(n376), .ZN(n379) );
  XNOR2_X2 U451 ( .A(G122), .B(G107), .ZN(n386) );
  XOR2_X1 U452 ( .A(KEYINPUT9), .B(n386), .Z(n378) );
  XNOR2_X1 U453 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U454 ( .A(n408), .B(n380), .ZN(n627) );
  NAND2_X1 U455 ( .A1(n486), .A2(n487), .ZN(n382) );
  XNOR2_X1 U456 ( .A(n382), .B(KEYINPUT106), .ZN(n505) );
  XNOR2_X1 U457 ( .A(n383), .B(KEYINPUT3), .ZN(n385) );
  XNOR2_X1 U458 ( .A(G101), .B(KEYINPUT73), .ZN(n384) );
  XNOR2_X1 U459 ( .A(n385), .B(n384), .ZN(n414) );
  XNOR2_X1 U460 ( .A(n386), .B(KEYINPUT16), .ZN(n388) );
  XNOR2_X1 U461 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U462 ( .A(n414), .B(n389), .ZN(n711) );
  XNOR2_X1 U463 ( .A(KEYINPUT75), .B(G110), .ZN(n422) );
  XNOR2_X1 U464 ( .A(n390), .B(n422), .ZN(n392) );
  XNOR2_X1 U465 ( .A(n392), .B(n391), .ZN(n400) );
  XNOR2_X1 U466 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n394) );
  NAND2_X1 U467 ( .A1(n722), .A2(G224), .ZN(n393) );
  XNOR2_X1 U468 ( .A(n394), .B(n393), .ZN(n398) );
  XNOR2_X1 U469 ( .A(KEYINPUT18), .B(KEYINPUT81), .ZN(n396) );
  XNOR2_X1 U470 ( .A(KEYINPUT91), .B(KEYINPUT93), .ZN(n395) );
  XNOR2_X1 U471 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U472 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U473 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U474 ( .A(n711), .B(n401), .ZN(n599) );
  XNOR2_X1 U475 ( .A(KEYINPUT15), .B(G902), .ZN(n432) );
  INV_X1 U476 ( .A(n432), .ZN(n587) );
  OR2_X2 U477 ( .A1(n599), .A2(n587), .ZN(n404) );
  OR2_X1 U478 ( .A1(G237), .A2(G902), .ZN(n402) );
  XNOR2_X1 U479 ( .A(KEYINPUT78), .B(n402), .ZN(n416) );
  NAND2_X1 U480 ( .A1(n416), .A2(G210), .ZN(n403) );
  NOR2_X1 U481 ( .A1(n505), .A2(n541), .ZN(n462) );
  XNOR2_X1 U482 ( .A(KEYINPUT4), .B(G137), .ZN(n405) );
  XNOR2_X1 U483 ( .A(n406), .B(n405), .ZN(n407) );
  NAND2_X1 U484 ( .A1(n409), .A2(G210), .ZN(n410) );
  XNOR2_X1 U485 ( .A(n410), .B(KEYINPUT5), .ZN(n412) );
  XNOR2_X1 U486 ( .A(G113), .B(KEYINPUT79), .ZN(n411) );
  XNOR2_X1 U487 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U488 ( .A(n414), .B(n413), .ZN(n415) );
  NAND2_X1 U489 ( .A1(n416), .A2(G214), .ZN(n418) );
  INV_X1 U490 ( .A(KEYINPUT94), .ZN(n417) );
  XNOR2_X1 U491 ( .A(n418), .B(n417), .ZN(n463) );
  INV_X1 U492 ( .A(n463), .ZN(n681) );
  NAND2_X1 U493 ( .A1(n545), .A2(n681), .ZN(n420) );
  XOR2_X1 U494 ( .A(KEYINPUT30), .B(KEYINPUT108), .Z(n419) );
  XNOR2_X1 U495 ( .A(n420), .B(n419), .ZN(n461) );
  XNOR2_X1 U496 ( .A(G140), .B(KEYINPUT96), .ZN(n421) );
  XNOR2_X1 U497 ( .A(n422), .B(n421), .ZN(n427) );
  XNOR2_X1 U498 ( .A(G101), .B(G104), .ZN(n423) );
  XNOR2_X1 U499 ( .A(G107), .B(n423), .ZN(n425) );
  NAND2_X1 U500 ( .A1(n722), .A2(G227), .ZN(n424) );
  XNOR2_X1 U501 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U502 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U503 ( .A(n429), .B(n428), .ZN(n633) );
  INV_X1 U504 ( .A(G469), .ZN(n430) );
  XNOR2_X2 U505 ( .A(n431), .B(n430), .ZN(n547) );
  NAND2_X1 U506 ( .A1(G234), .A2(n432), .ZN(n433) );
  XNOR2_X1 U507 ( .A(KEYINPUT20), .B(n433), .ZN(n446) );
  NAND2_X1 U508 ( .A1(n446), .A2(G221), .ZN(n434) );
  XNOR2_X1 U509 ( .A(n434), .B(KEYINPUT21), .ZN(n669) );
  XNOR2_X1 U510 ( .A(n669), .B(KEYINPUT98), .ZN(n474) );
  XOR2_X1 U511 ( .A(KEYINPUT74), .B(KEYINPUT24), .Z(n436) );
  XNOR2_X1 U512 ( .A(KEYINPUT97), .B(KEYINPUT23), .ZN(n435) );
  XNOR2_X1 U513 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U514 ( .A(n717), .B(n437), .ZN(n444) );
  NAND2_X1 U515 ( .A1(n438), .A2(G221), .ZN(n442) );
  XOR2_X1 U516 ( .A(G110), .B(G128), .Z(n440) );
  XNOR2_X1 U517 ( .A(G119), .B(G137), .ZN(n439) );
  XNOR2_X1 U518 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U519 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U520 ( .A(n444), .B(n443), .ZN(n622) );
  INV_X1 U521 ( .A(G902), .ZN(n445) );
  NAND2_X1 U522 ( .A1(n622), .A2(n445), .ZN(n450) );
  NAND2_X1 U523 ( .A1(n446), .A2(G217), .ZN(n448) );
  XNOR2_X1 U524 ( .A(KEYINPUT25), .B(KEYINPUT80), .ZN(n447) );
  XNOR2_X1 U525 ( .A(n448), .B(n447), .ZN(n449) );
  OR2_X1 U526 ( .A1(n474), .A2(n668), .ZN(n663) );
  XOR2_X1 U527 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n452) );
  NAND2_X1 U528 ( .A1(G234), .A2(G237), .ZN(n451) );
  XNOR2_X1 U529 ( .A(n452), .B(n451), .ZN(n456) );
  NAND2_X1 U530 ( .A1(G952), .A2(n456), .ZN(n697) );
  NOR2_X1 U531 ( .A1(G953), .A2(n697), .ZN(n454) );
  INV_X1 U532 ( .A(KEYINPUT95), .ZN(n453) );
  XNOR2_X1 U533 ( .A(n454), .B(n453), .ZN(n468) );
  AND2_X1 U534 ( .A1(G953), .A2(G902), .ZN(n455) );
  NAND2_X1 U535 ( .A1(n456), .A2(n455), .ZN(n466) );
  XOR2_X1 U536 ( .A(n466), .B(KEYINPUT107), .Z(n457) );
  NOR2_X1 U537 ( .A1(G900), .A2(n457), .ZN(n458) );
  OR2_X1 U538 ( .A1(n468), .A2(n458), .ZN(n482) );
  NAND2_X1 U539 ( .A1(n498), .A2(n482), .ZN(n459) );
  NOR2_X1 U540 ( .A1(n547), .A2(n459), .ZN(n460) );
  AND2_X1 U541 ( .A1(n461), .A2(n460), .ZN(n550) );
  NAND2_X1 U542 ( .A1(n462), .A2(n550), .ZN(n564) );
  XNOR2_X1 U543 ( .A(n564), .B(G143), .ZN(G45) );
  OR2_X2 U544 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X2 U545 ( .A(n465), .B(KEYINPUT19), .ZN(n566) );
  NOR2_X1 U546 ( .A1(n466), .A2(G898), .ZN(n467) );
  OR2_X1 U547 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U548 ( .A1(n566), .A2(n469), .ZN(n472) );
  INV_X1 U549 ( .A(KEYINPUT90), .ZN(n470) );
  XNOR2_X1 U550 ( .A(n470), .B(KEYINPUT0), .ZN(n471) );
  NOR2_X1 U551 ( .A1(n487), .A2(n486), .ZN(n473) );
  XNOR2_X1 U552 ( .A(KEYINPUT105), .B(n473), .ZN(n685) );
  NOR2_X1 U553 ( .A1(n474), .A2(n685), .ZN(n475) );
  NAND2_X1 U554 ( .A1(n503), .A2(n475), .ZN(n477) );
  XOR2_X1 U555 ( .A(KEYINPUT76), .B(KEYINPUT22), .Z(n476) );
  XNOR2_X2 U556 ( .A(n477), .B(n476), .ZN(n513) );
  INV_X1 U557 ( .A(n513), .ZN(n481) );
  NOR2_X1 U558 ( .A1(n350), .A2(n668), .ZN(n479) );
  XNOR2_X1 U559 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n478) );
  XNOR2_X2 U560 ( .A(n547), .B(n478), .ZN(n664) );
  NAND2_X1 U561 ( .A1(n479), .A2(n664), .ZN(n480) );
  NOR2_X1 U562 ( .A1(n481), .A2(n480), .ZN(n534) );
  XOR2_X1 U563 ( .A(G101), .B(n534), .Z(G3) );
  XNOR2_X1 U564 ( .A(G140), .B(KEYINPUT116), .ZN(n492) );
  INV_X1 U565 ( .A(n482), .ZN(n483) );
  NOR2_X1 U566 ( .A1(n483), .A2(n669), .ZN(n484) );
  XNOR2_X1 U567 ( .A(n484), .B(KEYINPUT72), .ZN(n485) );
  NAND2_X1 U568 ( .A1(n668), .A2(n485), .ZN(n543) );
  XNOR2_X1 U569 ( .A(n486), .B(KEYINPUT102), .ZN(n530) );
  INV_X1 U570 ( .A(n487), .ZN(n531) );
  NAND2_X1 U571 ( .A1(n530), .A2(n531), .ZN(n532) );
  NOR2_X1 U572 ( .A1(n543), .A2(n532), .ZN(n488) );
  NAND2_X1 U573 ( .A1(n681), .A2(n488), .ZN(n489) );
  NOR2_X2 U574 ( .A1(n510), .A2(n489), .ZN(n556) );
  NAND2_X1 U575 ( .A1(n556), .A2(n664), .ZN(n490) );
  XOR2_X1 U576 ( .A(KEYINPUT43), .B(n490), .Z(n491) );
  INV_X1 U577 ( .A(n541), .ZN(n555) );
  NOR2_X1 U578 ( .A1(n491), .A2(n555), .ZN(n580) );
  XOR2_X1 U579 ( .A(n492), .B(n580), .Z(G42) );
  INV_X1 U580 ( .A(n664), .ZN(n559) );
  NOR2_X1 U581 ( .A1(n559), .A2(n672), .ZN(n493) );
  NAND2_X1 U582 ( .A1(n513), .A2(n493), .ZN(n494) );
  XOR2_X1 U583 ( .A(KEYINPUT65), .B(n494), .Z(n496) );
  INV_X1 U584 ( .A(n668), .ZN(n495) );
  NOR2_X2 U585 ( .A1(n496), .A2(n495), .ZN(n515) );
  XOR2_X1 U586 ( .A(n515), .B(G110), .Z(G12) );
  XNOR2_X1 U587 ( .A(n502), .B(n501), .ZN(n690) );
  NAND2_X1 U588 ( .A1(n690), .A2(n528), .ZN(n504) );
  XNOR2_X1 U589 ( .A(n504), .B(KEYINPUT34), .ZN(n506) );
  XOR2_X1 U590 ( .A(KEYINPUT86), .B(KEYINPUT35), .Z(n507) );
  XNOR2_X1 U591 ( .A(n509), .B(KEYINPUT67), .ZN(n518) );
  NAND2_X1 U592 ( .A1(n510), .A2(n668), .ZN(n511) );
  NOR2_X1 U593 ( .A1(n511), .A2(n664), .ZN(n512) );
  NAND2_X1 U594 ( .A1(n513), .A2(n512), .ZN(n514) );
  XOR2_X1 U595 ( .A(KEYINPUT32), .B(n514), .Z(n728) );
  NOR2_X1 U596 ( .A1(n518), .A2(n517), .ZN(n539) );
  INV_X1 U597 ( .A(n620), .ZN(n519) );
  NAND2_X1 U598 ( .A1(n520), .A2(n519), .ZN(n521) );
  NAND2_X1 U599 ( .A1(n521), .A2(KEYINPUT44), .ZN(n537) );
  NAND2_X1 U600 ( .A1(n672), .A2(n498), .ZN(n522) );
  NOR2_X1 U601 ( .A1(n664), .A2(n522), .ZN(n677) );
  NAND2_X1 U602 ( .A1(n677), .A2(n528), .ZN(n524) );
  XNOR2_X1 U603 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n523) );
  XNOR2_X1 U604 ( .A(n524), .B(n523), .ZN(n655) );
  INV_X1 U605 ( .A(n672), .ZN(n525) );
  NAND2_X1 U606 ( .A1(n525), .A2(n498), .ZN(n526) );
  NOR2_X1 U607 ( .A1(n526), .A2(n547), .ZN(n527) );
  NAND2_X1 U608 ( .A1(n528), .A2(n527), .ZN(n640) );
  NAND2_X1 U609 ( .A1(n655), .A2(n640), .ZN(n529) );
  XOR2_X1 U610 ( .A(KEYINPUT100), .B(n529), .Z(n533) );
  NOR2_X1 U611 ( .A1(n531), .A2(n530), .ZN(n646) );
  INV_X1 U612 ( .A(n653), .ZN(n650) );
  NOR2_X1 U613 ( .A1(n533), .A2(n687), .ZN(n535) );
  NOR2_X1 U614 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U615 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U616 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U617 ( .A(n540), .B(KEYINPUT45), .ZN(n592) );
  INV_X1 U618 ( .A(n592), .ZN(n584) );
  XNOR2_X1 U619 ( .A(n541), .B(KEYINPUT38), .ZN(n682) );
  NAND2_X1 U620 ( .A1(n682), .A2(n681), .ZN(n686) );
  NOR2_X1 U621 ( .A1(n685), .A2(n686), .ZN(n542) );
  XNOR2_X1 U622 ( .A(n542), .B(KEYINPUT41), .ZN(n699) );
  INV_X1 U623 ( .A(n543), .ZN(n544) );
  NAND2_X1 U624 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U625 ( .A(n546), .B(KEYINPUT28), .ZN(n548) );
  NOR2_X1 U626 ( .A1(n699), .A2(n568), .ZN(n549) );
  XNOR2_X1 U627 ( .A(n549), .B(KEYINPUT42), .ZN(n730) );
  NAND2_X1 U628 ( .A1(n550), .A2(n682), .ZN(n551) );
  XNOR2_X1 U629 ( .A(n551), .B(KEYINPUT39), .ZN(n582) );
  AND2_X1 U630 ( .A1(n582), .A2(n650), .ZN(n552) );
  XNOR2_X1 U631 ( .A(n552), .B(KEYINPUT40), .ZN(n729) );
  NOR2_X1 U632 ( .A1(n730), .A2(n729), .ZN(n554) );
  XNOR2_X1 U633 ( .A(KEYINPUT87), .B(KEYINPUT46), .ZN(n553) );
  XNOR2_X1 U634 ( .A(n554), .B(n553), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n556), .A2(n555), .ZN(n558) );
  XNOR2_X1 U636 ( .A(KEYINPUT36), .B(KEYINPUT89), .ZN(n557) );
  XNOR2_X1 U637 ( .A(n558), .B(n557), .ZN(n560) );
  NAND2_X1 U638 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U639 ( .A1(n687), .A2(KEYINPUT47), .ZN(n563) );
  NAND2_X1 U640 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U641 ( .A(n565), .B(KEYINPUT84), .ZN(n572) );
  INV_X1 U642 ( .A(n566), .ZN(n567) );
  NAND2_X1 U643 ( .A1(n651), .A2(n687), .ZN(n569) );
  AND2_X1 U644 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U645 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U646 ( .A(n574), .B(KEYINPUT71), .ZN(n575) );
  NOR2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n579) );
  XNOR2_X1 U648 ( .A(n579), .B(n578), .ZN(n581) );
  NAND2_X1 U649 ( .A1(n582), .A2(n646), .ZN(n658) );
  NAND2_X1 U650 ( .A1(n353), .A2(n351), .ZN(n720) );
  INV_X1 U651 ( .A(n720), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n586) );
  INV_X1 U653 ( .A(KEYINPUT2), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n659), .A2(n587), .ZN(n588) );
  XNOR2_X1 U655 ( .A(n588), .B(KEYINPUT64), .ZN(n595) );
  NAND2_X1 U656 ( .A1(n658), .A2(KEYINPUT2), .ZN(n590) );
  XNOR2_X1 U657 ( .A(n590), .B(KEYINPUT83), .ZN(n591) );
  NAND2_X1 U658 ( .A1(n589), .A2(n591), .ZN(n594) );
  BUF_X1 U659 ( .A(n592), .Z(n593) );
  NOR2_X1 U660 ( .A1(n594), .A2(n593), .ZN(n660) );
  NOR2_X2 U661 ( .A1(n595), .A2(n660), .ZN(n621) );
  NAND2_X1 U662 ( .A1(n621), .A2(G210), .ZN(n601) );
  XOR2_X1 U663 ( .A(KEYINPUT124), .B(KEYINPUT54), .Z(n597) );
  XNOR2_X1 U664 ( .A(KEYINPUT55), .B(KEYINPUT85), .ZN(n596) );
  XNOR2_X1 U665 ( .A(n597), .B(n596), .ZN(n598) );
  XNOR2_X1 U666 ( .A(n599), .B(n598), .ZN(n600) );
  XNOR2_X1 U667 ( .A(n601), .B(n600), .ZN(n603) );
  INV_X1 U668 ( .A(G952), .ZN(n602) );
  NAND2_X1 U669 ( .A1(n602), .A2(G953), .ZN(n625) );
  NAND2_X1 U670 ( .A1(n603), .A2(n625), .ZN(n605) );
  INV_X1 U671 ( .A(KEYINPUT56), .ZN(n604) );
  XNOR2_X1 U672 ( .A(n605), .B(n604), .ZN(G51) );
  NAND2_X1 U673 ( .A1(n621), .A2(G472), .ZN(n609) );
  XOR2_X1 U674 ( .A(KEYINPUT110), .B(KEYINPUT62), .Z(n607) );
  XNOR2_X1 U675 ( .A(n606), .B(n607), .ZN(n608) );
  XNOR2_X1 U676 ( .A(n609), .B(n608), .ZN(n610) );
  NAND2_X1 U677 ( .A1(n610), .A2(n625), .ZN(n612) );
  XOR2_X1 U678 ( .A(KEYINPUT111), .B(KEYINPUT63), .Z(n611) );
  XNOR2_X1 U679 ( .A(n612), .B(n611), .ZN(G57) );
  NAND2_X1 U680 ( .A1(n621), .A2(G475), .ZN(n616) );
  XNOR2_X1 U681 ( .A(KEYINPUT92), .B(KEYINPUT59), .ZN(n613) );
  XNOR2_X1 U682 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U683 ( .A(n616), .B(n615), .ZN(n617) );
  NAND2_X1 U684 ( .A1(n617), .A2(n625), .ZN(n619) );
  INV_X1 U685 ( .A(KEYINPUT60), .ZN(n618) );
  XNOR2_X1 U686 ( .A(n619), .B(n618), .ZN(G60) );
  XOR2_X1 U687 ( .A(n354), .B(G122), .Z(G24) );
  NAND2_X1 U688 ( .A1(n631), .A2(G217), .ZN(n624) );
  XOR2_X1 U689 ( .A(KEYINPUT126), .B(n622), .Z(n623) );
  XNOR2_X1 U690 ( .A(n624), .B(n623), .ZN(n626) );
  INV_X1 U691 ( .A(n625), .ZN(n636) );
  NOR2_X1 U692 ( .A1(n626), .A2(n636), .ZN(G66) );
  NAND2_X1 U693 ( .A1(n631), .A2(G478), .ZN(n629) );
  XOR2_X1 U694 ( .A(KEYINPUT125), .B(n627), .Z(n628) );
  XNOR2_X1 U695 ( .A(n629), .B(n628), .ZN(n630) );
  NOR2_X1 U696 ( .A1(n630), .A2(n636), .ZN(G63) );
  NAND2_X1 U697 ( .A1(n631), .A2(G469), .ZN(n635) );
  XOR2_X1 U698 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n632) );
  XNOR2_X1 U699 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U700 ( .A(n635), .B(n634), .ZN(n637) );
  NOR2_X1 U701 ( .A1(n637), .A2(n636), .ZN(G54) );
  NOR2_X1 U702 ( .A1(n640), .A2(n653), .ZN(n638) );
  XOR2_X1 U703 ( .A(KEYINPUT112), .B(n638), .Z(n639) );
  XNOR2_X1 U704 ( .A(G104), .B(n639), .ZN(G6) );
  INV_X1 U705 ( .A(n646), .ZN(n656) );
  NOR2_X1 U706 ( .A1(n640), .A2(n656), .ZN(n645) );
  XOR2_X1 U707 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n642) );
  XNOR2_X1 U708 ( .A(G107), .B(KEYINPUT26), .ZN(n641) );
  XNOR2_X1 U709 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U710 ( .A(KEYINPUT27), .B(n643), .ZN(n644) );
  XNOR2_X1 U711 ( .A(n645), .B(n644), .ZN(G9) );
  XOR2_X1 U712 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n648) );
  NAND2_X1 U713 ( .A1(n651), .A2(n646), .ZN(n647) );
  XNOR2_X1 U714 ( .A(n648), .B(n647), .ZN(n649) );
  XOR2_X1 U715 ( .A(G128), .B(n649), .Z(G30) );
  NAND2_X1 U716 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U717 ( .A(n652), .B(G146), .ZN(G48) );
  NOR2_X1 U718 ( .A1(n653), .A2(n655), .ZN(n654) );
  XOR2_X1 U719 ( .A(G113), .B(n654), .Z(G15) );
  NOR2_X1 U720 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U721 ( .A(G116), .B(n657), .Z(G18) );
  XNOR2_X1 U722 ( .A(G134), .B(n658), .ZN(G36) );
  INV_X1 U723 ( .A(n659), .ZN(n661) );
  NOR2_X1 U724 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U725 ( .A1(n662), .A2(G953), .ZN(n704) );
  NAND2_X1 U726 ( .A1(n664), .A2(n663), .ZN(n667) );
  XNOR2_X1 U727 ( .A(KEYINPUT119), .B(KEYINPUT50), .ZN(n665) );
  XOR2_X1 U728 ( .A(n665), .B(KEYINPUT118), .Z(n666) );
  XNOR2_X1 U729 ( .A(n667), .B(n666), .ZN(n675) );
  XOR2_X1 U730 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n671) );
  NAND2_X1 U731 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U732 ( .A(n671), .B(n670), .ZN(n673) );
  NOR2_X1 U733 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U734 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U735 ( .A(KEYINPUT120), .B(n676), .Z(n678) );
  NOR2_X1 U736 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U737 ( .A(KEYINPUT51), .B(n679), .Z(n680) );
  NOR2_X1 U738 ( .A1(n699), .A2(n680), .ZN(n693) );
  NOR2_X1 U739 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U740 ( .A(KEYINPUT121), .B(n683), .Z(n684) );
  NOR2_X1 U741 ( .A1(n685), .A2(n684), .ZN(n689) );
  NOR2_X1 U742 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U743 ( .A1(n689), .A2(n688), .ZN(n691) );
  INV_X1 U744 ( .A(n690), .ZN(n698) );
  NOR2_X1 U745 ( .A1(n691), .A2(n698), .ZN(n692) );
  NOR2_X1 U746 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U747 ( .A(n694), .B(KEYINPUT52), .ZN(n695) );
  XNOR2_X1 U748 ( .A(KEYINPUT122), .B(n695), .ZN(n696) );
  NOR2_X1 U749 ( .A1(n697), .A2(n696), .ZN(n701) );
  NOR2_X1 U750 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U751 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U752 ( .A(KEYINPUT123), .B(n702), .Z(n703) );
  NAND2_X1 U753 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U754 ( .A(KEYINPUT53), .B(n705), .Z(G75) );
  NOR2_X1 U755 ( .A1(n593), .A2(G953), .ZN(n710) );
  NAND2_X1 U756 ( .A1(G953), .A2(G224), .ZN(n706) );
  XNOR2_X1 U757 ( .A(KEYINPUT61), .B(n706), .ZN(n707) );
  NAND2_X1 U758 ( .A1(n707), .A2(G898), .ZN(n708) );
  XNOR2_X1 U759 ( .A(n708), .B(KEYINPUT127), .ZN(n709) );
  NOR2_X1 U760 ( .A1(n710), .A2(n709), .ZN(n715) );
  XNOR2_X1 U761 ( .A(n711), .B(G110), .ZN(n713) );
  NOR2_X1 U762 ( .A1(n722), .A2(G898), .ZN(n712) );
  NOR2_X1 U763 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U764 ( .A(n715), .B(n714), .Z(G69) );
  XOR2_X1 U765 ( .A(n716), .B(n717), .Z(n721) );
  XNOR2_X1 U766 ( .A(n721), .B(G227), .ZN(n718) );
  NAND2_X1 U767 ( .A1(G900), .A2(n718), .ZN(n719) );
  NAND2_X1 U768 ( .A1(n719), .A2(G953), .ZN(n725) );
  XNOR2_X1 U769 ( .A(n720), .B(n721), .ZN(n723) );
  NAND2_X1 U770 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U771 ( .A1(n725), .A2(n724), .ZN(G72) );
  XOR2_X1 U772 ( .A(G125), .B(KEYINPUT37), .Z(n726) );
  XNOR2_X1 U773 ( .A(n727), .B(n726), .ZN(G27) );
  XOR2_X1 U774 ( .A(G119), .B(n728), .Z(G21) );
  XOR2_X1 U775 ( .A(n729), .B(G131), .Z(G33) );
  XOR2_X1 U776 ( .A(G137), .B(n730), .Z(G39) );
endmodule

