

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U553 ( .A(n533), .B(KEYINPUT65), .ZN(n597) );
  NOR2_X2 U554 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X2 U555 ( .A(n612), .B(n611), .ZN(n615) );
  NOR2_X2 U556 ( .A1(n597), .A2(n598), .ZN(n521) );
  NAND2_X1 U557 ( .A1(n759), .A2(n758), .ZN(n761) );
  NOR2_X1 U558 ( .A1(n608), .A2(n606), .ZN(G160) );
  NOR2_X1 U559 ( .A1(n701), .A2(n700), .ZN(n520) );
  INV_X1 U560 ( .A(KEYINPUT26), .ZN(n627) );
  NOR2_X1 U561 ( .A1(n609), .A2(n725), .ZN(n610) );
  INV_X1 U562 ( .A(KEYINPUT93), .ZN(n636) );
  XNOR2_X1 U563 ( .A(n637), .B(n636), .ZN(n645) );
  INV_X1 U564 ( .A(KEYINPUT95), .ZN(n668) );
  INV_X1 U565 ( .A(G2104), .ZN(n533) );
  NOR2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n539) );
  NOR2_X1 U567 ( .A1(G543), .A2(n526), .ZN(n522) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n795) );
  INV_X1 U569 ( .A(KEYINPUT40), .ZN(n760) );
  BUF_X1 U570 ( .A(n762), .Z(G164) );
  XNOR2_X1 U571 ( .A(G651), .B(KEYINPUT67), .ZN(n526) );
  XOR2_X1 U572 ( .A(KEYINPUT1), .B(n522), .Z(n791) );
  NAND2_X1 U573 ( .A1(G62), .A2(n791), .ZN(n525) );
  XOR2_X1 U574 ( .A(KEYINPUT0), .B(G543), .Z(n575) );
  NOR2_X1 U575 ( .A1(G651), .A2(n575), .ZN(n523) );
  XNOR2_X1 U576 ( .A(KEYINPUT64), .B(n523), .ZN(n792) );
  NAND2_X1 U577 ( .A1(G50), .A2(n792), .ZN(n524) );
  NAND2_X1 U578 ( .A1(n525), .A2(n524), .ZN(n532) );
  NAND2_X1 U579 ( .A1(G88), .A2(n795), .ZN(n529) );
  NOR2_X1 U580 ( .A1(n575), .A2(n526), .ZN(n527) );
  XNOR2_X1 U581 ( .A(KEYINPUT68), .B(n527), .ZN(n789) );
  NAND2_X1 U582 ( .A1(G75), .A2(n789), .ZN(n528) );
  NAND2_X1 U583 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U584 ( .A(KEYINPUT83), .B(n530), .Z(n531) );
  NOR2_X1 U585 ( .A1(n532), .A2(n531), .ZN(G166) );
  INV_X1 U586 ( .A(G2105), .ZN(n598) );
  AND2_X1 U587 ( .A1(n598), .A2(G101), .ZN(n534) );
  NAND2_X1 U588 ( .A1(n597), .A2(n534), .ZN(n535) );
  XOR2_X1 U589 ( .A(n535), .B(KEYINPUT23), .Z(n537) );
  NAND2_X1 U590 ( .A1(n521), .A2(G125), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U592 ( .A(n538), .B(KEYINPUT66), .ZN(n608) );
  XOR2_X2 U593 ( .A(KEYINPUT17), .B(n539), .Z(n877) );
  NAND2_X1 U594 ( .A1(G137), .A2(n877), .ZN(n541) );
  AND2_X1 U595 ( .A1(G2105), .A2(G2104), .ZN(n874) );
  NAND2_X1 U596 ( .A1(G113), .A2(n874), .ZN(n540) );
  NAND2_X1 U597 ( .A1(n541), .A2(n540), .ZN(n606) );
  NAND2_X1 U598 ( .A1(n789), .A2(G78), .ZN(n542) );
  XOR2_X1 U599 ( .A(KEYINPUT70), .B(n542), .Z(n547) );
  NAND2_X1 U600 ( .A1(G65), .A2(n791), .ZN(n544) );
  NAND2_X1 U601 ( .A1(G53), .A2(n792), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U603 ( .A(KEYINPUT71), .B(n545), .Z(n546) );
  NOR2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n795), .A2(G91), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(G299) );
  NAND2_X1 U607 ( .A1(G90), .A2(n795), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G77), .A2(n789), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U610 ( .A(KEYINPUT9), .B(n552), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n792), .A2(G52), .ZN(n554) );
  NAND2_X1 U612 ( .A1(G64), .A2(n791), .ZN(n553) );
  AND2_X1 U613 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n556), .A2(n555), .ZN(G301) );
  NAND2_X1 U615 ( .A1(n795), .A2(G89), .ZN(n557) );
  XNOR2_X1 U616 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U617 ( .A1(G76), .A2(n789), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U619 ( .A(n560), .B(KEYINPUT5), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G63), .A2(n791), .ZN(n562) );
  NAND2_X1 U621 ( .A1(G51), .A2(n792), .ZN(n561) );
  NAND2_X1 U622 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U623 ( .A(KEYINPUT6), .B(n563), .Z(n564) );
  NAND2_X1 U624 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U625 ( .A(n566), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U626 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U627 ( .A(G166), .ZN(G303) );
  NAND2_X1 U628 ( .A1(n792), .A2(G48), .ZN(n573) );
  NAND2_X1 U629 ( .A1(G86), .A2(n795), .ZN(n568) );
  NAND2_X1 U630 ( .A1(G61), .A2(n791), .ZN(n567) );
  NAND2_X1 U631 ( .A1(n568), .A2(n567), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n789), .A2(G73), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT2), .B(n569), .Z(n570) );
  NOR2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U636 ( .A(n574), .B(KEYINPUT82), .ZN(G305) );
  NAND2_X1 U637 ( .A1(G87), .A2(n575), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G74), .A2(G651), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U640 ( .A1(n791), .A2(n578), .ZN(n580) );
  NAND2_X1 U641 ( .A1(G49), .A2(n792), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n580), .A2(n579), .ZN(G288) );
  NAND2_X1 U643 ( .A1(G72), .A2(n789), .ZN(n582) );
  NAND2_X1 U644 ( .A1(n795), .A2(G85), .ZN(n581) );
  NAND2_X1 U645 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT69), .B(n583), .ZN(n587) );
  NAND2_X1 U647 ( .A1(n792), .A2(G47), .ZN(n585) );
  NAND2_X1 U648 ( .A1(G60), .A2(n791), .ZN(n584) );
  AND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U650 ( .A1(n587), .A2(n586), .ZN(G290) );
  NAND2_X1 U651 ( .A1(G8), .A2(G166), .ZN(n588) );
  NOR2_X1 U652 ( .A1(G2090), .A2(n588), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n589), .B(KEYINPUT97), .ZN(n687) );
  NAND2_X1 U654 ( .A1(G79), .A2(n789), .ZN(n591) );
  NAND2_X1 U655 ( .A1(G54), .A2(n792), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U657 ( .A1(G66), .A2(n791), .ZN(n593) );
  NAND2_X1 U658 ( .A1(G92), .A2(n795), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U660 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U661 ( .A(KEYINPUT15), .B(n596), .Z(n1008) );
  AND2_X1 U662 ( .A1(n598), .A2(n597), .ZN(n709) );
  NAND2_X1 U663 ( .A1(G102), .A2(n709), .ZN(n600) );
  NAND2_X1 U664 ( .A1(G114), .A2(n874), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U666 ( .A1(G138), .A2(n877), .ZN(n602) );
  NAND2_X1 U667 ( .A1(G126), .A2(n521), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U669 ( .A1(n604), .A2(n603), .ZN(n762) );
  NOR2_X2 U670 ( .A1(n762), .A2(G1384), .ZN(n726) );
  INV_X1 U671 ( .A(n726), .ZN(n609) );
  INV_X1 U672 ( .A(G40), .ZN(n605) );
  OR2_X1 U673 ( .A1(n606), .A2(n605), .ZN(n607) );
  OR2_X1 U674 ( .A1(n608), .A2(n607), .ZN(n725) );
  XNOR2_X1 U675 ( .A(n610), .B(KEYINPUT88), .ZN(n640) );
  NAND2_X1 U676 ( .A1(G2067), .A2(n640), .ZN(n612) );
  INV_X1 U677 ( .A(KEYINPUT92), .ZN(n611) );
  AND2_X1 U678 ( .A1(n726), .A2(G40), .ZN(n613) );
  NAND2_X1 U679 ( .A1(n613), .A2(G160), .ZN(n671) );
  INV_X1 U680 ( .A(n671), .ZN(n653) );
  INV_X1 U681 ( .A(G1348), .ZN(n977) );
  NOR2_X1 U682 ( .A1(n653), .A2(n977), .ZN(n614) );
  OR2_X1 U683 ( .A1(n1008), .A2(n616), .ZN(n635) );
  NAND2_X1 U684 ( .A1(n1008), .A2(n616), .ZN(n633) );
  NAND2_X1 U685 ( .A1(G56), .A2(n791), .ZN(n617) );
  XOR2_X1 U686 ( .A(KEYINPUT14), .B(n617), .Z(n624) );
  NAND2_X1 U687 ( .A1(G81), .A2(n795), .ZN(n618) );
  XNOR2_X1 U688 ( .A(n618), .B(KEYINPUT72), .ZN(n619) );
  XNOR2_X1 U689 ( .A(n619), .B(KEYINPUT12), .ZN(n621) );
  NAND2_X1 U690 ( .A1(G68), .A2(n789), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U692 ( .A(KEYINPUT13), .B(n622), .Z(n623) );
  NOR2_X1 U693 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U694 ( .A1(G43), .A2(n792), .ZN(n625) );
  NAND2_X1 U695 ( .A1(n626), .A2(n625), .ZN(n1027) );
  INV_X1 U696 ( .A(G1996), .ZN(n829) );
  NOR2_X1 U697 ( .A1(n671), .A2(n829), .ZN(n628) );
  XNOR2_X1 U698 ( .A(n628), .B(n627), .ZN(n630) );
  NAND2_X1 U699 ( .A1(n671), .A2(G1341), .ZN(n629) );
  NAND2_X1 U700 ( .A1(n630), .A2(n629), .ZN(n631) );
  OR2_X1 U701 ( .A1(n1027), .A2(n631), .ZN(n632) );
  NAND2_X1 U702 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n635), .A2(n634), .ZN(n637) );
  XOR2_X1 U704 ( .A(KEYINPUT27), .B(KEYINPUT89), .Z(n639) );
  NAND2_X1 U705 ( .A1(G2072), .A2(n640), .ZN(n638) );
  XNOR2_X1 U706 ( .A(n639), .B(n638), .ZN(n643) );
  INV_X1 U707 ( .A(n640), .ZN(n652) );
  NAND2_X1 U708 ( .A1(n652), .A2(G1956), .ZN(n641) );
  XOR2_X1 U709 ( .A(KEYINPUT90), .B(n641), .Z(n642) );
  NOR2_X1 U710 ( .A1(n643), .A2(n642), .ZN(n646) );
  INV_X1 U711 ( .A(G299), .ZN(n1010) );
  NAND2_X1 U712 ( .A1(n646), .A2(n1010), .ZN(n644) );
  NAND2_X1 U713 ( .A1(n645), .A2(n644), .ZN(n650) );
  NOR2_X1 U714 ( .A1(n646), .A2(n1010), .ZN(n648) );
  XNOR2_X1 U715 ( .A(KEYINPUT28), .B(KEYINPUT91), .ZN(n647) );
  XNOR2_X1 U716 ( .A(n648), .B(n647), .ZN(n649) );
  NAND2_X1 U717 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U718 ( .A(n651), .B(KEYINPUT29), .ZN(n657) );
  XOR2_X1 U719 ( .A(G2078), .B(KEYINPUT25), .Z(n934) );
  NOR2_X1 U720 ( .A1(n934), .A2(n652), .ZN(n655) );
  NOR2_X1 U721 ( .A1(n653), .A2(G1961), .ZN(n654) );
  NOR2_X1 U722 ( .A1(n655), .A2(n654), .ZN(n658) );
  NOR2_X1 U723 ( .A1(G301), .A2(n658), .ZN(n656) );
  NOR2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n667) );
  AND2_X1 U725 ( .A1(G301), .A2(n658), .ZN(n663) );
  NAND2_X1 U726 ( .A1(G8), .A2(n671), .ZN(n700) );
  NOR2_X1 U727 ( .A1(G1966), .A2(n700), .ZN(n681) );
  NOR2_X1 U728 ( .A1(G2084), .A2(n671), .ZN(n679) );
  NOR2_X1 U729 ( .A1(n681), .A2(n679), .ZN(n659) );
  NAND2_X1 U730 ( .A1(G8), .A2(n659), .ZN(n660) );
  XNOR2_X1 U731 ( .A(KEYINPUT30), .B(n660), .ZN(n661) );
  NOR2_X1 U732 ( .A1(G168), .A2(n661), .ZN(n662) );
  NOR2_X1 U733 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U734 ( .A(KEYINPUT31), .B(n664), .ZN(n665) );
  XNOR2_X1 U735 ( .A(KEYINPUT94), .B(n665), .ZN(n666) );
  NOR2_X1 U736 ( .A1(n667), .A2(n666), .ZN(n669) );
  XNOR2_X1 U737 ( .A(n669), .B(n668), .ZN(n680) );
  INV_X1 U738 ( .A(n680), .ZN(n670) );
  NAND2_X1 U739 ( .A1(n670), .A2(G286), .ZN(n676) );
  NOR2_X1 U740 ( .A1(G1971), .A2(n700), .ZN(n673) );
  NOR2_X1 U741 ( .A1(G2090), .A2(n671), .ZN(n672) );
  NOR2_X1 U742 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n674), .A2(G303), .ZN(n675) );
  NAND2_X1 U744 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U745 ( .A1(n677), .A2(G8), .ZN(n678) );
  XNOR2_X1 U746 ( .A(n678), .B(KEYINPUT32), .ZN(n685) );
  NAND2_X1 U747 ( .A1(G8), .A2(n679), .ZN(n683) );
  NOR2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U751 ( .A(KEYINPUT96), .B(n686), .ZN(n699) );
  NAND2_X1 U752 ( .A1(n687), .A2(n699), .ZN(n688) );
  NAND2_X1 U753 ( .A1(n688), .A2(n700), .ZN(n689) );
  XNOR2_X1 U754 ( .A(n689), .B(KEYINPUT98), .ZN(n693) );
  NOR2_X1 U755 ( .A1(G1981), .A2(G305), .ZN(n690) );
  XOR2_X1 U756 ( .A(n690), .B(KEYINPUT24), .Z(n691) );
  OR2_X1 U757 ( .A1(n700), .A2(n691), .ZN(n692) );
  AND2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n749) );
  NOR2_X1 U759 ( .A1(G1976), .A2(G288), .ZN(n696) );
  NAND2_X1 U760 ( .A1(n696), .A2(KEYINPUT33), .ZN(n694) );
  NOR2_X1 U761 ( .A1(n700), .A2(n694), .ZN(n705) );
  NOR2_X1 U762 ( .A1(G1971), .A2(G303), .ZN(n695) );
  NOR2_X1 U763 ( .A1(n696), .A2(n695), .ZN(n1020) );
  INV_X1 U764 ( .A(KEYINPUT33), .ZN(n697) );
  AND2_X1 U765 ( .A1(n1020), .A2(n697), .ZN(n698) );
  NAND2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U767 ( .A1(G1976), .A2(G288), .ZN(n1007) );
  INV_X1 U768 ( .A(n1007), .ZN(n701) );
  OR2_X1 U769 ( .A1(KEYINPUT33), .A2(n520), .ZN(n702) );
  NAND2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U771 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U772 ( .A(G1981), .B(G305), .Z(n1022) );
  NAND2_X1 U773 ( .A1(n706), .A2(n1022), .ZN(n747) );
  NAND2_X1 U774 ( .A1(G141), .A2(n877), .ZN(n708) );
  NAND2_X1 U775 ( .A1(G117), .A2(n874), .ZN(n707) );
  NAND2_X1 U776 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U777 ( .A1(n709), .A2(G105), .ZN(n710) );
  XOR2_X1 U778 ( .A(KEYINPUT38), .B(n710), .Z(n711) );
  NOR2_X1 U779 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U780 ( .A1(n521), .A2(G129), .ZN(n713) );
  NAND2_X1 U781 ( .A1(n714), .A2(n713), .ZN(n885) );
  NOR2_X1 U782 ( .A1(G1996), .A2(n885), .ZN(n954) );
  AND2_X1 U783 ( .A1(n885), .A2(G1996), .ZN(n724) );
  NAND2_X1 U784 ( .A1(G107), .A2(n874), .ZN(n716) );
  NAND2_X1 U785 ( .A1(G119), .A2(n521), .ZN(n715) );
  NAND2_X1 U786 ( .A1(n716), .A2(n715), .ZN(n721) );
  NAND2_X1 U787 ( .A1(G95), .A2(n709), .ZN(n718) );
  NAND2_X1 U788 ( .A1(G131), .A2(n877), .ZN(n717) );
  NAND2_X1 U789 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U790 ( .A(KEYINPUT86), .B(n719), .ZN(n720) );
  NOR2_X1 U791 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U792 ( .A(n722), .B(KEYINPUT87), .Z(n870) );
  INV_X1 U793 ( .A(G1991), .ZN(n925) );
  NOR2_X1 U794 ( .A1(n870), .A2(n925), .ZN(n723) );
  OR2_X1 U795 ( .A1(n724), .A2(n723), .ZN(n962) );
  NOR2_X1 U796 ( .A1(n726), .A2(n725), .ZN(n751) );
  NAND2_X1 U797 ( .A1(n962), .A2(n751), .ZN(n752) );
  INV_X1 U798 ( .A(n752), .ZN(n730) );
  NOR2_X1 U799 ( .A1(G1986), .A2(G290), .ZN(n728) );
  AND2_X1 U800 ( .A1(n925), .A2(n870), .ZN(n727) );
  XOR2_X1 U801 ( .A(KEYINPUT99), .B(n727), .Z(n961) );
  NOR2_X1 U802 ( .A1(n728), .A2(n961), .ZN(n729) );
  NOR2_X1 U803 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U804 ( .A1(n954), .A2(n731), .ZN(n732) );
  XNOR2_X1 U805 ( .A(n732), .B(KEYINPUT39), .ZN(n743) );
  NAND2_X1 U806 ( .A1(G104), .A2(n709), .ZN(n734) );
  NAND2_X1 U807 ( .A1(G140), .A2(n877), .ZN(n733) );
  NAND2_X1 U808 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U809 ( .A(KEYINPUT34), .B(n735), .ZN(n741) );
  NAND2_X1 U810 ( .A1(n521), .A2(G128), .ZN(n736) );
  XOR2_X1 U811 ( .A(KEYINPUT85), .B(n736), .Z(n738) );
  NAND2_X1 U812 ( .A1(n874), .A2(G116), .ZN(n737) );
  NAND2_X1 U813 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U814 ( .A(KEYINPUT35), .B(n739), .Z(n740) );
  NOR2_X1 U815 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U816 ( .A(KEYINPUT36), .B(n742), .ZN(n890) );
  XNOR2_X1 U817 ( .A(G2067), .B(KEYINPUT37), .ZN(n744) );
  NOR2_X1 U818 ( .A1(n890), .A2(n744), .ZN(n958) );
  NAND2_X1 U819 ( .A1(n751), .A2(n958), .ZN(n753) );
  NAND2_X1 U820 ( .A1(n743), .A2(n753), .ZN(n745) );
  NAND2_X1 U821 ( .A1(n890), .A2(n744), .ZN(n960) );
  NAND2_X1 U822 ( .A1(n745), .A2(n960), .ZN(n746) );
  NAND2_X1 U823 ( .A1(n746), .A2(n751), .ZN(n750) );
  AND2_X1 U824 ( .A1(n747), .A2(n750), .ZN(n748) );
  NAND2_X1 U825 ( .A1(n749), .A2(n748), .ZN(n759) );
  INV_X1 U826 ( .A(n750), .ZN(n757) );
  XNOR2_X1 U827 ( .A(G1986), .B(G290), .ZN(n1014) );
  AND2_X1 U828 ( .A1(n1014), .A2(n751), .ZN(n755) );
  NAND2_X1 U829 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U830 ( .A1(n755), .A2(n754), .ZN(n756) );
  OR2_X1 U831 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U832 ( .A(n761), .B(n760), .ZN(G329) );
  AND2_X1 U833 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U834 ( .A(G57), .ZN(G237) );
  INV_X1 U835 ( .A(G132), .ZN(G219) );
  INV_X1 U836 ( .A(G82), .ZN(G220) );
  NAND2_X1 U837 ( .A1(G7), .A2(G661), .ZN(n763) );
  XOR2_X1 U838 ( .A(n763), .B(KEYINPUT10), .Z(n921) );
  NAND2_X1 U839 ( .A1(n921), .A2(G567), .ZN(n764) );
  XOR2_X1 U840 ( .A(KEYINPUT11), .B(n764), .Z(G234) );
  INV_X1 U841 ( .A(G860), .ZN(n770) );
  OR2_X1 U842 ( .A1(n1027), .A2(n770), .ZN(G153) );
  NAND2_X1 U843 ( .A1(G868), .A2(G301), .ZN(n766) );
  OR2_X1 U844 ( .A1(n1008), .A2(G868), .ZN(n765) );
  NAND2_X1 U845 ( .A1(n766), .A2(n765), .ZN(G284) );
  INV_X1 U846 ( .A(G868), .ZN(n808) );
  NAND2_X1 U847 ( .A1(n1010), .A2(n808), .ZN(n767) );
  XNOR2_X1 U848 ( .A(n767), .B(KEYINPUT73), .ZN(n769) );
  NOR2_X1 U849 ( .A1(n808), .A2(G286), .ZN(n768) );
  NOR2_X1 U850 ( .A1(n769), .A2(n768), .ZN(G297) );
  NAND2_X1 U851 ( .A1(n770), .A2(G559), .ZN(n771) );
  NAND2_X1 U852 ( .A1(n771), .A2(n1008), .ZN(n772) );
  XNOR2_X1 U853 ( .A(n772), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U854 ( .A1(G868), .A2(n1027), .ZN(n773) );
  XNOR2_X1 U855 ( .A(KEYINPUT74), .B(n773), .ZN(n776) );
  NAND2_X1 U856 ( .A1(G868), .A2(n1008), .ZN(n774) );
  NOR2_X1 U857 ( .A1(G559), .A2(n774), .ZN(n775) );
  NOR2_X1 U858 ( .A1(n776), .A2(n775), .ZN(G282) );
  NAND2_X1 U859 ( .A1(G99), .A2(n709), .ZN(n778) );
  NAND2_X1 U860 ( .A1(G111), .A2(n874), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n778), .A2(n777), .ZN(n784) );
  NAND2_X1 U862 ( .A1(n521), .A2(G123), .ZN(n779) );
  XNOR2_X1 U863 ( .A(n779), .B(KEYINPUT18), .ZN(n781) );
  NAND2_X1 U864 ( .A1(G135), .A2(n877), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U866 ( .A(KEYINPUT75), .B(n782), .Z(n783) );
  NOR2_X1 U867 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U868 ( .A(KEYINPUT76), .B(n785), .Z(n945) );
  XNOR2_X1 U869 ( .A(n945), .B(G2096), .ZN(n786) );
  NOR2_X1 U870 ( .A1(G2100), .A2(n786), .ZN(n787) );
  XNOR2_X1 U871 ( .A(KEYINPUT77), .B(n787), .ZN(G156) );
  NAND2_X1 U872 ( .A1(G559), .A2(n1008), .ZN(n788) );
  XNOR2_X1 U873 ( .A(n788), .B(n1027), .ZN(n916) );
  NAND2_X1 U874 ( .A1(n789), .A2(G80), .ZN(n790) );
  XNOR2_X1 U875 ( .A(n790), .B(KEYINPUT80), .ZN(n800) );
  NAND2_X1 U876 ( .A1(G67), .A2(n791), .ZN(n794) );
  NAND2_X1 U877 ( .A1(G55), .A2(n792), .ZN(n793) );
  NAND2_X1 U878 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U879 ( .A1(G93), .A2(n795), .ZN(n796) );
  XNOR2_X1 U880 ( .A(KEYINPUT79), .B(n796), .ZN(n797) );
  NOR2_X1 U881 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U882 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U883 ( .A(KEYINPUT81), .B(n801), .Z(n919) );
  XOR2_X1 U884 ( .A(n919), .B(KEYINPUT19), .Z(n803) );
  XOR2_X1 U885 ( .A(G288), .B(G299), .Z(n802) );
  XNOR2_X1 U886 ( .A(n803), .B(n802), .ZN(n804) );
  XOR2_X1 U887 ( .A(G303), .B(n804), .Z(n806) );
  XNOR2_X1 U888 ( .A(G290), .B(G305), .ZN(n805) );
  XNOR2_X1 U889 ( .A(n806), .B(n805), .ZN(n893) );
  XNOR2_X1 U890 ( .A(n916), .B(n893), .ZN(n807) );
  NAND2_X1 U891 ( .A1(n807), .A2(G868), .ZN(n810) );
  NAND2_X1 U892 ( .A1(n808), .A2(n919), .ZN(n809) );
  NAND2_X1 U893 ( .A1(n810), .A2(n809), .ZN(G295) );
  XOR2_X1 U894 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n812) );
  NAND2_X1 U895 ( .A1(G2078), .A2(G2084), .ZN(n811) );
  XNOR2_X1 U896 ( .A(n812), .B(n811), .ZN(n813) );
  NAND2_X1 U897 ( .A1(G2090), .A2(n813), .ZN(n814) );
  XNOR2_X1 U898 ( .A(KEYINPUT21), .B(n814), .ZN(n815) );
  NAND2_X1 U899 ( .A1(n815), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U900 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U901 ( .A1(G220), .A2(G219), .ZN(n816) );
  XOR2_X1 U902 ( .A(KEYINPUT22), .B(n816), .Z(n817) );
  NOR2_X1 U903 ( .A1(G218), .A2(n817), .ZN(n818) );
  NAND2_X1 U904 ( .A1(G96), .A2(n818), .ZN(n914) );
  NAND2_X1 U905 ( .A1(n914), .A2(G2106), .ZN(n822) );
  NAND2_X1 U906 ( .A1(G69), .A2(G120), .ZN(n819) );
  NOR2_X1 U907 ( .A1(G237), .A2(n819), .ZN(n820) );
  NAND2_X1 U908 ( .A1(G108), .A2(n820), .ZN(n915) );
  NAND2_X1 U909 ( .A1(n915), .A2(G567), .ZN(n821) );
  NAND2_X1 U910 ( .A1(n822), .A2(n821), .ZN(n828) );
  NAND2_X1 U911 ( .A1(G661), .A2(G483), .ZN(n823) );
  NOR2_X1 U912 ( .A1(n828), .A2(n823), .ZN(n826) );
  NAND2_X1 U913 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n921), .ZN(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U916 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n825) );
  XNOR2_X1 U918 ( .A(KEYINPUT102), .B(n825), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(G188) );
  INV_X1 U920 ( .A(n828), .ZN(G319) );
  XOR2_X1 U921 ( .A(KEYINPUT104), .B(G1981), .Z(n831) );
  XOR2_X1 U922 ( .A(n829), .B(G1991), .Z(n830) );
  XNOR2_X1 U923 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U924 ( .A(n832), .B(KEYINPUT41), .Z(n834) );
  XNOR2_X1 U925 ( .A(G1986), .B(G1971), .ZN(n833) );
  XNOR2_X1 U926 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U927 ( .A(G1956), .B(G1961), .Z(n836) );
  XNOR2_X1 U928 ( .A(G1976), .B(G1966), .ZN(n835) );
  XNOR2_X1 U929 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U930 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U931 ( .A(KEYINPUT105), .B(G2474), .ZN(n839) );
  XNOR2_X1 U932 ( .A(n840), .B(n839), .ZN(G229) );
  XOR2_X1 U933 ( .A(KEYINPUT42), .B(G2072), .Z(n842) );
  XNOR2_X1 U934 ( .A(G2084), .B(G2078), .ZN(n841) );
  XNOR2_X1 U935 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U936 ( .A(n843), .B(G2100), .Z(n845) );
  XNOR2_X1 U937 ( .A(G2067), .B(G2090), .ZN(n844) );
  XNOR2_X1 U938 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U939 ( .A(G2096), .B(KEYINPUT43), .Z(n847) );
  XNOR2_X1 U940 ( .A(G2678), .B(KEYINPUT103), .ZN(n846) );
  XNOR2_X1 U941 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U942 ( .A(n849), .B(n848), .Z(G227) );
  NAND2_X1 U943 ( .A1(n874), .A2(G112), .ZN(n850) );
  XOR2_X1 U944 ( .A(KEYINPUT107), .B(n850), .Z(n852) );
  NAND2_X1 U945 ( .A1(n709), .A2(G100), .ZN(n851) );
  NAND2_X1 U946 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U947 ( .A(KEYINPUT108), .B(n853), .ZN(n859) );
  NAND2_X1 U948 ( .A1(G124), .A2(n521), .ZN(n854) );
  XNOR2_X1 U949 ( .A(n854), .B(KEYINPUT44), .ZN(n855) );
  XNOR2_X1 U950 ( .A(n855), .B(KEYINPUT106), .ZN(n857) );
  NAND2_X1 U951 ( .A1(G136), .A2(n877), .ZN(n856) );
  NAND2_X1 U952 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U953 ( .A1(n859), .A2(n858), .ZN(G162) );
  XOR2_X1 U954 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n861) );
  XNOR2_X1 U955 ( .A(KEYINPUT111), .B(KEYINPUT110), .ZN(n860) );
  XNOR2_X1 U956 ( .A(n861), .B(n860), .ZN(n869) );
  NAND2_X1 U957 ( .A1(G103), .A2(n709), .ZN(n863) );
  NAND2_X1 U958 ( .A1(G139), .A2(n877), .ZN(n862) );
  NAND2_X1 U959 ( .A1(n863), .A2(n862), .ZN(n868) );
  NAND2_X1 U960 ( .A1(G115), .A2(n874), .ZN(n865) );
  NAND2_X1 U961 ( .A1(G127), .A2(n521), .ZN(n864) );
  NAND2_X1 U962 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U963 ( .A(KEYINPUT47), .B(n866), .Z(n867) );
  NOR2_X1 U964 ( .A1(n868), .A2(n867), .ZN(n947) );
  XOR2_X1 U965 ( .A(n869), .B(n947), .Z(n872) );
  XNOR2_X1 U966 ( .A(G164), .B(n870), .ZN(n871) );
  XNOR2_X1 U967 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U968 ( .A(n945), .B(n873), .ZN(n889) );
  NAND2_X1 U969 ( .A1(G118), .A2(n874), .ZN(n876) );
  NAND2_X1 U970 ( .A1(G130), .A2(n521), .ZN(n875) );
  NAND2_X1 U971 ( .A1(n876), .A2(n875), .ZN(n883) );
  NAND2_X1 U972 ( .A1(G106), .A2(n709), .ZN(n879) );
  NAND2_X1 U973 ( .A1(G142), .A2(n877), .ZN(n878) );
  NAND2_X1 U974 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U975 ( .A(KEYINPUT45), .B(n880), .ZN(n881) );
  XNOR2_X1 U976 ( .A(KEYINPUT109), .B(n881), .ZN(n882) );
  NOR2_X1 U977 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U978 ( .A(n884), .B(G162), .Z(n887) );
  XOR2_X1 U979 ( .A(G160), .B(n885), .Z(n886) );
  XNOR2_X1 U980 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U981 ( .A(n889), .B(n888), .ZN(n891) );
  XOR2_X1 U982 ( .A(n891), .B(n890), .Z(n892) );
  NOR2_X1 U983 ( .A1(G37), .A2(n892), .ZN(G395) );
  XOR2_X1 U984 ( .A(n893), .B(G286), .Z(n895) );
  XOR2_X1 U985 ( .A(G301), .B(n1008), .Z(n894) );
  XNOR2_X1 U986 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U987 ( .A(n896), .B(n1027), .ZN(n897) );
  NOR2_X1 U988 ( .A1(G37), .A2(n897), .ZN(G397) );
  XNOR2_X1 U989 ( .A(G2454), .B(G2443), .ZN(n907) );
  XOR2_X1 U990 ( .A(G2430), .B(KEYINPUT100), .Z(n899) );
  XNOR2_X1 U991 ( .A(G2446), .B(KEYINPUT101), .ZN(n898) );
  XNOR2_X1 U992 ( .A(n899), .B(n898), .ZN(n903) );
  XOR2_X1 U993 ( .A(G2451), .B(G2427), .Z(n901) );
  XOR2_X1 U994 ( .A(n977), .B(G1341), .Z(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U996 ( .A(n903), .B(n902), .Z(n905) );
  XNOR2_X1 U997 ( .A(G2435), .B(G2438), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U999 ( .A(n907), .B(n906), .ZN(n908) );
  NAND2_X1 U1000 ( .A1(n908), .A2(G14), .ZN(n920) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n920), .ZN(n911) );
  NOR2_X1 U1002 ( .A1(G229), .A2(G227), .ZN(n909) );
  XNOR2_X1 U1003 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1004 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1006 ( .A1(n913), .A2(n912), .ZN(G225) );
  XOR2_X1 U1007 ( .A(KEYINPUT112), .B(G225), .Z(G308) );
  INV_X1 U1009 ( .A(G120), .ZN(G236) );
  INV_X1 U1010 ( .A(G96), .ZN(G221) );
  INV_X1 U1011 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(G325) );
  INV_X1 U1013 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1014 ( .A(KEYINPUT78), .B(n916), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(G860), .A2(n917), .ZN(n918) );
  XOR2_X1 U1016 ( .A(n919), .B(n918), .Z(G145) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  INV_X1 U1018 ( .A(n920), .ZN(G401) );
  INV_X1 U1019 ( .A(n921), .ZN(G223) );
  INV_X1 U1020 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U1021 ( .A(KEYINPUT115), .B(G2090), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(n922), .B(G35), .ZN(n941) );
  XOR2_X1 U1023 ( .A(KEYINPUT117), .B(G34), .Z(n924) );
  XNOR2_X1 U1024 ( .A(G2084), .B(KEYINPUT54), .ZN(n923) );
  XNOR2_X1 U1025 ( .A(n924), .B(n923), .ZN(n939) );
  XOR2_X1 U1026 ( .A(n925), .B(G25), .Z(n927) );
  XNOR2_X1 U1027 ( .A(G33), .B(G2072), .ZN(n926) );
  NOR2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n933) );
  XOR2_X1 U1029 ( .A(G32), .B(G1996), .Z(n928) );
  NAND2_X1 U1030 ( .A1(n928), .A2(G28), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(KEYINPUT116), .B(G2067), .ZN(n929) );
  XNOR2_X1 U1032 ( .A(G26), .B(n929), .ZN(n930) );
  NOR2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(G27), .B(n934), .ZN(n935) );
  NOR2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(n937), .B(KEYINPUT53), .ZN(n938) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n944) );
  NOR2_X1 U1040 ( .A1(G29), .A2(KEYINPUT55), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n942), .ZN(n943) );
  NAND2_X1 U1042 ( .A1(G11), .A2(n943), .ZN(n976) );
  INV_X1 U1043 ( .A(KEYINPUT55), .ZN(n970) );
  OR2_X1 U1044 ( .A1(n970), .A2(n944), .ZN(n974) );
  XNOR2_X1 U1045 ( .A(G160), .B(G2084), .ZN(n946) );
  NAND2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n968) );
  XNOR2_X1 U1047 ( .A(G2072), .B(n947), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(G164), .B(G2078), .ZN(n948) );
  XNOR2_X1 U1049 ( .A(n948), .B(KEYINPUT114), .ZN(n949) );
  NAND2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1051 ( .A(n951), .B(KEYINPUT50), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(G2090), .B(G162), .ZN(n952) );
  XNOR2_X1 U1053 ( .A(n952), .B(KEYINPUT113), .ZN(n953) );
  NOR2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1055 ( .A(KEYINPUT51), .B(n955), .ZN(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n966) );
  INV_X1 U1057 ( .A(n958), .ZN(n959) );
  NAND2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n964) );
  OR2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n969), .B(KEYINPUT52), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(G29), .A2(n972), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n1036) );
  XOR2_X1 U1068 ( .A(KEYINPUT59), .B(n977), .Z(n978) );
  XNOR2_X1 U1069 ( .A(n978), .B(G4), .ZN(n986) );
  XNOR2_X1 U1070 ( .A(G1956), .B(G20), .ZN(n984) );
  XNOR2_X1 U1071 ( .A(G1341), .B(G19), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(n979), .B(KEYINPUT120), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(G6), .B(G1981), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(KEYINPUT121), .B(n982), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(KEYINPUT60), .B(n987), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(G21), .B(G1966), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(KEYINPUT122), .B(n988), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1082 ( .A(KEYINPUT123), .B(n991), .Z(n1000) );
  XOR2_X1 U1083 ( .A(G1986), .B(KEYINPUT125), .Z(n992) );
  XNOR2_X1 U1084 ( .A(G24), .B(n992), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(G1976), .B(G23), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(G22), .B(G1971), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1088 ( .A(KEYINPUT124), .B(n995), .Z(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1090 ( .A(KEYINPUT58), .B(n998), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(G5), .B(G1961), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1094 ( .A(KEYINPUT61), .B(n1003), .Z(n1004) );
  NOR2_X1 U1095 ( .A1(G16), .A2(n1004), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(KEYINPUT126), .B(n1005), .ZN(n1033) );
  NAND2_X1 U1097 ( .A1(G1971), .A2(G303), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1018) );
  XNOR2_X1 U1099 ( .A(n1008), .B(KEYINPUT118), .ZN(n1009) );
  XOR2_X1 U1100 ( .A(n1009), .B(G1348), .Z(n1012) );
  XOR2_X1 U1101 ( .A(G1956), .B(n1010), .Z(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(G1961), .B(G171), .Z(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(KEYINPUT119), .B(n1021), .ZN(n1026) );
  XNOR2_X1 U1109 ( .A(G1966), .B(G168), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1111 ( .A(n1024), .B(KEYINPUT57), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(G1341), .B(n1027), .ZN(n1028) );
  NOR2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(KEYINPUT56), .B(G16), .Z(n1030) );
  NOR2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1117 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1118 ( .A(KEYINPUT127), .B(n1034), .Z(n1035) );
  NAND2_X1 U1119 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1120 ( .A(KEYINPUT62), .B(n1037), .ZN(G150) );
  INV_X1 U1121 ( .A(G150), .ZN(G311) );
endmodule

