

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757;

  NAND2_X1 U368 ( .A1(n700), .A2(n701), .ZN(n599) );
  XOR2_X1 U369 ( .A(G131), .B(KEYINPUT69), .Z(n347) );
  NOR2_X2 U370 ( .A1(n594), .A2(n595), .ZN(n596) );
  NOR2_X2 U371 ( .A1(n594), .A2(n581), .ZN(n366) );
  NAND2_X2 U372 ( .A1(n614), .A2(n615), .ZN(n420) );
  XNOR2_X2 U373 ( .A(n400), .B(n355), .ZN(n531) );
  OR2_X2 U374 ( .A1(n729), .A2(G902), .ZN(n400) );
  XNOR2_X2 U375 ( .A(n492), .B(n491), .ZN(n584) );
  AND2_X1 U376 ( .A1(n425), .A2(n693), .ZN(n740) );
  INV_X1 U377 ( .A(n562), .ZN(n700) );
  AND2_X1 U378 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U379 ( .A1(n417), .A2(n416), .ZN(n602) );
  XNOR2_X1 U380 ( .A(n347), .B(n434), .ZN(n459) );
  XNOR2_X1 U381 ( .A(G146), .B(KEYINPUT68), .ZN(n434) );
  XNOR2_X1 U382 ( .A(G146), .B(G125), .ZN(n510) );
  NOR2_X1 U383 ( .A1(n599), .A2(n699), .ZN(n706) );
  XNOR2_X1 U384 ( .A(n366), .B(n360), .ZN(n607) );
  XNOR2_X1 U385 ( .A(n543), .B(n542), .ZN(n568) );
  NAND2_X1 U386 ( .A1(n541), .A2(n540), .ZN(n543) );
  NOR2_X1 U387 ( .A1(n667), .A2(n739), .ZN(n669) );
  NOR2_X1 U388 ( .A1(n650), .A2(n739), .ZN(n652) );
  AND2_X1 U389 ( .A1(n635), .A2(G475), .ZN(n421) );
  NOR2_X1 U390 ( .A1(n544), .A2(n568), .ZN(n683) );
  XNOR2_X2 U391 ( .A(n569), .B(n429), .ZN(n600) );
  NOR2_X1 U392 ( .A1(n695), .A2(n523), .ZN(n536) );
  XNOR2_X1 U393 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n443) );
  XNOR2_X1 U394 ( .A(n472), .B(n473), .ZN(n742) );
  NAND2_X1 U395 ( .A1(n368), .A2(n367), .ZN(n625) );
  AND2_X1 U396 ( .A1(n683), .A2(n359), .ZN(n547) );
  NOR2_X1 U397 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U398 ( .A(n379), .B(n556), .ZN(n378) );
  XOR2_X1 U399 ( .A(KEYINPUT100), .B(KEYINPUT11), .Z(n436) );
  XOR2_X1 U400 ( .A(G140), .B(G104), .Z(n475) );
  AND2_X1 U401 ( .A1(n740), .A2(n620), .ZN(n361) );
  INV_X1 U402 ( .A(KEYINPUT116), .ZN(n365) );
  NOR2_X1 U403 ( .A1(n710), .A2(n709), .ZN(n431) );
  XNOR2_X1 U404 ( .A(n541), .B(KEYINPUT38), .ZN(n710) );
  INV_X1 U405 ( .A(n532), .ZN(n522) );
  NOR2_X1 U406 ( .A1(n584), .A2(n695), .ZN(n701) );
  XNOR2_X1 U407 ( .A(n461), .B(n460), .ZN(n472) );
  XNOR2_X1 U408 ( .A(n459), .B(n432), .ZN(n461) );
  XOR2_X1 U409 ( .A(G137), .B(KEYINPUT4), .Z(n432) );
  XNOR2_X1 U410 ( .A(n408), .B(n407), .ZN(n504) );
  XNOR2_X1 U411 ( .A(G119), .B(G116), .ZN(n407) );
  XNOR2_X1 U412 ( .A(n462), .B(G113), .ZN(n408) );
  INV_X1 U413 ( .A(KEYINPUT3), .ZN(n462) );
  XNOR2_X1 U414 ( .A(n427), .B(n426), .ZN(n627) );
  XNOR2_X1 U415 ( .A(n485), .B(n487), .ZN(n426) );
  XNOR2_X1 U416 ( .A(n483), .B(n486), .ZN(n427) );
  XNOR2_X1 U417 ( .A(n381), .B(n440), .ZN(n664) );
  XNOR2_X1 U418 ( .A(n382), .B(n384), .ZN(n381) );
  XNOR2_X1 U419 ( .A(n380), .B(n456), .ZN(n546) );
  INV_X1 U420 ( .A(KEYINPUT101), .ZN(n456) );
  NAND2_X1 U421 ( .A1(n531), .A2(n701), .ZN(n595) );
  BUF_X1 U422 ( .A(n562), .Z(n606) );
  NAND2_X1 U423 ( .A1(n636), .A2(n348), .ZN(n403) );
  AND2_X1 U424 ( .A1(n399), .A2(n353), .ZN(n398) );
  NAND2_X1 U425 ( .A1(G237), .A2(G234), .ZN(n496) );
  INV_X1 U426 ( .A(n706), .ZN(n362) );
  XNOR2_X1 U427 ( .A(n705), .B(KEYINPUT115), .ZN(n363) );
  XNOR2_X1 U428 ( .A(n376), .B(n375), .ZN(n425) );
  INV_X1 U429 ( .A(KEYINPUT84), .ZN(n375) );
  NAND2_X1 U430 ( .A1(n378), .A2(n377), .ZN(n376) );
  XNOR2_X1 U431 ( .A(n383), .B(n437), .ZN(n382) );
  XNOR2_X1 U432 ( .A(n436), .B(n435), .ZN(n383) );
  XNOR2_X1 U433 ( .A(G143), .B(G113), .ZN(n435) );
  INV_X1 U434 ( .A(n459), .ZN(n384) );
  XNOR2_X1 U435 ( .A(G140), .B(G125), .ZN(n438) );
  XNOR2_X1 U436 ( .A(n452), .B(n451), .ZN(n514) );
  INV_X1 U437 ( .A(G128), .ZN(n451) );
  XNOR2_X1 U438 ( .A(G143), .B(KEYINPUT64), .ZN(n452) );
  XNOR2_X1 U439 ( .A(KEYINPUT88), .B(KEYINPUT4), .ZN(n507) );
  XNOR2_X1 U440 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n508) );
  INV_X1 U441 ( .A(KEYINPUT104), .ZN(n374) );
  OR2_X1 U442 ( .A1(n538), .A2(n548), .ZN(n393) );
  INV_X1 U443 ( .A(KEYINPUT36), .ZN(n395) );
  XNOR2_X1 U444 ( .A(n531), .B(n530), .ZN(n562) );
  XNOR2_X1 U445 ( .A(G107), .B(G116), .ZN(n448) );
  XOR2_X1 U446 ( .A(G122), .B(KEYINPUT9), .Z(n446) );
  XNOR2_X1 U447 ( .A(n514), .B(G134), .ZN(n460) );
  XNOR2_X1 U448 ( .A(n742), .B(n477), .ZN(n729) );
  XOR2_X1 U449 ( .A(KEYINPUT41), .B(n528), .Z(n722) );
  AND2_X1 U450 ( .A1(n501), .A2(n404), .ZN(n519) );
  AND2_X1 U451 ( .A1(n502), .A2(n405), .ZN(n404) );
  INV_X1 U452 ( .A(n606), .ZN(n394) );
  NOR2_X1 U453 ( .A1(n393), .A2(n395), .ZN(n392) );
  NOR2_X1 U454 ( .A1(n595), .A2(n532), .ZN(n501) );
  XNOR2_X1 U455 ( .A(n527), .B(KEYINPUT108), .ZN(n544) );
  NOR2_X1 U456 ( .A1(n627), .A2(G902), .ZN(n492) );
  XNOR2_X1 U457 ( .A(n455), .B(G478), .ZN(n545) );
  XNOR2_X1 U458 ( .A(n442), .B(n441), .ZN(n551) );
  INV_X2 U459 ( .A(G953), .ZN(n750) );
  XNOR2_X1 U460 ( .A(n506), .B(n503), .ZN(n409) );
  NAND2_X1 U461 ( .A1(n387), .A2(n385), .ZN(n691) );
  NAND2_X1 U462 ( .A1(n386), .A2(n392), .ZN(n385) );
  NAND2_X1 U463 ( .A1(n388), .A2(n394), .ZN(n387) );
  AND2_X1 U464 ( .A1(n391), .A2(n394), .ZN(n386) );
  XNOR2_X1 U465 ( .A(n583), .B(KEYINPUT32), .ZN(n643) );
  XNOR2_X1 U466 ( .A(n546), .B(KEYINPUT105), .ZN(n682) );
  NAND2_X1 U467 ( .A1(n402), .A2(n401), .ZN(n369) );
  XNOR2_X1 U468 ( .A(n403), .B(n640), .ZN(n402) );
  INV_X1 U469 ( .A(KEYINPUT118), .ZN(n371) );
  AND2_X1 U470 ( .A1(n635), .A2(G472), .ZN(n348) );
  AND2_X1 U471 ( .A1(n425), .A2(n357), .ZN(n349) );
  AND2_X1 U472 ( .A1(n363), .A2(n362), .ZN(n350) );
  XOR2_X1 U473 ( .A(G137), .B(G146), .Z(n351) );
  XOR2_X1 U474 ( .A(KEYINPUT94), .B(KEYINPUT80), .Z(n352) );
  AND2_X1 U475 ( .A1(n555), .A2(n554), .ZN(n353) );
  AND2_X1 U476 ( .A1(n688), .A2(n418), .ZN(n354) );
  XOR2_X1 U477 ( .A(n478), .B(KEYINPUT70), .Z(n355) );
  AND2_X1 U478 ( .A1(n635), .A2(G217), .ZN(n356) );
  AND2_X1 U479 ( .A1(n693), .A2(n619), .ZN(n357) );
  AND2_X1 U480 ( .A1(n724), .A2(n723), .ZN(n358) );
  AND2_X1 U481 ( .A1(n714), .A2(n423), .ZN(n359) );
  XOR2_X1 U482 ( .A(KEYINPUT73), .B(KEYINPUT22), .Z(n360) );
  XNOR2_X1 U483 ( .A(n409), .B(n504), .ZN(n659) );
  INV_X1 U484 ( .A(KEYINPUT99), .ZN(n418) );
  XNOR2_X1 U485 ( .A(n631), .B(KEYINPUT87), .ZN(n739) );
  INV_X1 U486 ( .A(n739), .ZN(n401) );
  NAND2_X1 U487 ( .A1(n361), .A2(n653), .ZN(n368) );
  NAND2_X1 U488 ( .A1(n364), .A2(n718), .ZN(n719) );
  XNOR2_X1 U489 ( .A(n708), .B(n365), .ZN(n364) );
  NOR2_X2 U490 ( .A1(G953), .A2(n727), .ZN(n728) );
  NOR2_X1 U491 ( .A1(n726), .A2(n358), .ZN(n370) );
  INV_X1 U492 ( .A(KEYINPUT82), .ZN(n367) );
  AND2_X1 U493 ( .A1(n414), .A2(n714), .ZN(n413) );
  NAND2_X2 U494 ( .A1(n626), .A2(KEYINPUT2), .ZN(n635) );
  XNOR2_X1 U495 ( .A(n369), .B(KEYINPUT63), .ZN(G57) );
  AND2_X2 U496 ( .A1(n643), .A2(n642), .ZN(n611) );
  AND2_X2 U497 ( .A1(n370), .A2(n725), .ZN(n372) );
  XNOR2_X2 U498 ( .A(n372), .B(n371), .ZN(n727) );
  NAND2_X1 U499 ( .A1(n373), .A2(n537), .ZN(n563) );
  XNOR2_X1 U500 ( .A(n599), .B(n374), .ZN(n373) );
  INV_X1 U501 ( .A(n645), .ZN(n377) );
  NAND2_X1 U502 ( .A1(n398), .A2(n396), .ZN(n379) );
  NAND2_X1 U503 ( .A1(n545), .A2(n551), .ZN(n380) );
  NAND2_X1 U504 ( .A1(n389), .A2(n390), .ZN(n388) );
  NAND2_X1 U505 ( .A1(n393), .A2(n395), .ZN(n389) );
  NAND2_X1 U506 ( .A1(n539), .A2(n395), .ZN(n390) );
  INV_X1 U507 ( .A(n539), .ZN(n391) );
  NOR2_X1 U508 ( .A1(n538), .A2(n539), .ZN(n557) );
  XNOR2_X1 U509 ( .A(n397), .B(KEYINPUT46), .ZN(n396) );
  NOR2_X1 U510 ( .A1(n756), .A2(n755), .ZN(n397) );
  XNOR2_X1 U511 ( .A(n691), .B(KEYINPUT85), .ZN(n399) );
  NAND2_X1 U512 ( .A1(n501), .A2(n502), .ZN(n406) );
  INV_X1 U513 ( .A(n710), .ZN(n405) );
  NOR2_X1 U514 ( .A1(n406), .A2(n548), .ZN(n549) );
  XNOR2_X2 U515 ( .A(n576), .B(n575), .ZN(n757) );
  XNOR2_X2 U516 ( .A(n411), .B(n410), .ZN(n503) );
  XNOR2_X2 U517 ( .A(KEYINPUT76), .B(G110), .ZN(n410) );
  XNOR2_X2 U518 ( .A(G107), .B(G101), .ZN(n411) );
  NAND2_X1 U519 ( .A1(n672), .A2(n354), .ZN(n412) );
  XNOR2_X2 U520 ( .A(n598), .B(KEYINPUT98), .ZN(n672) );
  NAND2_X1 U521 ( .A1(n413), .A2(n412), .ZN(n416) );
  NAND2_X1 U522 ( .A1(n415), .A2(KEYINPUT99), .ZN(n414) );
  INV_X1 U523 ( .A(n688), .ZN(n415) );
  NOR2_X1 U524 ( .A1(n672), .A2(n418), .ZN(n417) );
  XNOR2_X2 U525 ( .A(n601), .B(n419), .ZN(n688) );
  INV_X1 U526 ( .A(KEYINPUT31), .ZN(n419) );
  AND2_X2 U527 ( .A1(n740), .A2(n653), .ZN(n626) );
  XNOR2_X2 U528 ( .A(n420), .B(n617), .ZN(n653) );
  AND2_X1 U529 ( .A1(n636), .A2(n635), .ZN(n735) );
  NAND2_X1 U530 ( .A1(n636), .A2(n356), .ZN(n629) );
  NAND2_X1 U531 ( .A1(n636), .A2(n421), .ZN(n666) );
  NAND2_X1 U532 ( .A1(n636), .A2(n422), .ZN(n649) );
  AND2_X1 U533 ( .A1(n635), .A2(G210), .ZN(n422) );
  NAND2_X1 U534 ( .A1(n683), .A2(n714), .ZN(n424) );
  INV_X1 U535 ( .A(KEYINPUT47), .ZN(n423) );
  NAND2_X1 U536 ( .A1(n424), .A2(KEYINPUT47), .ZN(n553) );
  NAND2_X1 U537 ( .A1(n653), .A2(n349), .ZN(n623) );
  NAND2_X2 U538 ( .A1(n625), .A2(n624), .ZN(n636) );
  XNOR2_X2 U539 ( .A(n518), .B(n517), .ZN(n541) );
  OR2_X2 U540 ( .A1(n647), .A2(n620), .ZN(n518) );
  NAND2_X1 U541 ( .A1(n428), .A2(n536), .ZN(n525) );
  AND2_X1 U542 ( .A1(n534), .A2(n522), .ZN(n428) );
  XOR2_X1 U543 ( .A(KEYINPUT67), .B(KEYINPUT0), .Z(n429) );
  XOR2_X1 U544 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n430) );
  XOR2_X1 U545 ( .A(n466), .B(n465), .Z(n433) );
  INV_X1 U546 ( .A(KEYINPUT48), .ZN(n556) );
  INV_X1 U547 ( .A(n741), .ZN(n486) );
  INV_X1 U548 ( .A(KEYINPUT28), .ZN(n524) );
  XNOR2_X1 U549 ( .A(n467), .B(n433), .ZN(n468) );
  INV_X1 U550 ( .A(KEYINPUT7), .ZN(n447) );
  XNOR2_X1 U551 ( .A(n472), .B(n468), .ZN(n639) );
  XNOR2_X1 U552 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U553 ( .A(n450), .B(n449), .ZN(n454) );
  INV_X1 U554 ( .A(KEYINPUT122), .ZN(n633) );
  NOR2_X1 U555 ( .A1(G953), .A2(G237), .ZN(n463) );
  NAND2_X1 U556 ( .A1(G214), .A2(n463), .ZN(n437) );
  XNOR2_X2 U557 ( .A(G122), .B(G104), .ZN(n505) );
  XNOR2_X1 U558 ( .A(n505), .B(KEYINPUT12), .ZN(n439) );
  XNOR2_X1 U559 ( .A(KEYINPUT10), .B(n438), .ZN(n741) );
  XNOR2_X1 U560 ( .A(n439), .B(n741), .ZN(n440) );
  INV_X1 U561 ( .A(G902), .ZN(n469) );
  NAND2_X1 U562 ( .A1(n664), .A2(n469), .ZN(n442) );
  XOR2_X1 U563 ( .A(KEYINPUT13), .B(G475), .Z(n441) );
  NAND2_X1 U564 ( .A1(n750), .A2(G234), .ZN(n444) );
  XNOR2_X1 U565 ( .A(n444), .B(n443), .ZN(n484) );
  NAND2_X1 U566 ( .A1(G217), .A2(n484), .ZN(n445) );
  XNOR2_X1 U567 ( .A(n446), .B(n445), .ZN(n450) );
  INV_X1 U568 ( .A(n460), .ZN(n453) );
  XNOR2_X1 U569 ( .A(n454), .B(n453), .ZN(n736) );
  NOR2_X1 U570 ( .A1(n736), .A2(G902), .ZN(n455) );
  INV_X1 U571 ( .A(G237), .ZN(n457) );
  NAND2_X1 U572 ( .A1(n469), .A2(n457), .ZN(n516) );
  NAND2_X1 U573 ( .A1(n516), .A2(G214), .ZN(n458) );
  XNOR2_X1 U574 ( .A(n458), .B(KEYINPUT89), .ZN(n709) );
  NAND2_X1 U575 ( .A1(n463), .A2(G210), .ZN(n464) );
  XNOR2_X1 U576 ( .A(n504), .B(n464), .ZN(n467) );
  XOR2_X1 U577 ( .A(KEYINPUT97), .B(KEYINPUT75), .Z(n466) );
  XNOR2_X1 U578 ( .A(G101), .B(KEYINPUT5), .ZN(n465) );
  NAND2_X1 U579 ( .A1(n639), .A2(n469), .ZN(n470) );
  INV_X1 U580 ( .A(G472), .ZN(n637) );
  XNOR2_X1 U581 ( .A(n470), .B(n637), .ZN(n521) );
  NOR2_X1 U582 ( .A1(n709), .A2(n521), .ZN(n471) );
  XNOR2_X1 U583 ( .A(KEYINPUT30), .B(n471), .ZN(n502) );
  INV_X1 U584 ( .A(KEYINPUT92), .ZN(n473) );
  NAND2_X1 U585 ( .A1(G227), .A2(n750), .ZN(n474) );
  XNOR2_X1 U586 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U587 ( .A(n503), .B(n476), .Z(n477) );
  INV_X1 U588 ( .A(G469), .ZN(n478) );
  XNOR2_X1 U589 ( .A(G119), .B(G128), .ZN(n479) );
  XNOR2_X1 U590 ( .A(n351), .B(n479), .ZN(n482) );
  XNOR2_X1 U591 ( .A(G110), .B(KEYINPUT93), .ZN(n480) );
  XNOR2_X1 U592 ( .A(n352), .B(n480), .ZN(n481) );
  XNOR2_X1 U593 ( .A(n482), .B(n481), .ZN(n483) );
  NAND2_X1 U594 ( .A1(G221), .A2(n484), .ZN(n485) );
  XNOR2_X1 U595 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n487) );
  XOR2_X1 U596 ( .A(KEYINPUT77), .B(KEYINPUT25), .Z(n490) );
  XNOR2_X1 U597 ( .A(G902), .B(KEYINPUT15), .ZN(n618) );
  NAND2_X1 U598 ( .A1(n618), .A2(G234), .ZN(n488) );
  XNOR2_X1 U599 ( .A(n488), .B(KEYINPUT20), .ZN(n493) );
  AND2_X1 U600 ( .A1(n493), .A2(G217), .ZN(n489) );
  XNOR2_X1 U601 ( .A(n490), .B(n489), .ZN(n491) );
  AND2_X1 U602 ( .A1(n493), .A2(G221), .ZN(n495) );
  XNOR2_X1 U603 ( .A(KEYINPUT95), .B(KEYINPUT21), .ZN(n494) );
  XNOR2_X1 U604 ( .A(n495), .B(n494), .ZN(n695) );
  XNOR2_X1 U605 ( .A(n496), .B(KEYINPUT14), .ZN(n497) );
  NAND2_X1 U606 ( .A1(G952), .A2(n497), .ZN(n721) );
  NOR2_X1 U607 ( .A1(n721), .A2(G953), .ZN(n565) );
  NAND2_X1 U608 ( .A1(n497), .A2(G902), .ZN(n498) );
  XOR2_X1 U609 ( .A(n498), .B(KEYINPUT91), .Z(n564) );
  OR2_X1 U610 ( .A1(n750), .A2(n564), .ZN(n499) );
  NOR2_X1 U611 ( .A1(G900), .A2(n499), .ZN(n500) );
  NOR2_X1 U612 ( .A1(n565), .A2(n500), .ZN(n532) );
  XNOR2_X1 U613 ( .A(n505), .B(KEYINPUT16), .ZN(n506) );
  XNOR2_X1 U614 ( .A(n508), .B(n507), .ZN(n512) );
  NAND2_X1 U615 ( .A1(n750), .A2(G224), .ZN(n509) );
  XNOR2_X1 U616 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U617 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U618 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U619 ( .A(n659), .B(n515), .ZN(n647) );
  INV_X1 U620 ( .A(n618), .ZN(n620) );
  AND2_X1 U621 ( .A1(n516), .A2(G210), .ZN(n517) );
  INV_X1 U622 ( .A(n541), .ZN(n548) );
  XNOR2_X1 U623 ( .A(n519), .B(KEYINPUT39), .ZN(n561) );
  NOR2_X1 U624 ( .A1(n546), .A2(n561), .ZN(n520) );
  XNOR2_X1 U625 ( .A(n520), .B(KEYINPUT40), .ZN(n756) );
  INV_X1 U626 ( .A(n521), .ZN(n534) );
  INV_X1 U627 ( .A(n584), .ZN(n523) );
  XNOR2_X1 U628 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U629 ( .A1(n526), .A2(n531), .ZN(n527) );
  INV_X1 U630 ( .A(n545), .ZN(n550) );
  NOR2_X1 U631 ( .A1(n551), .A2(n550), .ZN(n712) );
  NAND2_X1 U632 ( .A1(n431), .A2(n712), .ZN(n528) );
  NOR2_X1 U633 ( .A1(n544), .A2(n722), .ZN(n529) );
  XNOR2_X1 U634 ( .A(n529), .B(KEYINPUT42), .ZN(n755) );
  INV_X1 U635 ( .A(KEYINPUT1), .ZN(n530) );
  NOR2_X1 U636 ( .A1(n532), .A2(n709), .ZN(n533) );
  NAND2_X1 U637 ( .A1(n682), .A2(n533), .ZN(n539) );
  INV_X1 U638 ( .A(n534), .ZN(n699) );
  INV_X1 U639 ( .A(KEYINPUT6), .ZN(n535) );
  XNOR2_X1 U640 ( .A(n699), .B(n535), .ZN(n604) );
  INV_X1 U641 ( .A(n604), .ZN(n537) );
  NAND2_X1 U642 ( .A1(n537), .A2(n536), .ZN(n538) );
  INV_X1 U643 ( .A(n709), .ZN(n540) );
  INV_X1 U644 ( .A(KEYINPUT19), .ZN(n542) );
  OR2_X1 U645 ( .A1(n551), .A2(n545), .ZN(n689) );
  NAND2_X1 U646 ( .A1(n689), .A2(n546), .ZN(n714) );
  XOR2_X1 U647 ( .A(n547), .B(KEYINPUT74), .Z(n555) );
  XOR2_X1 U648 ( .A(KEYINPUT107), .B(n549), .Z(n552) );
  AND2_X1 U649 ( .A1(n551), .A2(n550), .ZN(n572) );
  NAND2_X1 U650 ( .A1(n552), .A2(n572), .ZN(n681) );
  AND2_X1 U651 ( .A1(n553), .A2(n681), .ZN(n554) );
  XOR2_X1 U652 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n559) );
  NAND2_X1 U653 ( .A1(n557), .A2(n606), .ZN(n558) );
  XNOR2_X1 U654 ( .A(n559), .B(n558), .ZN(n560) );
  NOR2_X1 U655 ( .A1(n560), .A2(n541), .ZN(n645) );
  OR2_X1 U656 ( .A1(n561), .A2(n689), .ZN(n693) );
  XNOR2_X2 U657 ( .A(n563), .B(n430), .ZN(n723) );
  XOR2_X1 U658 ( .A(G898), .B(KEYINPUT90), .Z(n656) );
  NAND2_X1 U659 ( .A1(G953), .A2(n656), .ZN(n660) );
  NOR2_X1 U660 ( .A1(n564), .A2(n660), .ZN(n566) );
  NOR2_X1 U661 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X2 U662 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U663 ( .A1(n723), .A2(n600), .ZN(n571) );
  XOR2_X1 U664 ( .A(KEYINPUT72), .B(KEYINPUT34), .Z(n570) );
  XNOR2_X1 U665 ( .A(n571), .B(n570), .ZN(n573) );
  NAND2_X1 U666 ( .A1(n573), .A2(n572), .ZN(n576) );
  INV_X1 U667 ( .A(KEYINPUT78), .ZN(n574) );
  XNOR2_X1 U668 ( .A(n574), .B(KEYINPUT35), .ZN(n575) );
  INV_X1 U669 ( .A(KEYINPUT103), .ZN(n577) );
  XNOR2_X1 U670 ( .A(n584), .B(n577), .ZN(n696) );
  INV_X1 U671 ( .A(n696), .ZN(n603) );
  OR2_X1 U672 ( .A1(n606), .A2(n603), .ZN(n579) );
  XNOR2_X1 U673 ( .A(n604), .B(KEYINPUT79), .ZN(n578) );
  NOR2_X1 U674 ( .A1(n579), .A2(n578), .ZN(n582) );
  INV_X1 U675 ( .A(n600), .ZN(n594) );
  INV_X1 U676 ( .A(n695), .ZN(n580) );
  NAND2_X1 U677 ( .A1(n712), .A2(n580), .ZN(n581) );
  NAND2_X1 U678 ( .A1(n582), .A2(n607), .ZN(n583) );
  AND2_X1 U679 ( .A1(n584), .A2(n699), .ZN(n585) );
  AND2_X1 U680 ( .A1(n606), .A2(n585), .ZN(n586) );
  NAND2_X1 U681 ( .A1(n586), .A2(n607), .ZN(n642) );
  XNOR2_X1 U682 ( .A(n611), .B(KEYINPUT86), .ZN(n587) );
  NAND2_X1 U683 ( .A1(n757), .A2(n587), .ZN(n589) );
  NOR2_X1 U684 ( .A1(KEYINPUT65), .A2(KEYINPUT44), .ZN(n588) );
  NAND2_X1 U685 ( .A1(n589), .A2(n588), .ZN(n593) );
  OR2_X1 U686 ( .A1(n611), .A2(KEYINPUT65), .ZN(n590) );
  AND2_X1 U687 ( .A1(n590), .A2(KEYINPUT44), .ZN(n591) );
  NAND2_X1 U688 ( .A1(n757), .A2(n591), .ZN(n592) );
  NAND2_X1 U689 ( .A1(n593), .A2(n592), .ZN(n615) );
  XNOR2_X1 U690 ( .A(n596), .B(KEYINPUT96), .ZN(n597) );
  NAND2_X1 U691 ( .A1(n597), .A2(n699), .ZN(n598) );
  NAND2_X1 U692 ( .A1(n706), .A2(n600), .ZN(n601) );
  XNOR2_X1 U693 ( .A(KEYINPUT102), .B(n602), .ZN(n610) );
  AND2_X1 U694 ( .A1(n604), .A2(n603), .ZN(n605) );
  AND2_X1 U695 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U696 ( .A1(n608), .A2(n607), .ZN(n670) );
  INV_X1 U697 ( .A(n670), .ZN(n609) );
  NOR2_X1 U698 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U699 ( .A1(n611), .A2(KEYINPUT65), .ZN(n612) );
  AND2_X1 U700 ( .A1(n613), .A2(n612), .ZN(n614) );
  INV_X1 U701 ( .A(KEYINPUT83), .ZN(n616) );
  XNOR2_X1 U702 ( .A(n616), .B(KEYINPUT45), .ZN(n617) );
  AND2_X1 U703 ( .A1(KEYINPUT82), .A2(n620), .ZN(n619) );
  INV_X1 U704 ( .A(KEYINPUT2), .ZN(n621) );
  OR2_X1 U705 ( .A1(n618), .A2(n621), .ZN(n622) );
  INV_X1 U706 ( .A(n627), .ZN(n628) );
  XNOR2_X1 U707 ( .A(n629), .B(n628), .ZN(n632) );
  INV_X1 U708 ( .A(G952), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n630), .A2(G953), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n401), .ZN(n634) );
  XNOR2_X1 U711 ( .A(n634), .B(n633), .ZN(G66) );
  XOR2_X1 U712 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n638) );
  XNOR2_X1 U713 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U714 ( .A(G110), .B(KEYINPUT112), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n642), .B(n641), .ZN(G12) );
  XNOR2_X1 U716 ( .A(G119), .B(KEYINPUT127), .ZN(n644) );
  XOR2_X1 U717 ( .A(n644), .B(n643), .Z(G21) );
  XOR2_X1 U718 ( .A(G140), .B(n645), .Z(G42) );
  XOR2_X1 U719 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n646) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n649), .B(n648), .ZN(n650) );
  XOR2_X1 U722 ( .A(KEYINPUT119), .B(KEYINPUT56), .Z(n651) );
  XNOR2_X1 U723 ( .A(n652), .B(n651), .ZN(G51) );
  AND2_X1 U724 ( .A1(n653), .A2(n750), .ZN(n658) );
  NAND2_X1 U725 ( .A1(G953), .A2(G224), .ZN(n654) );
  XOR2_X1 U726 ( .A(KEYINPUT61), .B(n654), .Z(n655) );
  NOR2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U729 ( .A1(n659), .A2(n660), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n662), .B(n661), .ZN(G69) );
  XNOR2_X1 U731 ( .A(KEYINPUT66), .B(KEYINPUT59), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U734 ( .A(KEYINPUT121), .B(KEYINPUT60), .Z(n668) );
  XNOR2_X1 U735 ( .A(n669), .B(n668), .ZN(G60) );
  XNOR2_X1 U736 ( .A(G101), .B(KEYINPUT110), .ZN(n671) );
  XNOR2_X1 U737 ( .A(n671), .B(n670), .ZN(G3) );
  INV_X1 U738 ( .A(n682), .ZN(n686) );
  NOR2_X1 U739 ( .A1(n672), .A2(n686), .ZN(n673) );
  XOR2_X1 U740 ( .A(G104), .B(n673), .Z(G6) );
  NOR2_X1 U741 ( .A1(n689), .A2(n672), .ZN(n677) );
  XOR2_X1 U742 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n675) );
  XNOR2_X1 U743 ( .A(G107), .B(KEYINPUT111), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U745 ( .A(n677), .B(n676), .ZN(G9) );
  XOR2_X1 U746 ( .A(G128), .B(KEYINPUT29), .Z(n680) );
  INV_X1 U747 ( .A(n689), .ZN(n678) );
  NAND2_X1 U748 ( .A1(n683), .A2(n678), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n680), .B(n679), .ZN(G30) );
  XNOR2_X1 U750 ( .A(G143), .B(n681), .ZN(G45) );
  XOR2_X1 U751 ( .A(G146), .B(KEYINPUT113), .Z(n685) );
  NAND2_X1 U752 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U753 ( .A(n685), .B(n684), .ZN(G48) );
  NOR2_X1 U754 ( .A1(n686), .A2(n688), .ZN(n687) );
  XOR2_X1 U755 ( .A(G113), .B(n687), .Z(G15) );
  NOR2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U757 ( .A(G116), .B(n690), .Z(G18) );
  XNOR2_X1 U758 ( .A(G125), .B(n691), .ZN(n692) );
  XNOR2_X1 U759 ( .A(n692), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U760 ( .A(G134), .B(KEYINPUT114), .ZN(n694) );
  XNOR2_X1 U761 ( .A(n694), .B(n693), .ZN(G36) );
  NAND2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U763 ( .A(KEYINPUT49), .B(n697), .Z(n698) );
  NAND2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n704) );
  XNOR2_X1 U765 ( .A(n702), .B(KEYINPUT50), .ZN(n703) );
  NOR2_X1 U766 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U767 ( .A(KEYINPUT51), .B(n350), .Z(n707) );
  NOR2_X1 U768 ( .A1(n722), .A2(n707), .ZN(n708) );
  NAND2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U770 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U771 ( .A(KEYINPUT117), .B(n713), .Z(n716) );
  NAND2_X1 U772 ( .A1(n431), .A2(n714), .ZN(n715) );
  NAND2_X1 U773 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U774 ( .A1(n723), .A2(n717), .ZN(n718) );
  XOR2_X1 U775 ( .A(KEYINPUT52), .B(n719), .Z(n720) );
  NOR2_X1 U776 ( .A1(n721), .A2(n720), .ZN(n726) );
  XNOR2_X1 U777 ( .A(n626), .B(KEYINPUT2), .ZN(n725) );
  INV_X1 U778 ( .A(n722), .ZN(n724) );
  XNOR2_X1 U779 ( .A(KEYINPUT53), .B(n728), .ZN(G75) );
  NAND2_X1 U780 ( .A1(n735), .A2(G469), .ZN(n733) );
  XOR2_X1 U781 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n731) );
  XNOR2_X1 U782 ( .A(n729), .B(KEYINPUT120), .ZN(n730) );
  XNOR2_X1 U783 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U784 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U785 ( .A1(n739), .A2(n734), .ZN(G54) );
  NAND2_X1 U786 ( .A1(n735), .A2(G478), .ZN(n737) );
  XNOR2_X1 U787 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U788 ( .A1(n739), .A2(n738), .ZN(G63) );
  INV_X1 U789 ( .A(n740), .ZN(n744) );
  XNOR2_X1 U790 ( .A(n742), .B(n741), .ZN(n743) );
  XNOR2_X1 U791 ( .A(n743), .B(KEYINPUT123), .ZN(n747) );
  XOR2_X1 U792 ( .A(n744), .B(n747), .Z(n745) );
  XNOR2_X1 U793 ( .A(KEYINPUT124), .B(n745), .ZN(n746) );
  NOR2_X1 U794 ( .A1(G953), .A2(n746), .ZN(n753) );
  XNOR2_X1 U795 ( .A(n747), .B(G227), .ZN(n748) );
  XNOR2_X1 U796 ( .A(n748), .B(KEYINPUT125), .ZN(n749) );
  NAND2_X1 U797 ( .A1(n749), .A2(G900), .ZN(n751) );
  NOR2_X1 U798 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U799 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U800 ( .A(KEYINPUT126), .B(n754), .ZN(G72) );
  XOR2_X1 U801 ( .A(n755), .B(G137), .Z(G39) );
  XOR2_X1 U802 ( .A(n756), .B(G131), .Z(G33) );
  XNOR2_X1 U803 ( .A(n757), .B(G122), .ZN(G24) );
endmodule

