//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n607, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT65), .Z(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  XOR2_X1   g032(.A(G325), .B(KEYINPUT67), .Z(G261));
  AOI22_X1  g033(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G137), .ZN(new_n465));
  NAND2_X1  g040(.A1(G101), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n464), .A2(new_n467), .ZN(G160));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(new_n460), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(new_n460), .B2(G112), .ZN(new_n478));
  NOR2_X1   g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT68), .Z(new_n480));
  OAI211_X1 g055(.A(new_n475), .B(new_n477), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  INV_X1    g057(.A(KEYINPUT72), .ZN(new_n483));
  OR2_X1    g058(.A1(KEYINPUT69), .A2(G114), .ZN(new_n484));
  NAND2_X1  g059(.A1(KEYINPUT69), .A2(G114), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n484), .A2(G2105), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n486), .A2(KEYINPUT70), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(KEYINPUT70), .B1(new_n486), .B2(new_n488), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n461), .A2(G126), .A3(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n460), .A2(KEYINPUT71), .A3(G138), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n473), .A2(KEYINPUT4), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n460), .A2(KEYINPUT71), .A3(G138), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n495), .B1(new_n461), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n492), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n483), .B1(new_n491), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT4), .B1(new_n473), .B2(new_n493), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n461), .A2(new_n495), .A3(new_n496), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n500), .A2(new_n501), .B1(new_n476), .B2(G126), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT69), .A2(G114), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT69), .A2(G114), .ZN(new_n505));
  NOR3_X1   g080(.A1(new_n504), .A2(new_n505), .A3(new_n460), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n503), .B1(new_n506), .B2(new_n487), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n486), .A2(KEYINPUT70), .A3(new_n488), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n502), .A2(new_n509), .A3(KEYINPUT72), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n499), .A2(new_n510), .ZN(G164));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n520), .B(new_n522), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n517), .A2(new_n518), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n515), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  AOI22_X1  g104(.A1(new_n516), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n516), .A2(G543), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n531), .A2(new_n512), .B1(new_n532), .B2(G51), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(new_n532), .A2(G52), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OAI221_X1 g115(.A(new_n538), .B1(new_n539), .B2(new_n525), .C1(new_n514), .C2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n542), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(G171));
  AOI22_X1  g120(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n514), .ZN(new_n547));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n517), .A2(new_n548), .B1(new_n525), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n532), .A2(G53), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n512), .A2(G65), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n514), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n525), .B(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n562), .B1(new_n564), .B2(G91), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n559), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  NOR2_X1   g142(.A1(new_n525), .A2(new_n563), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT74), .B1(new_n512), .B2(new_n516), .ZN(new_n569));
  OAI21_X1  g144(.A(G87), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT75), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n512), .A2(G74), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G651), .B1(new_n532), .B2(G49), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n574), .B(G87), .C1(new_n568), .C2(new_n569), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n571), .A2(new_n573), .A3(new_n575), .ZN(G288));
  AOI22_X1  g151(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G48), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n577), .A2(new_n514), .B1(new_n578), .B2(new_n517), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(G86), .B2(new_n564), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n514), .ZN(new_n583));
  INV_X1    g158(.A(G47), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n517), .A2(new_n584), .B1(new_n525), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(new_n564), .A2(G92), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n520), .A2(new_n522), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(new_n532), .B2(G54), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n589), .A2(KEYINPUT10), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n590), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n598), .B2(G171), .ZN(G284));
  OAI21_X1  g175(.A(new_n599), .B1(new_n598), .B2(G171), .ZN(G321));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  INV_X1    g177(.A(G299), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G297));
  XOR2_X1   g179(.A(G297), .B(KEYINPUT76), .Z(G280));
  INV_X1    g180(.A(new_n597), .ZN(new_n606));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G860), .ZN(G148));
  INV_X1    g183(.A(new_n551), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(new_n598), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n597), .A2(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(new_n598), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n474), .A2(G2104), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2100), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n476), .A2(G123), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT77), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n474), .A2(G135), .ZN(new_n621));
  OR2_X1    g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n622), .B(G2104), .C1(G111), .C2(new_n460), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n476), .A2(KEYINPUT77), .A3(G123), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n620), .A2(new_n621), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G2096), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n617), .A2(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT78), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2430), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT14), .ZN(new_n634));
  XOR2_X1   g209(.A(G2451), .B(G2454), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n634), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2443), .B(G2446), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n641), .A2(G14), .ZN(G401));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT79), .ZN(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  AND2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT80), .Z(new_n650));
  OR2_X1    g225(.A1(new_n650), .A2(KEYINPUT18), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n646), .B1(KEYINPUT17), .B2(new_n648), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n644), .A2(new_n645), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT17), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n653), .B1(new_n654), .B2(new_n647), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n647), .B(KEYINPUT81), .Z(new_n656));
  AOI22_X1  g231(.A1(new_n652), .A2(new_n655), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n650), .A2(KEYINPUT18), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n651), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT82), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(new_n626), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(G2100), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n675), .C1(new_n673), .C2(new_n672), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(G1986), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1991), .B(G1996), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT83), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT22), .B(G1981), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  NOR2_X1   g258(.A1(G16), .A2(G23), .ZN(new_n684));
  INV_X1    g259(.A(G288), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(G16), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT33), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G22), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n689), .ZN(new_n691));
  INV_X1    g266(.A(G1971), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n689), .A2(G6), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(new_n580), .B2(new_n689), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT32), .B(G1981), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n688), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT34), .Z(new_n699));
  INV_X1    g274(.A(KEYINPUT84), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n689), .A2(G24), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n587), .B2(new_n689), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1986), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n476), .A2(G119), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n474), .A2(G131), .ZN(new_n705));
  NOR2_X1   g280(.A1(G95), .A2(G2105), .ZN(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(new_n460), .B2(G107), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n704), .B(new_n705), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  MUX2_X1   g283(.A(G25), .B(new_n708), .S(G29), .Z(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT35), .B(G1991), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n703), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n699), .A2(new_n700), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n699), .A2(new_n713), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(KEYINPUT85), .ZN(new_n716));
  OAI211_X1 g291(.A(KEYINPUT36), .B(new_n714), .C1(new_n716), .C2(new_n700), .ZN(new_n717));
  NOR2_X1   g292(.A1(G171), .A2(new_n689), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G5), .B2(new_n689), .ZN(new_n719));
  INV_X1    g294(.A(G1961), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G32), .ZN(new_n722));
  NAND2_X1  g297(.A1(G105), .A2(G2104), .ZN(new_n723));
  INV_X1    g298(.A(G141), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n473), .B2(new_n724), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n725), .A2(new_n460), .B1(new_n476), .B2(G129), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n722), .B1(new_n731), .B2(new_n721), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT93), .Z(new_n733));
  XOR2_X1   g308(.A(KEYINPUT27), .B(G1996), .Z(new_n734));
  AOI22_X1  g309(.A1(new_n719), .A2(new_n720), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT29), .B(G2090), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n721), .A2(G35), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n721), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT96), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n735), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G16), .A2(G21), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G168), .B2(G16), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(G1966), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT28), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n721), .A2(G26), .ZN(new_n745));
  AOI22_X1  g320(.A1(G128), .A2(new_n476), .B1(new_n474), .B2(G140), .ZN(new_n746));
  OAI21_X1  g321(.A(G2104), .B1(new_n460), .B2(G116), .ZN(new_n747));
  NOR2_X1   g322(.A1(G104), .A2(G2105), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT86), .Z(new_n749));
  OAI21_X1  g324(.A(new_n746), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  AOI211_X1 g325(.A(new_n744), .B(new_n745), .C1(new_n750), .C2(G29), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n744), .B2(new_n745), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT87), .B(G2067), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT88), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n752), .B(new_n754), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n689), .A2(KEYINPUT23), .A3(G20), .ZN(new_n756));
  AOI21_X1  g331(.A(KEYINPUT23), .B1(new_n689), .B2(G20), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n756), .B(new_n757), .C1(G299), .C2(G16), .ZN(new_n758));
  INV_X1    g333(.A(G1956), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n740), .A2(new_n743), .A3(new_n755), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n739), .A2(new_n736), .ZN(new_n762));
  INV_X1    g337(.A(G34), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n763), .A2(KEYINPUT24), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(KEYINPUT24), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n721), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G160), .B2(new_n721), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G2084), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G11), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n762), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G19), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n551), .B2(G16), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n770), .B1(G1341), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n719), .A2(new_n720), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n733), .A2(new_n734), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n625), .A2(new_n721), .ZN(new_n776));
  INV_X1    g351(.A(G28), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(KEYINPUT30), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT94), .ZN(new_n779));
  AOI211_X1 g354(.A(G29), .B(new_n779), .C1(KEYINPUT30), .C2(new_n777), .ZN(new_n780));
  NOR4_X1   g355(.A1(new_n774), .A2(new_n775), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n717), .A2(new_n761), .A3(new_n773), .A4(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n767), .A2(G2084), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT95), .Z(new_n784));
  NOR2_X1   g359(.A1(G4), .A2(G16), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n606), .B2(G16), .ZN(new_n786));
  NOR2_X1   g361(.A1(G29), .A2(G33), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT25), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n474), .A2(G139), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT89), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT90), .Z(new_n794));
  OAI21_X1  g369(.A(new_n792), .B1(new_n460), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT91), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n787), .B1(new_n796), .B2(G29), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n784), .B1(G1348), .B2(new_n786), .C1(new_n797), .C2(G2072), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n742), .A2(G1966), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n782), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n797), .A2(G2072), .B1(G1348), .B2(new_n786), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n772), .A2(G1341), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n716), .A2(KEYINPUT36), .ZN(new_n804));
  NOR2_X1   g379(.A1(G27), .A2(G29), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G164), .B2(G29), .ZN(new_n806));
  INV_X1    g381(.A(G2078), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n802), .A2(new_n803), .A3(new_n804), .A4(new_n808), .ZN(G150));
  INV_X1    g384(.A(G150), .ZN(G311));
  AOI22_X1  g385(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT97), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(new_n514), .ZN(new_n813));
  INV_X1    g388(.A(G55), .ZN(new_n814));
  INV_X1    g389(.A(G93), .ZN(new_n815));
  OAI22_X1  g390(.A1(new_n517), .A2(new_n814), .B1(new_n525), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT99), .B(G860), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT37), .Z(new_n821));
  NOR2_X1   g396(.A1(new_n597), .A2(new_n607), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT38), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT39), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n551), .B1(new_n818), .B2(KEYINPUT98), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n818), .A2(KEYINPUT98), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n825), .B(new_n826), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n824), .B(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n821), .B1(new_n828), .B2(new_n819), .ZN(G145));
  XNOR2_X1  g404(.A(new_n796), .B(new_n731), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT100), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n491), .A2(new_n498), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(KEYINPUT100), .B1(new_n502), .B2(new_n509), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n708), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n830), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n625), .B(G160), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G162), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n476), .A2(G130), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n474), .A2(G142), .ZN(new_n840));
  NOR2_X1   g415(.A1(G106), .A2(G2105), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(new_n460), .B2(G118), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n839), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n750), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n615), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n838), .B(new_n845), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n836), .B(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(G37), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT40), .Z(G395));
  NAND2_X1  g424(.A1(new_n818), .A2(new_n598), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n827), .B(new_n611), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n597), .B(G299), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT101), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n606), .A2(G299), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(KEYINPUT101), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT41), .ZN(new_n857));
  INV_X1    g432(.A(new_n852), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n855), .A2(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n851), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n855), .B2(new_n851), .ZN(new_n862));
  XNOR2_X1  g437(.A(G303), .B(new_n587), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n685), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n580), .B(KEYINPUT103), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT42), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n862), .B(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n850), .B1(new_n868), .B2(new_n598), .ZN(G295));
  OAI21_X1  g444(.A(new_n850), .B1(new_n868), .B2(new_n598), .ZN(G331));
  XNOR2_X1  g445(.A(G171), .B(G286), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n827), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(new_n855), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n860), .B2(new_n872), .ZN(new_n874));
  AOI21_X1  g449(.A(G37), .B1(new_n874), .B2(new_n866), .ZN(new_n875));
  INV_X1    g450(.A(new_n872), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n855), .B1(new_n876), .B2(new_n856), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n872), .A2(new_n857), .A3(new_n858), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n875), .B1(new_n879), .B2(new_n866), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT43), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT104), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n874), .A2(new_n866), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n884), .A2(new_n875), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n880), .A2(KEYINPUT43), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(new_n886), .B2(new_n885), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n883), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(G397));
  NOR2_X1   g467(.A1(new_n750), .A2(G2067), .ZN(new_n893));
  INV_X1    g468(.A(G1384), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n832), .B2(new_n833), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT45), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(G40), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n464), .A2(new_n467), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G1996), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OR3_X1    g478(.A1(new_n903), .A2(KEYINPUT105), .A3(new_n730), .ZN(new_n904));
  INV_X1    g479(.A(G2067), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n750), .B(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n902), .B2(new_n731), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT105), .B1(new_n903), .B2(new_n730), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n904), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT106), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n708), .A2(new_n710), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT125), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n893), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT126), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n917), .A3(new_n901), .ZN(new_n918));
  INV_X1    g493(.A(new_n903), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n919), .A2(KEYINPUT46), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(KEYINPUT46), .ZN(new_n921));
  INV_X1    g496(.A(new_n906), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n901), .B1(new_n730), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT47), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n708), .B(new_n710), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n901), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n911), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(G290), .A2(G1986), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n901), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT48), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n918), .A2(new_n925), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT123), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n831), .B1(new_n491), .B2(new_n498), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n502), .A2(new_n509), .A3(KEYINPUT100), .ZN(new_n936));
  AOI21_X1  g511(.A(G1384), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n900), .B1(new_n937), .B2(KEYINPUT45), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n499), .A2(new_n894), .A3(new_n510), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n896), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n807), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT53), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(G2078), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n895), .B2(new_n896), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n946), .A2(KEYINPUT122), .A3(new_n938), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT122), .B1(new_n946), .B2(new_n938), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n943), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n939), .A2(KEYINPUT50), .ZN(new_n950));
  AOI21_X1  g525(.A(G1384), .B1(new_n502), .B2(new_n509), .ZN(new_n951));
  XOR2_X1   g526(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n900), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT114), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT114), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n950), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n720), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT121), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n950), .A2(new_n954), .A3(new_n957), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n957), .B1(new_n950), .B2(new_n954), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(KEYINPUT121), .A3(new_n720), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n949), .B1(new_n961), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT54), .B1(new_n966), .B2(G301), .ZN(new_n967));
  INV_X1    g542(.A(new_n943), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT120), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n962), .A2(new_n963), .A3(G1961), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n894), .B1(new_n491), .B2(new_n498), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n896), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n972), .B(new_n899), .C1(new_n939), .C2(new_n896), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(new_n945), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n969), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n974), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n959), .A2(KEYINPUT120), .A3(new_n976), .ZN(new_n977));
  AOI211_X1 g552(.A(G171), .B(new_n968), .C1(new_n975), .C2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n934), .B1(new_n967), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n977), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(G301), .A3(new_n943), .ZN(new_n981));
  INV_X1    g556(.A(new_n948), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n946), .A2(new_n938), .A3(KEYINPUT122), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n982), .A2(new_n983), .B1(new_n942), .B2(new_n941), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n970), .A2(KEYINPUT121), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n959), .A2(new_n960), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(G171), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n981), .A2(new_n988), .A3(KEYINPUT123), .A4(KEYINPUT54), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n979), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT119), .ZN(new_n991));
  NAND2_X1  g566(.A1(G286), .A2(G8), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n992), .B(KEYINPUT117), .Z(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G8), .ZN(new_n995));
  INV_X1    g570(.A(G1966), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n973), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G2084), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n950), .A2(new_n954), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n995), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n994), .B1(new_n1000), .B2(KEYINPUT118), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1000), .A2(KEYINPUT118), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n991), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT51), .B1(new_n1000), .B2(new_n994), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1004), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1007), .A2(KEYINPUT119), .A3(new_n1002), .A4(new_n1001), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n997), .A2(new_n999), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n994), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n499), .A2(new_n1013), .A3(new_n894), .A4(new_n510), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n971), .A2(new_n952), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(new_n1015), .A3(new_n899), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n759), .ZN(new_n1017));
  OAI211_X1 g592(.A(KEYINPUT45), .B(new_n894), .C1(new_n832), .C2(new_n833), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT56), .B(G2072), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n940), .A2(new_n1018), .A3(new_n899), .A4(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n1021));
  XNOR2_X1  g596(.A(G299), .B(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1017), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1348), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n964), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n951), .A2(new_n899), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(G2067), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n597), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1022), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1023), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT115), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1033), .B(new_n1023), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1022), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(KEYINPUT61), .A3(new_n1023), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n938), .A2(new_n902), .A3(new_n940), .ZN(new_n1039));
  XOR2_X1   g614(.A(KEYINPUT58), .B(G1341), .Z(new_n1040));
  NAND2_X1  g615(.A1(new_n1026), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n609), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1037), .A2(new_n1023), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT61), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1017), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1045), .B(new_n1047), .C1(new_n1049), .C2(new_n1030), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1038), .B(new_n1044), .C1(new_n1048), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n606), .A2(KEYINPUT60), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n606), .A2(KEYINPUT60), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1025), .A2(new_n1028), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1032), .B(new_n1034), .C1(new_n1052), .C2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1981), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G73), .A2(G543), .ZN(new_n1061));
  INV_X1    g636(.A(G61), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n592), .B2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1063), .A2(G651), .B1(new_n532), .B2(G48), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT110), .B(G86), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n512), .A2(new_n516), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1060), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n580), .B2(new_n1060), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT49), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n1070));
  AOI211_X1 g645(.A(G1981), .B(new_n579), .C1(G86), .C2(new_n564), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(new_n1067), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n995), .B1(new_n951), .B2(new_n899), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n571), .A2(G1976), .A3(new_n573), .A4(new_n575), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(KEYINPUT109), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1976), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1026), .A2(G288), .A3(G8), .A4(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1076), .B1(new_n1079), .B2(new_n1078), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1074), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1018), .A2(new_n899), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n939), .A2(new_n896), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n692), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G2090), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n950), .A2(new_n954), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n995), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(G303), .A2(G8), .ZN(new_n1090));
  XOR2_X1   g665(.A(new_n1090), .B(KEYINPUT55), .Z(new_n1091));
  AOI21_X1  g666(.A(new_n1083), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1014), .A2(new_n1015), .A3(new_n899), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1087), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n995), .B1(new_n1086), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT111), .B1(new_n1095), .B2(new_n1091), .ZN(new_n1096));
  AOI21_X1  g671(.A(G1971), .B1(new_n938), .B2(new_n940), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1016), .A2(G2090), .ZN(new_n1098));
  OAI21_X1  g673(.A(G8), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT111), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1091), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1092), .A2(new_n1096), .A3(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n984), .B(G301), .C1(new_n985), .C2(new_n986), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n968), .B1(new_n975), .B2(new_n977), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(G301), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1103), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n990), .A2(new_n1012), .A3(new_n1059), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1074), .A2(new_n1077), .A3(new_n685), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(G1981), .B2(G305), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n1073), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1088), .ZN(new_n1114));
  OAI211_X1 g689(.A(G8), .B(new_n1091), .C1(new_n1097), .C2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1113), .B1(new_n1115), .B2(new_n1083), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1000), .A2(G168), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1092), .A2(new_n1118), .A3(new_n1096), .A4(new_n1102), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT112), .B(KEYINPUT63), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT63), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1069), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1124), .A2(KEYINPUT109), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1123), .B1(new_n1125), .B2(new_n1080), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1115), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1128), .A2(new_n1118), .ZN(new_n1129));
  OAI211_X1 g704(.A(KEYINPUT113), .B(new_n1117), .C1(new_n1121), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT113), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1119), .A2(new_n1120), .B1(new_n1128), .B2(new_n1118), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1132), .B2(new_n1116), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1109), .A2(new_n1110), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1110), .B1(new_n1109), .B2(new_n1134), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1103), .B1(new_n1012), .B2(KEYINPUT62), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1009), .A2(new_n1138), .A3(new_n1011), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1105), .A2(G301), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1135), .A2(new_n1136), .A3(new_n1141), .ZN(new_n1142));
  AND2_X1   g717(.A1(G290), .A2(G1986), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n901), .B1(new_n929), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n928), .A2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT107), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n933), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n933), .B(KEYINPUT127), .C1(new_n1142), .C2(new_n1146), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g726(.A1(new_n848), .A2(G401), .A3(G229), .ZN(new_n1153));
  NAND4_X1  g727(.A1(new_n890), .A2(G319), .A3(new_n662), .A4(new_n1153), .ZN(G225));
  INV_X1    g728(.A(G225), .ZN(G308));
endmodule


