//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n212), .B(new_n217), .C1(G107), .C2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G116), .A2(G270), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n206), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n204), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT64), .ZN(new_n233));
  OAI21_X1  g0033(.A(G50), .B1(G58), .B2(G68), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n209), .B(new_n230), .C1(new_n233), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n252), .B(new_n231), .C1(G1), .C2(new_n204), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(new_n221), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G13), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n256), .A2(new_n204), .A3(G1), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G50), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR3_X1   g0063(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n261), .A2(new_n263), .B1(new_n264), .B2(new_n204), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n226), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT8), .B(G58), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(KEYINPUT66), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n204), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n265), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n252), .A2(new_n231), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n255), .B(new_n260), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT70), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT66), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT8), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n278), .A3(G58), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n226), .A2(KEYINPUT8), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n270), .B(new_n279), .C1(new_n282), .C2(new_n277), .ZN(new_n283));
  INV_X1    g0083(.A(new_n264), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n284), .A2(G20), .B1(G150), .B2(new_n262), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n259), .B1(new_n286), .B2(new_n272), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(KEYINPUT70), .A3(new_n255), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n276), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G1), .A3(G13), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT65), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n291), .A2(KEYINPUT65), .A3(new_n292), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G226), .ZN(new_n298));
  OR2_X1    g0098(.A1(KEYINPUT3), .A2(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(KEYINPUT3), .A2(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G1698), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G222), .ZN(new_n303));
  INV_X1    g0103(.A(G223), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n301), .B(new_n303), .C1(new_n304), .C2(new_n302), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n305), .B(new_n306), .C1(G77), .C2(new_n301), .ZN(new_n307));
  INV_X1    g0107(.A(G274), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n292), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n298), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n289), .A2(KEYINPUT9), .B1(G190), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT9), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n276), .A2(new_n288), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n311), .A2(G200), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n313), .A2(new_n314), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT70), .B1(new_n287), .B2(new_n255), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n273), .B1(new_n283), .B2(new_n285), .ZN(new_n320));
  NOR4_X1   g0120(.A1(new_n320), .A2(new_n275), .A3(new_n254), .A4(new_n259), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT9), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n312), .A2(G190), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n322), .A2(new_n323), .A3(new_n316), .A4(new_n317), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT10), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n312), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n311), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n274), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n309), .B1(new_n297), .B2(G244), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n302), .A2(G232), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n301), .B(new_n336), .C1(new_n211), .C2(new_n302), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(G107), .B2(new_n301), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n335), .B1(new_n291), .B2(new_n338), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n339), .A2(G200), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n257), .A2(new_n223), .ZN(new_n341));
  XOR2_X1   g0141(.A(new_n341), .B(KEYINPUT68), .Z(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT15), .B(G87), .Z(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n344), .A2(new_n269), .B1(new_n204), .B2(new_n223), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n267), .B(KEYINPUT67), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(new_n262), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n342), .B1(new_n223), .B2(new_n253), .C1(new_n347), .C2(new_n273), .ZN(new_n348));
  INV_X1    g0148(.A(G190), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n339), .A2(new_n349), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n340), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n339), .A2(G179), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n339), .A2(new_n330), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(new_n348), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n356), .A2(KEYINPUT69), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(KEYINPUT69), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n334), .A2(new_n357), .A3(KEYINPUT71), .A4(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT16), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n299), .A2(new_n204), .A3(new_n300), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT7), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(KEYINPUT3), .A2(G33), .ZN(new_n364));
  NOR2_X1   g0164(.A1(KEYINPUT3), .A2(G33), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n210), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n226), .A2(new_n210), .ZN(new_n369));
  NOR2_X1   g0169(.A1(G58), .A2(G68), .ZN(new_n370));
  OAI21_X1  g0170(.A(G20), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n262), .A2(G159), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n360), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT7), .B1(new_n366), .B2(new_n204), .ZN(new_n375));
  NOR4_X1   g0175(.A1(new_n364), .A2(new_n365), .A3(new_n362), .A4(G20), .ZN(new_n376));
  OAI21_X1  g0176(.A(G68), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n373), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(KEYINPUT16), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n374), .A2(new_n379), .A3(new_n272), .ZN(new_n380));
  INV_X1    g0180(.A(new_n268), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n381), .A2(new_n253), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n257), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n304), .A2(new_n302), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n301), .B(new_n385), .C1(G226), .C2(new_n302), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n309), .B1(new_n388), .B2(new_n306), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n293), .A2(new_n227), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G200), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(G190), .A3(new_n391), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n384), .A2(KEYINPUT17), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT17), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n380), .A2(new_n394), .A3(new_n382), .A4(new_n383), .ZN(new_n397));
  INV_X1    g0197(.A(new_n393), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n395), .A2(KEYINPUT75), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT75), .B1(new_n395), .B2(new_n399), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n291), .B1(new_n386), .B2(new_n387), .ZN(new_n402));
  NOR4_X1   g0202(.A1(new_n402), .A2(G179), .A3(new_n309), .A4(new_n390), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n330), .B2(new_n392), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n404), .A2(new_n405), .A3(KEYINPUT18), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT18), .B1(new_n404), .B2(new_n405), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n400), .A2(new_n401), .A3(new_n408), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n359), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT14), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n291), .A2(KEYINPUT65), .A3(new_n292), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT65), .B1(new_n291), .B2(new_n292), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT73), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT73), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n295), .A2(new_n415), .A3(new_n296), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n416), .A3(G238), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n222), .A2(new_n302), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n227), .A2(G1698), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n418), .B(new_n419), .C1(new_n364), .C2(new_n365), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G97), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT72), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT72), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n420), .A2(new_n424), .A3(new_n421), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n306), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n417), .A2(new_n310), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT13), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n417), .A2(new_n426), .A3(new_n429), .A4(new_n310), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n411), .B1(new_n431), .B2(G169), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI211_X1 g0233(.A(KEYINPUT14), .B(new_n330), .C1(new_n428), .C2(new_n430), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n431), .A2(new_n328), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n263), .A2(new_n221), .B1(new_n204), .B2(G68), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n269), .A2(new_n223), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n272), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  XOR2_X1   g0241(.A(KEYINPUT74), .B(KEYINPUT11), .Z(new_n442));
  XNOR2_X1  g0242(.A(new_n441), .B(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n253), .A2(new_n210), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n257), .A2(new_n210), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT12), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n445), .B(new_n446), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n443), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n438), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n431), .A2(G200), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n451), .B(new_n448), .C1(new_n349), .C2(new_n431), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n334), .A2(new_n357), .A3(new_n358), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT71), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n410), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT24), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n204), .B(G87), .C1(new_n364), .C2(new_n365), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT22), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT22), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n301), .A2(new_n462), .A3(new_n204), .A4(G87), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT82), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G116), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G20), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT23), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n204), .B2(G107), .ZN(new_n469));
  INV_X1    g0269(.A(G107), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(KEYINPUT23), .A3(G20), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n467), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n464), .A2(new_n465), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n465), .B1(new_n464), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n459), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n464), .A2(new_n472), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT82), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(KEYINPUT24), .A3(new_n473), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n476), .A2(new_n479), .A3(new_n272), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT25), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n258), .B2(G107), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n257), .A2(KEYINPUT25), .A3(new_n470), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n203), .A2(G33), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(new_n231), .A3(new_n252), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(new_n257), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n482), .A2(new_n483), .B1(G107), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G41), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n203), .B(G45), .C1(new_n489), .C2(KEYINPUT5), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT5), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(G41), .ZN(new_n492));
  OAI211_X1 g0292(.A(G264), .B(new_n291), .C1(new_n490), .C2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n214), .A2(new_n302), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n216), .A2(G1698), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(new_n496), .C1(new_n364), .C2(new_n365), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G294), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n497), .A2(KEYINPUT83), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT83), .B1(new_n497), .B2(new_n498), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n494), .B1(new_n501), .B2(new_n306), .ZN(new_n502));
  OAI21_X1  g0302(.A(G274), .B1(new_n491), .B2(G41), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n306), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n490), .A2(KEYINPUT76), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT76), .ZN(new_n506));
  INV_X1    g0306(.A(G45), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(G1), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n491), .A2(G41), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n504), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT77), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n490), .A2(KEYINPUT76), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n508), .A2(new_n506), .A3(new_n509), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT77), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(new_n504), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(G169), .B1(new_n502), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n497), .A2(new_n498), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT83), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n497), .A2(KEYINPUT83), .A3(new_n498), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n306), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n493), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n515), .A2(new_n516), .A3(new_n504), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n516), .B1(new_n515), .B2(new_n504), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n526), .A2(new_n529), .A3(G179), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n488), .A2(new_n520), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n533), .B(new_n204), .C1(G33), .C2(new_n215), .ZN(new_n534));
  INV_X1    g0334(.A(G116), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G20), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n272), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT20), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n534), .A2(KEYINPUT20), .A3(new_n272), .A4(new_n536), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n539), .A2(new_n540), .B1(G116), .B2(new_n486), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n257), .A2(new_n535), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n330), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n302), .A2(G257), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G264), .A2(G1698), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n544), .B(new_n545), .C1(new_n364), .C2(new_n365), .ZN(new_n546));
  INV_X1    g0346(.A(G303), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n299), .A2(new_n547), .A3(new_n300), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n306), .A3(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(G270), .B(new_n291), .C1(new_n490), .C2(new_n492), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n549), .B(new_n550), .C1(new_n527), .C2(new_n528), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n543), .A2(new_n551), .A3(KEYINPUT21), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT21), .B1(new_n543), .B2(new_n551), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT81), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n518), .A2(G179), .A3(new_n549), .A4(new_n550), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n541), .A2(new_n542), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n555), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n551), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n560), .A2(KEYINPUT81), .A3(G179), .A4(new_n557), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n557), .B1(new_n560), .B2(G190), .ZN(new_n563));
  INV_X1    g0363(.A(G200), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n563), .B1(new_n564), .B2(new_n560), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n532), .A2(new_n554), .A3(new_n562), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n508), .A2(new_n308), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n214), .B1(new_n507), .B2(G1), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n291), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n224), .A2(G1698), .ZN(new_n570));
  OAI221_X1 g0370(.A(new_n570), .B1(G238), .B2(G1698), .C1(new_n364), .C2(new_n365), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n571), .A2(new_n466), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n569), .B1(new_n572), .B2(new_n291), .ZN(new_n573));
  OAI21_X1  g0373(.A(KEYINPUT80), .B1(new_n573), .B2(new_n349), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n291), .B1(new_n571), .B2(new_n466), .ZN(new_n575));
  INV_X1    g0375(.A(new_n569), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT80), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(new_n578), .A3(G190), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n301), .A2(new_n204), .A3(G68), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n213), .A2(new_n215), .A3(new_n470), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n421), .A2(new_n204), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT19), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n421), .B2(G20), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n581), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(new_n272), .B1(new_n257), .B2(new_n344), .ZN(new_n588));
  OAI21_X1  g0388(.A(G200), .B1(new_n575), .B2(new_n576), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n486), .A2(G87), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT79), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT79), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n588), .A2(new_n589), .A3(new_n593), .A4(new_n590), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n580), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n486), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n588), .B1(new_n344), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n577), .A2(new_n328), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n597), .B(new_n598), .C1(G169), .C2(new_n577), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n214), .B1(new_n299), .B2(new_n300), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT4), .ZN(new_n602));
  OAI21_X1  g0402(.A(G1698), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(G244), .B1(new_n364), .B2(new_n365), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n604), .A2(new_n602), .B1(G33), .B2(G283), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n301), .A2(KEYINPUT4), .A3(G244), .A4(new_n302), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n306), .ZN(new_n608));
  OAI211_X1 g0408(.A(G257), .B(new_n291), .C1(new_n490), .C2(new_n492), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT78), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n518), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n330), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n517), .A2(new_n512), .B1(new_n607), .B2(new_n306), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(new_n328), .A3(new_n611), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT6), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n616), .A2(new_n215), .A3(G107), .ZN(new_n617));
  XNOR2_X1  g0417(.A(G97), .B(G107), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n617), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI22_X1  g0419(.A1(new_n619), .A2(new_n204), .B1(new_n223), .B2(new_n263), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n470), .B1(new_n363), .B2(new_n367), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n272), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n486), .A2(G97), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n257), .A2(new_n215), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n613), .A2(new_n615), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n612), .A2(G200), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n614), .A2(G190), .A3(new_n611), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n502), .A2(new_n518), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G200), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n502), .A2(G190), .A3(new_n518), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n480), .A2(new_n632), .A3(new_n633), .A4(new_n487), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n600), .A2(new_n626), .A3(new_n630), .A4(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n458), .A2(new_n566), .A3(new_n635), .ZN(G372));
  AND3_X1   g0436(.A1(new_n562), .A2(KEYINPUT87), .A3(new_n554), .ZN(new_n637));
  AOI21_X1  g0437(.A(KEYINPUT87), .B1(new_n562), .B2(new_n554), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n532), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n575), .A2(KEYINPUT84), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT84), .ZN(new_n641));
  AOI211_X1 g0441(.A(new_n641), .B(new_n291), .C1(new_n571), .C2(new_n466), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n569), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n643), .A2(KEYINPUT85), .A3(new_n330), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT85), .B1(new_n643), .B2(new_n330), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n598), .B(new_n597), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n587), .A2(new_n272), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n344), .A2(new_n257), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n590), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT86), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n643), .A2(G200), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n580), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n480), .A2(new_n632), .A3(new_n633), .A4(new_n487), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n626), .A2(new_n630), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n639), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n626), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n646), .A2(new_n659), .A3(new_n660), .A4(new_n653), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n595), .A2(new_n599), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT26), .B1(new_n662), .B2(new_n626), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n661), .A2(new_n663), .A3(new_n646), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n457), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n450), .A2(new_n355), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT75), .ZN(new_n668));
  INV_X1    g0468(.A(new_n399), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n397), .A2(new_n398), .A3(new_n396), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n395), .A2(KEYINPUT75), .A3(new_n399), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n667), .A2(new_n452), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n408), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n333), .B1(new_n675), .B2(new_n326), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n666), .A2(new_n676), .ZN(G369));
  NOR2_X1   g0477(.A1(new_n256), .A2(G20), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n203), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n557), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT88), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n565), .A2(new_n562), .A3(new_n554), .A4(new_n686), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n637), .A2(new_n638), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n687), .B1(new_n688), .B2(new_n686), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n684), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n480), .B2(new_n487), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n532), .B1(new_n655), .B2(new_n693), .ZN(new_n694));
  AOI211_X1 g0494(.A(new_n519), .B(new_n530), .C1(new_n480), .C2(new_n487), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n692), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n684), .B1(new_n562), .B2(new_n554), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n700), .A2(new_n696), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n207), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n582), .A2(G116), .ZN(new_n706));
  XOR2_X1   g0506(.A(new_n706), .B(KEYINPUT89), .Z(new_n707));
  NAND3_X1  g0507(.A1(new_n705), .A2(new_n707), .A3(G1), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n234), .B2(new_n705), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n655), .A2(new_n656), .A3(new_n662), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n562), .A2(new_n554), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n695), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n711), .A2(new_n713), .A3(new_n565), .A4(new_n692), .ZN(new_n714));
  XNOR2_X1  g0514(.A(KEYINPUT91), .B(KEYINPUT30), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n614), .A2(new_n502), .A3(new_n611), .A4(new_n577), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT90), .B1(new_n716), .B2(new_n556), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n551), .A2(new_n328), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n518), .A2(new_n608), .A3(new_n611), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT90), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n526), .A2(new_n573), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n718), .A2(new_n719), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n715), .B1(new_n717), .B2(new_n722), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n643), .A2(new_n328), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n551), .A3(new_n631), .A4(new_n612), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n718), .A2(new_n719), .A3(KEYINPUT30), .A4(new_n721), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n684), .B1(new_n723), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g0530(.A(KEYINPUT31), .B(new_n684), .C1(new_n723), .C2(new_n727), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n714), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G330), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n684), .B1(new_n658), .B2(new_n664), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT29), .ZN(new_n736));
  NOR4_X1   g0536(.A1(new_n713), .A2(new_n656), .A3(new_n655), .A4(new_n654), .ZN(new_n737));
  OAI21_X1  g0537(.A(KEYINPUT26), .B1(new_n654), .B2(new_n626), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n600), .A2(new_n660), .A3(new_n659), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(new_n646), .A3(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(KEYINPUT29), .B(new_n692), .C1(new_n737), .C2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n734), .B1(new_n736), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n710), .B1(new_n742), .B2(G1), .ZN(G364));
  XOR2_X1   g0543(.A(new_n690), .B(KEYINPUT92), .Z(new_n744));
  AOI21_X1  g0544(.A(new_n203), .B1(new_n678), .B2(G45), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n705), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(new_n689), .B2(G330), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n231), .B1(G20), .B2(new_n330), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n328), .A2(new_n564), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n204), .A2(G190), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G317), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT33), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n754), .A2(KEYINPUT33), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n753), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G179), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n751), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G329), .ZN(new_n761));
  INV_X1    g0561(.A(G283), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n564), .A2(G179), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n751), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n757), .B(new_n761), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n204), .B1(new_n758), .B2(G190), .ZN(new_n766));
  INV_X1    g0566(.A(G294), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G311), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n328), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n751), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n769), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n204), .A2(new_n349), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n750), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n301), .B(new_n773), .C1(G326), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n774), .A2(new_n763), .ZN(new_n778));
  INV_X1    g0578(.A(G322), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n774), .A2(new_n771), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n777), .B1(new_n547), .B2(new_n778), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n778), .A2(new_n213), .ZN(new_n782));
  INV_X1    g0582(.A(new_n764), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n366), .B(new_n782), .C1(G107), .C2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT93), .ZN(new_n785));
  INV_X1    g0585(.A(new_n766), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n785), .B1(G97), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n780), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G58), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n752), .A2(new_n210), .B1(new_n772), .B2(new_n223), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(G50), .B2(new_n776), .ZN(new_n791));
  INV_X1    g0591(.A(G159), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n759), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT32), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n787), .A2(new_n789), .A3(new_n791), .A4(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n749), .B1(new_n781), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n703), .A2(new_n301), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(new_n507), .B2(new_n235), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n247), .B2(new_n507), .ZN(new_n800));
  INV_X1    g0600(.A(G355), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n207), .A2(new_n301), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n800), .B1(G116), .B2(new_n207), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(G13), .A2(G33), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(G20), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n748), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n746), .ZN(new_n809));
  INV_X1    g0609(.A(new_n806), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n808), .B(new_n809), .C1(new_n689), .C2(new_n810), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n744), .A2(new_n747), .B1(new_n796), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT94), .ZN(G396));
  NAND2_X1  g0613(.A1(new_n355), .A2(KEYINPUT95), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT95), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n353), .A2(new_n348), .A3(new_n815), .A4(new_n354), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n351), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n735), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n355), .A2(new_n692), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n348), .A2(new_n684), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n734), .B(new_n818), .C1(new_n735), .C2(new_n822), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n823), .A2(KEYINPUT96), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n809), .B1(new_n823), .B2(KEYINPUT96), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n818), .B1(new_n735), .B2(new_n822), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n733), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT97), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n826), .A2(KEYINPUT97), .A3(new_n733), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n824), .A2(new_n825), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n772), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G143), .A2(new_n788), .B1(new_n832), .B2(G159), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n834), .B2(new_n775), .C1(new_n261), .C2(new_n752), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT34), .Z(new_n836));
  INV_X1    g0636(.A(new_n778), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n836), .B1(G50), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n366), .B1(new_n760), .B2(G132), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n786), .A2(G58), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n783), .A2(G68), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G311), .A2(new_n760), .B1(new_n786), .B2(G97), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n470), .B2(new_n778), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n366), .B1(new_n780), .B2(new_n767), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n213), .A2(new_n764), .B1(new_n772), .B2(new_n535), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n847), .B1(new_n762), .B2(new_n752), .C1(new_n547), .C2(new_n775), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n749), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n748), .A2(new_n804), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n746), .B(new_n849), .C1(new_n223), .C2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n805), .B2(new_n822), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n831), .A2(new_n852), .ZN(G384));
  NOR2_X1   g0653(.A1(new_n450), .A2(new_n684), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n404), .A2(new_n405), .ZN(new_n856));
  INV_X1    g0656(.A(new_n682), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n405), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n397), .A2(new_n398), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n855), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n860), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n405), .B1(new_n404), .B2(new_n857), .ZN(new_n863));
  XOR2_X1   g0663(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n409), .B2(new_n858), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(KEYINPUT38), .B(new_n867), .C1(new_n409), .C2(new_n858), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n864), .B1(new_n859), .B2(KEYINPUT101), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n862), .A2(new_n863), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n862), .A2(KEYINPUT101), .A3(new_n863), .A4(new_n864), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n669), .A2(new_n670), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n858), .B1(new_n674), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n869), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT39), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n871), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n872), .A2(KEYINPUT39), .B1(new_n882), .B2(KEYINPUT100), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n671), .A2(new_n674), .A3(new_n672), .ZN(new_n884));
  INV_X1    g0684(.A(new_n858), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n886), .B2(new_n867), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n869), .B(new_n866), .C1(new_n884), .C2(new_n885), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT100), .B(KEYINPUT39), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n854), .B1(new_n883), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n408), .A2(new_n682), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n814), .A2(new_n692), .A3(new_n816), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n735), .B2(new_n817), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n449), .A2(new_n684), .ZN(new_n897));
  NOR3_X1   g0697(.A1(new_n432), .A2(new_n434), .A3(new_n436), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n452), .B(new_n897), .C1(new_n898), .C2(new_n448), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n438), .A2(new_n449), .A3(new_n684), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n896), .A2(new_n901), .A3(new_n872), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n891), .A2(new_n892), .A3(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n736), .A2(new_n410), .A3(new_n456), .A4(new_n741), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n904), .A2(new_n676), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n903), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n871), .A2(new_n880), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n821), .B1(new_n899), .B2(new_n900), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n732), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT40), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(KEYINPUT102), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT102), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n909), .A2(new_n732), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n912), .A2(new_n872), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n457), .A2(new_n732), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n917), .B(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(G330), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n906), .B(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n203), .B2(new_n678), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT35), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n619), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(G116), .A3(new_n233), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT98), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n923), .B2(new_n619), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT36), .ZN(new_n928));
  OAI21_X1  g0728(.A(G77), .B1(new_n226), .B2(new_n210), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n929), .A2(new_n234), .B1(G50), .B2(new_n210), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(G1), .A3(new_n256), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n922), .A2(new_n928), .A3(new_n931), .ZN(G367));
  OR2_X1    g0732(.A1(new_n651), .A2(new_n692), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n933), .A2(new_n646), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n933), .A2(new_n646), .A3(new_n653), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n656), .B1(new_n625), .B2(new_n684), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n700), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n940), .B(new_n941), .Z(new_n942));
  AOI21_X1  g0742(.A(new_n659), .B1(new_n938), .B2(new_n695), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(new_n684), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n937), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n945), .B(new_n946), .Z(new_n947));
  OAI21_X1  g0747(.A(new_n939), .B1(new_n626), .B2(new_n692), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n691), .A2(new_n697), .A3(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n947), .B(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n704), .B(KEYINPUT41), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT104), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n698), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(KEYINPUT105), .B1(new_n697), .B2(new_n699), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(new_n700), .ZN(new_n956));
  MUX2_X1   g0756(.A(new_n690), .B(new_n744), .S(new_n956), .Z(new_n957));
  AND2_X1   g0757(.A1(new_n957), .A2(new_n742), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n701), .A2(new_n948), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT45), .Z(new_n960));
  NOR2_X1   g0760(.A1(new_n701), .A2(new_n948), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT44), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(new_n698), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n954), .B(new_n958), .C1(new_n964), .C2(new_n953), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n952), .B1(new_n965), .B2(new_n742), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n745), .B(KEYINPUT106), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n950), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n807), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n239), .A2(new_n798), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n969), .B(new_n970), .C1(new_n703), .C2(new_n343), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n366), .B1(new_n766), .B2(new_n470), .C1(new_n547), .C2(new_n780), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n783), .A2(G97), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n754), .B2(new_n759), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n972), .B(new_n974), .C1(G283), .C2(new_n832), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n837), .A2(G116), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT46), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n975), .B(new_n977), .C1(new_n767), .C2(new_n752), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n775), .A2(new_n770), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n301), .B1(new_n752), .B2(new_n792), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(G50), .B2(new_n832), .ZN(new_n981));
  AOI22_X1  g0781(.A1(G77), .A2(new_n783), .B1(new_n760), .B2(G137), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(new_n226), .C2(new_n778), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n776), .A2(G143), .B1(new_n786), .B2(G68), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n261), .B2(new_n780), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT107), .Z(new_n986));
  OAI22_X1  g0786(.A1(new_n978), .A2(new_n979), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n971), .B1(new_n988), .B2(new_n748), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n989), .B(new_n809), .C1(new_n810), .C2(new_n936), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n968), .A2(new_n990), .ZN(G387));
  NAND2_X1  g0791(.A1(new_n957), .A2(new_n967), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n697), .A2(new_n810), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G322), .A2(new_n776), .B1(new_n753), .B2(G311), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n547), .B2(new_n772), .C1(new_n754), .C2(new_n780), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT48), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n762), .B2(new_n766), .C1(new_n767), .C2(new_n778), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT49), .Z(new_n998));
  AOI21_X1  g0798(.A(new_n301), .B1(new_n760), .B2(G326), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n535), .B2(new_n764), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n344), .A2(new_n766), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n776), .A2(G159), .B1(new_n760), .B2(G150), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n221), .B2(new_n780), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1002), .B(new_n1004), .C1(G77), .C2(new_n837), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n268), .A2(new_n753), .B1(new_n832), .B2(G68), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT109), .Z(new_n1007));
  AND4_X1   g0807(.A1(new_n301), .A2(new_n1005), .A3(new_n973), .A4(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n748), .B1(new_n1001), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n346), .A2(new_n221), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT108), .Z(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g0812(.A(G45), .B1(new_n1011), .B2(KEYINPUT50), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(G68), .A2(G77), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n707), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n797), .B1(new_n243), .B2(new_n507), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n707), .B2(new_n802), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n1015), .A2(new_n1017), .B1(new_n470), .B2(new_n703), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1009), .B(new_n809), .C1(new_n969), .C2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n704), .B1(new_n957), .B2(new_n742), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n992), .B1(new_n993), .B2(new_n1019), .C1(new_n958), .C2(new_n1020), .ZN(G393));
  OR2_X1    g0821(.A1(new_n964), .A2(new_n958), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n965), .A2(new_n1022), .A3(new_n704), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n948), .A2(new_n810), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n807), .B1(new_n798), .B2(new_n250), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G97), .B2(new_n703), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n775), .A2(new_n754), .B1(new_n780), .B2(new_n770), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT52), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n764), .A2(new_n470), .B1(new_n759), .B2(new_n779), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n772), .A2(new_n767), .B1(new_n766), .B2(new_n535), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n366), .B1(new_n752), .B2(new_n547), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1028), .B(new_n1032), .C1(new_n762), .C2(new_n778), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n346), .A2(new_n832), .B1(G50), .B2(new_n753), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT110), .Z(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G68), .B2(new_n837), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n766), .A2(new_n223), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G87), .B2(new_n783), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n366), .B1(new_n760), .B2(G143), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1036), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n775), .A2(new_n261), .B1(new_n780), .B2(new_n792), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT51), .Z(new_n1042));
  OAI21_X1  g0842(.A(new_n1033), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n746), .B(new_n1026), .C1(new_n1043), .C2(new_n748), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n964), .A2(new_n967), .B1(new_n1024), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1023), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(KEYINPUT111), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT111), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1023), .A2(new_n1048), .A3(new_n1045), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(G390));
  NAND2_X1  g0850(.A1(new_n882), .A2(KEYINPUT100), .ZN(new_n1051));
  OAI21_X1  g0851(.A(KEYINPUT39), .B1(new_n887), .B2(new_n888), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n854), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n901), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1054), .B1(new_n895), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1053), .A2(new_n1056), .A3(new_n889), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n692), .B1(new_n737), .B2(new_n740), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n817), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n893), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n907), .B(new_n1054), .C1(new_n1061), .C2(new_n1055), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1057), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n732), .A2(new_n901), .A3(G330), .A4(new_n822), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1057), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n967), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1053), .A2(new_n804), .A3(new_n889), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n841), .B1(new_n535), .B2(new_n780), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1037), .B(new_n1071), .C1(G283), .C2(new_n776), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n366), .B1(new_n759), .B2(new_n767), .C1(new_n470), .C2(new_n752), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n782), .B(new_n1073), .C1(G97), .C2(new_n832), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n366), .B1(new_n783), .B2(G50), .ZN(new_n1076));
  INV_X1    g0876(.A(G125), .ZN(new_n1077));
  INV_X1    g0877(.A(G128), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1076), .B1(new_n1077), .B2(new_n759), .C1(new_n1078), .C2(new_n775), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G137), .B2(new_n753), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT54), .B(G143), .Z(new_n1081));
  AOI22_X1  g0881(.A1(G132), .A2(new_n788), .B1(new_n832), .B2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1080), .B(new_n1082), .C1(new_n792), .C2(new_n766), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n778), .A2(new_n261), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1075), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT116), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n746), .B1(new_n1088), .B2(new_n748), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n850), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1070), .B(new_n1089), .C1(new_n268), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1069), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT114), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n410), .A2(G330), .A3(new_n456), .A4(new_n732), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n904), .A2(new_n1094), .A3(new_n676), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n730), .A2(new_n731), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n566), .A2(new_n635), .A3(new_n684), .ZN(new_n1098));
  OAI211_X1 g0898(.A(G330), .B(new_n822), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n1055), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1065), .B1(KEYINPUT112), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT112), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1099), .A2(new_n1102), .A3(new_n1055), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n895), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT113), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n821), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1099), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1100), .A2(new_n1064), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1060), .B(new_n1108), .C1(new_n1109), .C2(new_n1107), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1093), .B(new_n1096), .C1(new_n1104), .C2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1100), .A2(KEYINPUT112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1113), .A2(new_n1064), .A3(new_n1103), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n896), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1109), .A2(new_n1107), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1108), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n1061), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1093), .B1(new_n1119), .B2(new_n1096), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1112), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1060), .B1(new_n1109), .B2(new_n1107), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1117), .A2(new_n1124), .B1(new_n1114), .B2(new_n896), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT114), .B1(new_n1125), .B2(new_n1095), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n1111), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n705), .B1(new_n1127), .B2(new_n1068), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1092), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(G378));
  INV_X1    g0930(.A(KEYINPUT55), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n326), .B2(new_n332), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n326), .A2(new_n1131), .A3(new_n332), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n289), .A2(new_n682), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(KEYINPUT55), .B(new_n333), .C1(new_n318), .C2(new_n325), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1135), .B1(new_n1132), .B2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n909), .A2(new_n732), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n913), .B1(new_n1145), .B2(new_n907), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1145), .A2(new_n914), .B1(new_n871), .B2(new_n870), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n912), .ZN(new_n1148));
  INV_X1    g0948(.A(G330), .ZN(new_n1149));
  OAI211_X1 g0949(.A(KEYINPUT119), .B(new_n1144), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT118), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1140), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1136), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n1132), .A2(new_n1138), .A3(new_n1135), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(KEYINPUT118), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT119), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(KEYINPUT118), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1152), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(G330), .A3(new_n917), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1150), .A2(new_n903), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n903), .B1(new_n1150), .B2(new_n1162), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1122), .B1(new_n1126), .B2(new_n1111), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n1095), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT57), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n705), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1165), .B(KEYINPUT57), .C1(new_n1166), .C2(new_n1095), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(KEYINPUT120), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1068), .B1(new_n1112), .B2(new_n1120), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n1096), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT120), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1173), .A2(new_n1174), .A3(KEYINPUT57), .A4(new_n1165), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1169), .A2(new_n1171), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n903), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1159), .B(new_n1143), .C1(new_n917), .C2(G330), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1161), .A2(G330), .A3(new_n917), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1150), .A2(new_n903), .A3(new_n1162), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n967), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1152), .A2(new_n804), .A3(new_n1158), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n746), .B1(new_n221), .B2(new_n850), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G128), .A2(new_n788), .B1(new_n832), .B2(G137), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n837), .A2(new_n1081), .B1(new_n786), .B2(G150), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(new_n1077), .C2(new_n775), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G132), .B2(new_n753), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT59), .ZN(new_n1189));
  AOI21_X1  g0989(.A(G33), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(G41), .B1(new_n760), .B2(G124), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G159), .B2(new_n783), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n1189), .B2(new_n1188), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n223), .A2(new_n778), .B1(new_n780), .B2(new_n470), .ZN(new_n1195));
  AOI211_X1 g0995(.A(G41), .B(new_n1195), .C1(G68), .C2(new_n786), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n301), .B1(new_n783), .B2(G58), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n832), .A2(new_n343), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n753), .A2(G97), .B1(new_n760), .B2(G283), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G116), .B2(new_n776), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT58), .Z(new_n1202));
  OAI21_X1  g1002(.A(new_n221), .B1(new_n364), .B2(G41), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1194), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1183), .B(new_n1184), .C1(new_n749), .C2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1182), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1176), .A2(new_n1207), .ZN(G375));
  NAND3_X1  g1008(.A1(new_n1115), .A2(new_n1118), .A3(new_n1095), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(KEYINPUT121), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT121), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1125), .A2(new_n1211), .A3(new_n1095), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1121), .A2(new_n951), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1119), .A2(new_n967), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1055), .A2(new_n804), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT122), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1002), .B1(G283), .B2(new_n788), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT123), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n772), .A2(new_n470), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n366), .B1(new_n752), .B2(new_n535), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n778), .A2(new_n215), .B1(new_n764), .B2(new_n223), .ZN(new_n1222));
  NOR4_X1   g1022(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(new_n767), .B2(new_n775), .C1(new_n547), .C2(new_n759), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n301), .B1(new_n780), .B2(new_n834), .C1(new_n792), .C2(new_n778), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n753), .A2(new_n1081), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n766), .A2(new_n221), .ZN(new_n1227));
  INV_X1    g1027(.A(G132), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n775), .A2(new_n1228), .B1(new_n764), .B2(new_n226), .ZN(new_n1229));
  NOR4_X1   g1029(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1229), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1230), .B1(new_n1078), .B2(new_n759), .C1(new_n261), .C2(new_n772), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n749), .B1(new_n1224), .B2(new_n1231), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n746), .B(new_n1232), .C1(new_n210), .C2(new_n850), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1217), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1215), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1214), .A2(new_n1236), .ZN(G381));
  NAND4_X1  g1037(.A1(new_n1047), .A2(new_n968), .A3(new_n990), .A4(new_n1049), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1176), .A2(new_n1129), .A3(new_n1207), .ZN(new_n1239));
  OR2_X1    g1039(.A1(G393), .A2(G396), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(G384), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1241), .A2(new_n1242), .A3(new_n1236), .A4(new_n1214), .ZN(G407));
  OAI211_X1 g1043(.A(G407), .B(G213), .C1(G343), .C2(new_n1239), .ZN(G409));
  NAND2_X1  g1044(.A1(G375), .A2(G378), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1182), .A2(KEYINPUT124), .A3(new_n1205), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT124), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1206), .A2(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1165), .B(new_n951), .C1(new_n1166), .C2(new_n1095), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1129), .A2(new_n1246), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n683), .A2(G213), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1125), .A2(KEYINPUT60), .A3(new_n1095), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1126), .A2(KEYINPUT60), .A3(new_n1111), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1256), .B1(new_n1257), .B2(new_n1213), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1242), .B(new_n1235), .C1(new_n1258), .C2(new_n704), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1213), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n704), .A3(new_n1255), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G384), .B1(new_n1261), .B2(new_n1236), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1254), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n705), .B(new_n1256), .C1(new_n1257), .C2(new_n1213), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1242), .B1(new_n1264), .B2(new_n1235), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1261), .A2(G384), .A3(new_n1236), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(KEYINPUT125), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n683), .A2(G213), .A3(G2897), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n1245), .A2(new_n1253), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1269), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT61), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G390), .A2(G387), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1238), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1240), .A2(KEYINPUT126), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1277), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1240), .A2(new_n1276), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(KEYINPUT126), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1274), .B(new_n1238), .C1(new_n1279), .C2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1252), .B1(G375), .B2(G378), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1284), .A2(KEYINPUT63), .A3(new_n1268), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1245), .A2(new_n1268), .A3(new_n1253), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1273), .A2(new_n1283), .A3(new_n1285), .A4(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1245), .A2(new_n1253), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1267), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT125), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1269), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1290), .A2(new_n1293), .A3(new_n1272), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT62), .ZN(new_n1298));
  AOI211_X1 g1098(.A(new_n1297), .B(new_n1298), .C1(new_n1284), .C2(new_n1268), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT62), .B1(new_n1286), .B2(KEYINPUT127), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1296), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1289), .B1(new_n1301), .B2(new_n1283), .ZN(G405));
  AND2_X1   g1102(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1245), .A2(new_n1239), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1304), .B1(new_n1262), .B2(new_n1259), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1245), .A2(new_n1268), .A3(new_n1239), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1303), .B(new_n1307), .ZN(G402));
endmodule


