//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n441, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n571, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n605, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1135, new_n1136;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  XOR2_X1   g007(.A(KEYINPUT66), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT67), .ZN(G220));
  XOR2_X1   g012(.A(KEYINPUT68), .B(G96), .Z(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT69), .B(G57), .ZN(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(new_n441), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT70), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT72), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(G2104), .ZN(new_n464));
  NOR3_X1   g039(.A1(new_n460), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n461), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT71), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n461), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n470), .B1(new_n461), .B2(new_n469), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n468), .B1(new_n475), .B2(G2105), .ZN(G160));
  NOR2_X1   g051(.A1(new_n463), .A2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT72), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n462), .A2(new_n463), .A3(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  OR3_X1    g058(.A1(new_n482), .A2(KEYINPUT73), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n485), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT73), .B1(new_n482), .B2(new_n483), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n484), .A2(new_n488), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NOR2_X1   g068(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT71), .B1(new_n477), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n461), .A2(new_n469), .A3(new_n470), .ZN(new_n496));
  AOI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(KEYINPUT4), .B1(new_n497), .B2(G138), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n478), .A2(new_n479), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n499), .A2(G126), .A3(G2105), .A4(new_n461), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT4), .A2(G138), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n499), .A2(new_n485), .A3(new_n461), .A4(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(new_n485), .B2(G114), .ZN(new_n503));
  NOR2_X1   g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT74), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OR2_X1    g080(.A1(G102), .A2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(G114), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G2105), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n506), .A2(new_n508), .A3(new_n509), .A4(G2104), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n500), .A2(new_n502), .A3(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n498), .A2(new_n512), .ZN(G164));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(new_n514), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  OAI221_X1 g101(.A(new_n517), .B1(new_n518), .B2(new_n524), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(G166));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT76), .ZN(new_n533));
  XOR2_X1   g108(.A(new_n533), .B(KEYINPUT7), .Z(new_n534));
  AOI22_X1  g109(.A1(new_n514), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n520), .A2(new_n522), .ZN(new_n536));
  INV_X1    g111(.A(G51), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n535), .A2(new_n536), .B1(new_n537), .B2(new_n515), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n534), .A2(new_n538), .ZN(G168));
  AOI22_X1  g114(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n525), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(KEYINPUT77), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n524), .A2(new_n543), .B1(new_n515), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n541), .A2(KEYINPUT77), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n542), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n525), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n524), .A2(new_n552), .B1(new_n515), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT78), .Z(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n516), .A2(G53), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(new_n524), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  XOR2_X1   g141(.A(KEYINPUT79), .B(G65), .Z(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n567), .B2(new_n536), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n565), .A2(G91), .B1(new_n568), .B2(G651), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n564), .A2(new_n569), .ZN(G299));
  XOR2_X1   g145(.A(new_n548), .B(KEYINPUT80), .Z(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  INV_X1    g148(.A(G166), .ZN(G303));
  NAND2_X1  g149(.A1(new_n565), .A2(G87), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n516), .A2(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  AOI22_X1  g153(.A1(new_n523), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n525), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  INV_X1    g156(.A(G48), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n524), .A2(new_n581), .B1(new_n515), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n516), .A2(G47), .ZN(new_n586));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI221_X1 g163(.A(new_n586), .B1(new_n587), .B2(new_n524), .C1(new_n525), .C2(new_n588), .ZN(G290));
  INV_X1    g164(.A(G92), .ZN(new_n590));
  OR3_X1    g165(.A1(new_n524), .A2(KEYINPUT10), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n536), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n516), .A2(G54), .B1(new_n594), .B2(G651), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT10), .B1(new_n524), .B2(new_n590), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n571), .B2(new_n598), .ZN(G284));
  OAI21_X1  g175(.A(new_n599), .B1(new_n571), .B2(new_n598), .ZN(G321));
  NAND2_X1  g176(.A1(G299), .A2(new_n598), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n598), .B2(G168), .ZN(G297));
  OAI21_X1  g178(.A(new_n602), .B1(new_n598), .B2(G168), .ZN(G280));
  INV_X1    g179(.A(new_n597), .ZN(new_n605));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI211_X1 g186(.A(G2104), .B(new_n485), .C1(new_n471), .C2(new_n472), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT13), .Z(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(G2100), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n487), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n481), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n485), .A2(G111), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT81), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n616), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND2_X1  g197(.A1(new_n614), .A2(G2100), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n615), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT82), .ZN(G156));
  XOR2_X1   g200(.A(G2427), .B(G2430), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT83), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2438), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT84), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n629), .B2(new_n627), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT85), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2443), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2446), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n636), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G14), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT86), .ZN(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n644), .B1(new_n648), .B2(KEYINPUT18), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n648), .A2(KEYINPUT17), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n646), .A2(new_n647), .ZN(new_n653));
  AOI21_X1  g228(.A(KEYINPUT18), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n651), .B(new_n654), .Z(G227));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  AOI21_X1  g235(.A(KEYINPUT87), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AND3_X1   g236(.A1(new_n659), .A2(new_n660), .A3(KEYINPUT87), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n659), .A2(new_n660), .ZN(new_n665));
  AOI22_X1  g240(.A1(new_n663), .A2(new_n664), .B1(new_n658), .B2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n665), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n659), .A2(new_n660), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(new_n657), .A3(new_n668), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n666), .B(new_n669), .C1(new_n664), .C2(new_n663), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT88), .B(G1981), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(G229));
  AND2_X1   g252(.A1(KEYINPUT90), .A2(G16), .ZN(new_n678));
  NOR2_X1   g253(.A1(KEYINPUT90), .A2(G16), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n680), .A2(G22), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(G166), .B2(new_n680), .ZN(new_n682));
  INV_X1    g257(.A(G1971), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(G16), .A2(G23), .ZN(new_n685));
  INV_X1    g260(.A(G288), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(G16), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT33), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G6), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n584), .B2(new_n690), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT92), .B(G1981), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT32), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n684), .A2(new_n689), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT93), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(KEYINPUT34), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(KEYINPUT34), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G25), .A2(G29), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n487), .A2(G131), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n481), .A2(G119), .ZN(new_n703));
  OR2_X1    g278(.A1(G95), .A2(G2105), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n704), .B(G2104), .C1(G107), .C2(new_n485), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n701), .B1(new_n707), .B2(G29), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT89), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT35), .B(G1991), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G24), .B(G290), .S(new_n680), .Z(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT91), .B(G1986), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  OR3_X1    g290(.A1(new_n700), .A2(KEYINPUT36), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(KEYINPUT36), .B1(new_n700), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n680), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n719), .A2(KEYINPUT23), .A3(G20), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT23), .ZN(new_n721));
  INV_X1    g296(.A(G20), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n680), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G299), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n720), .B(new_n723), .C1(new_n724), .C2(new_n690), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(G1956), .Z(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G26), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n487), .A2(G140), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n481), .A2(G128), .ZN(new_n730));
  OR2_X1    g305(.A1(G104), .A2(G2105), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n731), .B(G2104), .C1(G116), .C2(new_n485), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n728), .B1(new_n734), .B2(new_n727), .ZN(new_n735));
  MUX2_X1   g310(.A(new_n728), .B(new_n735), .S(KEYINPUT28), .Z(new_n736));
  INV_X1    g311(.A(KEYINPUT99), .ZN(new_n737));
  AND3_X1   g312(.A1(new_n500), .A2(new_n502), .A3(new_n511), .ZN(new_n738));
  OAI211_X1 g313(.A(G138), .B(new_n485), .C1(new_n471), .C2(new_n472), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT4), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G29), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n727), .A2(G27), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n737), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n737), .B2(new_n744), .ZN(new_n746));
  INV_X1    g321(.A(G2078), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n736), .A2(G2067), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(G171), .A2(G16), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G5), .B2(G16), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n726), .B(new_n748), .C1(G1961), .C2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G4), .A2(G16), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n605), .B2(G16), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G1348), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G28), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(G28), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n758), .A2(new_n759), .A3(new_n727), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n755), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n621), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n761), .B1(G29), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G1966), .ZN(new_n764));
  NAND2_X1  g339(.A1(G168), .A2(G16), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G16), .B2(G21), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n763), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n766), .A2(new_n764), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(KEYINPUT97), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT24), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(G34), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(G34), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G125), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n495), .B2(new_n496), .ZN(new_n775));
  INV_X1    g350(.A(new_n474), .ZN(new_n776));
  OAI21_X1  g351(.A(G2105), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n468), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n773), .B1(new_n779), .B2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G2084), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n768), .A2(KEYINPUT97), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n769), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n752), .A2(new_n767), .A3(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n736), .A2(G2067), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n719), .A2(G19), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n555), .B2(new_n719), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(G1341), .Z(new_n788));
  AND3_X1   g363(.A1(new_n784), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G29), .A2(G32), .ZN(new_n790));
  AOI22_X1  g365(.A1(G141), .A2(new_n487), .B1(new_n481), .B2(G129), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n485), .A2(G105), .A3(G2104), .ZN(new_n792));
  NAND3_X1  g367(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT95), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT26), .ZN(new_n795));
  AND3_X1   g370(.A1(new_n791), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT96), .Z(new_n797));
  AOI21_X1  g372(.A(new_n790), .B1(new_n797), .B2(G29), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT27), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G1996), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G1348), .B2(new_n754), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n746), .A2(new_n747), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n799), .A2(G1996), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n718), .A2(new_n789), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n751), .A2(G1961), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT98), .ZN(new_n807));
  OAI21_X1  g382(.A(G127), .B1(new_n471), .B2(new_n472), .ZN(new_n808));
  INV_X1    g383(.A(G115), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n460), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G2105), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT94), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n487), .A2(G139), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n485), .A2(G103), .A3(G2104), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT25), .Z(new_n815));
  NAND3_X1  g390(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  MUX2_X1   g391(.A(G33), .B(new_n816), .S(G29), .Z(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(G2072), .Z(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G29), .A2(G35), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G162), .B2(G29), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT29), .ZN(new_n822));
  INV_X1    g397(.A(G2090), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n805), .A2(new_n807), .A3(new_n819), .A4(new_n825), .ZN(G311));
  NOR2_X1   g401(.A1(new_n805), .A2(new_n825), .ZN(new_n827));
  INV_X1    g402(.A(new_n807), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n827), .A2(new_n828), .A3(new_n818), .ZN(G150));
  NAND2_X1  g404(.A1(new_n516), .A2(G55), .ZN(new_n830));
  INV_X1    g405(.A(G93), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  OAI221_X1 g407(.A(new_n830), .B1(new_n831), .B2(new_n524), .C1(new_n525), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G860), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n605), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT39), .Z(new_n839));
  INV_X1    g414(.A(KEYINPUT100), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n555), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT101), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n833), .B1(new_n555), .B2(new_n840), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n839), .B(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n836), .B1(new_n847), .B2(G860), .ZN(G145));
  XNOR2_X1  g423(.A(new_n706), .B(KEYINPUT103), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n849), .A2(new_n613), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n613), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n487), .A2(G142), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n481), .A2(G130), .ZN(new_n854));
  OR2_X1    g429(.A1(G106), .A2(G2105), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(G2104), .C1(G118), .C2(new_n485), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n850), .A2(new_n851), .A3(new_n857), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n797), .A2(new_n816), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n816), .A2(new_n796), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n859), .A2(new_n862), .A3(new_n863), .A4(new_n860), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n733), .B(new_n742), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n865), .A2(new_n868), .A3(new_n866), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n762), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n870), .A2(new_n871), .A3(new_n872), .A4(new_n621), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n492), .B(new_n779), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n874), .A2(new_n877), .A3(new_n875), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g458(.A1(new_n833), .A2(new_n598), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n846), .B(new_n608), .Z(new_n885));
  XNOR2_X1  g460(.A(G299), .B(new_n605), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n887), .A2(KEYINPUT41), .ZN(new_n888));
  XOR2_X1   g463(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n886), .B2(new_n885), .ZN(new_n892));
  XNOR2_X1  g467(.A(G166), .B(G305), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n686), .B(G290), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n892), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n884), .B1(new_n898), .B2(new_n598), .ZN(G295));
  OAI21_X1  g474(.A(new_n884), .B1(new_n898), .B2(new_n598), .ZN(G331));
  NOR2_X1   g475(.A1(new_n548), .A2(G168), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n571), .B2(G286), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT107), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT107), .B1(new_n844), .B2(new_n845), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n907), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n905), .A3(new_n903), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n910), .A3(new_n886), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n890), .B1(new_n908), .B2(new_n910), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n895), .ZN(new_n915));
  INV_X1    g490(.A(new_n895), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n912), .B2(new_n913), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n880), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n920));
  AOI21_X1  g495(.A(G37), .B1(new_n914), .B2(new_n895), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n886), .A2(new_n889), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n886), .A2(KEYINPUT41), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n906), .A2(new_n904), .A3(new_n907), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n903), .B1(new_n909), .B2(new_n905), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n922), .B(new_n923), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n911), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT108), .B1(new_n927), .B2(new_n916), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n929));
  AOI211_X1 g504(.A(new_n929), .B(new_n895), .C1(new_n926), .C2(new_n911), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n920), .B(new_n921), .C1(new_n928), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n919), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n918), .A2(new_n920), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n921), .B1(new_n928), .B2(new_n930), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n933), .B1(new_n934), .B2(new_n920), .ZN(new_n935));
  MUX2_X1   g510(.A(new_n932), .B(new_n935), .S(KEYINPUT44), .Z(G397));
  INV_X1    g511(.A(G1384), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(new_n498), .B2(new_n512), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(G160), .B2(G40), .ZN(new_n941));
  AND4_X1   g516(.A1(new_n940), .A2(new_n777), .A3(new_n778), .A4(G40), .ZN(new_n942));
  NOR4_X1   g517(.A1(new_n939), .A2(new_n941), .A3(new_n942), .A4(KEYINPUT45), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n943), .A2(KEYINPUT110), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(KEYINPUT110), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G2067), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n733), .B(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G1996), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n797), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(new_n950), .B2(new_n796), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n946), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n953), .A2(KEYINPUT112), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(KEYINPUT112), .ZN(new_n955));
  INV_X1    g530(.A(new_n946), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n706), .B(new_n710), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n954), .B(new_n955), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(G290), .A2(G1986), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(KEYINPUT111), .ZN(new_n960));
  NAND2_X1  g535(.A1(G290), .A2(G1986), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n960), .B(new_n961), .Z(new_n962));
  AOI21_X1  g537(.A(new_n958), .B1(new_n946), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT61), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT57), .ZN(new_n965));
  INV_X1    g540(.A(new_n569), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n965), .B1(new_n966), .B2(KEYINPUT118), .ZN(new_n967));
  XNOR2_X1  g542(.A(G299), .B(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G40), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT109), .B1(new_n779), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(G160), .A2(new_n940), .A3(G40), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT50), .B1(new_n742), .B2(new_n937), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n974), .B(G1384), .C1(new_n738), .C2(new_n741), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n971), .B(new_n972), .C1(new_n973), .C2(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(KEYINPUT116), .B(G1956), .Z(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT117), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT117), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n976), .A2(new_n981), .A3(new_n978), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n938), .B(KEYINPUT45), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n941), .A2(new_n942), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT56), .B(G2072), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n969), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n938), .A2(new_n974), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n742), .A2(KEYINPUT50), .A3(new_n937), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI211_X1 g566(.A(KEYINPUT117), .B(new_n977), .C1(new_n985), .C2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n981), .B1(new_n976), .B2(new_n978), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n969), .B(new_n987), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n964), .B1(new_n988), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n971), .A2(new_n939), .A3(new_n972), .ZN(new_n997));
  XOR2_X1   g572(.A(KEYINPUT58), .B(G1341), .Z(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n984), .A2(new_n985), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n999), .B1(new_n1000), .B2(G1996), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n555), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT59), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n996), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n994), .A2(KEYINPUT61), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n987), .B1(new_n992), .B2(new_n993), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n968), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT120), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1006), .A2(new_n1009), .A3(new_n968), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1005), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT121), .B1(new_n1004), .B2(new_n1011), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1006), .A2(new_n1009), .A3(new_n968), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1009), .B1(new_n1006), .B2(new_n968), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT61), .B(new_n994), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT121), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(new_n996), .A4(new_n1003), .ZN(new_n1017));
  INV_X1    g592(.A(new_n976), .ZN(new_n1018));
  OAI22_X1  g593(.A1(new_n1018), .A2(G1348), .B1(G2067), .B2(new_n997), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT119), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n1021));
  OAI221_X1 g596(.A(new_n1021), .B1(G2067), .B2(new_n997), .C1(new_n1018), .C2(G1348), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1023), .A2(KEYINPUT60), .A3(new_n597), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n597), .B1(new_n1023), .B2(KEYINPUT60), .ZN(new_n1025));
  OAI22_X1  g600(.A1(new_n1024), .A2(new_n1025), .B1(KEYINPUT60), .B2(new_n1023), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1012), .A2(new_n1017), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT122), .ZN(new_n1028));
  OAI22_X1  g603(.A1(new_n1013), .A2(new_n1014), .B1(new_n597), .B2(new_n1023), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n994), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1028), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n984), .A2(new_n985), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n747), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1018), .A2(G1961), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1035), .A2(KEYINPUT123), .ZN(new_n1040));
  OR3_X1    g615(.A1(new_n1000), .A2(KEYINPUT123), .A3(G2078), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(KEYINPUT53), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(G301), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n779), .A2(new_n970), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n984), .A2(KEYINPUT53), .A3(new_n747), .A4(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1037), .A2(new_n1038), .A3(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(new_n571), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1033), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n1048), .A2(KEYINPUT124), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1034), .A2(G1971), .B1(G2090), .B2(new_n976), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1050), .A2(KEYINPUT113), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G303), .A2(G8), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1052), .B(KEYINPUT55), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1050), .A2(KEYINPUT113), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1051), .A2(new_n1054), .A3(G8), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G305), .A2(G1981), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(KEYINPUT49), .ZN(new_n1058));
  OR2_X1    g633(.A1(G305), .A2(G1981), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT115), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  OR2_X1    g636(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n997), .A2(G8), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1976), .ZN(new_n1066));
  NOR2_X1   g641(.A1(G288), .A2(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1067), .A2(KEYINPUT114), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(KEYINPUT114), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1063), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT52), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1065), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n686), .A2(G1976), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1070), .A2(KEYINPUT52), .A3(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1050), .A2(G8), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1053), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1056), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1033), .B1(new_n1079), .B2(G301), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1046), .A2(G171), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1034), .A2(G1966), .B1(G2084), .B2(new_n976), .ZN(new_n1083));
  OAI21_X1  g658(.A(G8), .B1(new_n1083), .B2(G286), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT51), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1086), .B1(new_n1083), .B2(G286), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1048), .A2(KEYINPUT124), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1049), .A2(new_n1082), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1031), .A2(new_n1032), .A3(new_n1090), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1056), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1063), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1065), .A2(new_n1066), .A3(new_n686), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(new_n1059), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1056), .A2(new_n1075), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1083), .A2(G8), .A3(G168), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT63), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1051), .A2(G8), .A3(new_n1055), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1099), .B2(new_n1053), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n1092), .B(new_n1095), .C1(new_n1101), .C2(KEYINPUT63), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1088), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT125), .B1(new_n1088), .B2(KEYINPUT62), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1088), .A2(KEYINPUT62), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1106), .A2(G301), .A3(new_n1079), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1105), .A2(new_n1107), .B1(new_n1097), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1102), .B1(new_n1109), .B2(new_n1078), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n963), .B1(new_n1091), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n956), .B1(new_n796), .B2(new_n948), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n946), .A2(KEYINPUT46), .A3(new_n950), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT46), .B1(new_n946), .B2(new_n950), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT47), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n954), .A2(new_n955), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n707), .A2(new_n710), .ZN(new_n1118));
  OAI22_X1  g693(.A1(new_n1117), .A2(new_n1118), .B1(G2067), .B2(new_n733), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1119), .A2(new_n946), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n946), .A2(new_n959), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT48), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n958), .B(new_n1123), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1116), .B(new_n1120), .C1(new_n1122), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1111), .A2(new_n1125), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g701(.A(G401), .ZN(new_n1128));
  INV_X1    g702(.A(G229), .ZN(new_n1129));
  NAND4_X1  g703(.A1(new_n932), .A2(new_n882), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g704(.A(G227), .ZN(new_n1131));
  NAND2_X1  g705(.A1(new_n1131), .A2(G319), .ZN(new_n1132));
  XOR2_X1   g706(.A(new_n1132), .B(KEYINPUT127), .Z(new_n1133));
  NOR2_X1   g707(.A1(new_n1130), .A2(new_n1133), .ZN(G308));
  AND2_X1   g708(.A1(new_n882), .A2(new_n1129), .ZN(new_n1135));
  INV_X1    g709(.A(new_n1133), .ZN(new_n1136));
  NAND4_X1  g710(.A1(new_n1135), .A2(new_n1128), .A3(new_n932), .A4(new_n1136), .ZN(G225));
endmodule


