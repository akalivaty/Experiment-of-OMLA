

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733;

  NAND2_X2 U366 ( .A1(n371), .A2(n368), .ZN(n579) );
  XNOR2_X2 U367 ( .A(n570), .B(n569), .ZN(n727) );
  AND2_X2 U368 ( .A1(n583), .A2(n568), .ZN(n570) );
  XNOR2_X2 U369 ( .A(n549), .B(KEYINPUT1), .ZN(n583) );
  XNOR2_X2 U370 ( .A(n430), .B(n391), .ZN(n549) );
  NAND2_X1 U371 ( .A1(n394), .A2(n732), .ZN(n381) );
  INV_X1 U372 ( .A(n656), .ZN(n390) );
  OR2_X2 U373 ( .A1(n609), .A2(G902), .ZN(n441) );
  OR2_X1 U374 ( .A1(n676), .A2(n556), .ZN(n553) );
  XNOR2_X1 U375 ( .A(n534), .B(KEYINPUT74), .ZN(n559) );
  NOR2_X1 U376 ( .A1(n566), .A2(n580), .ZN(n567) );
  NAND2_X1 U377 ( .A1(n533), .A2(n399), .ZN(n534) );
  AND2_X1 U378 ( .A1(n501), .A2(n384), .ZN(n383) );
  XNOR2_X1 U379 ( .A(n400), .B(KEYINPUT75), .ZN(n399) );
  XNOR2_X1 U380 ( .A(n363), .B(n362), .ZN(n508) );
  XNOR2_X1 U381 ( .A(n545), .B(KEYINPUT6), .ZN(n562) );
  INV_X1 U382 ( .A(KEYINPUT64), .ZN(n414) );
  XNOR2_X1 U383 ( .A(G113), .B(KEYINPUT69), .ZN(n377) );
  XNOR2_X1 U384 ( .A(G137), .B(G131), .ZN(n423) );
  AND2_X2 U385 ( .A1(n549), .A2(n390), .ZN(n529) );
  BUF_X1 U386 ( .A(n535), .Z(n585) );
  NOR2_X2 U387 ( .A1(n695), .A2(G902), .ZN(n402) );
  XNOR2_X1 U388 ( .A(n460), .B(n461), .ZN(n591) );
  XNOR2_X1 U389 ( .A(n366), .B(n365), .ZN(n695) );
  XNOR2_X1 U390 ( .A(n376), .B(n432), .ZN(n457) );
  XOR2_X1 U391 ( .A(KEYINPUT3), .B(G119), .Z(n432) );
  XNOR2_X1 U392 ( .A(n377), .B(n431), .ZN(n376) );
  INV_X1 U393 ( .A(G116), .ZN(n431) );
  XOR2_X1 U394 ( .A(G146), .B(G125), .Z(n451) );
  NAND2_X1 U395 ( .A1(n493), .A2(G221), .ZN(n367) );
  INV_X1 U396 ( .A(KEYINPUT33), .ZN(n392) );
  NAND2_X1 U397 ( .A1(n508), .A2(n562), .ZN(n393) );
  XNOR2_X1 U398 ( .A(KEYINPUT66), .B(KEYINPUT4), .ZN(n452) );
  XNOR2_X1 U399 ( .A(KEYINPUT65), .B(G101), .ZN(n435) );
  INV_X1 U400 ( .A(KEYINPUT44), .ZN(n378) );
  XOR2_X1 U401 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n449) );
  INV_X1 U402 ( .A(KEYINPUT39), .ZN(n373) );
  OR2_X1 U403 ( .A1(n646), .A2(n373), .ZN(n372) );
  XNOR2_X1 U404 ( .A(n375), .B(n348), .ZN(n535) );
  NAND2_X1 U405 ( .A1(n591), .A2(n589), .ZN(n375) );
  XNOR2_X1 U406 ( .A(n544), .B(KEYINPUT68), .ZN(n564) );
  INV_X1 U407 ( .A(KEYINPUT28), .ZN(n546) );
  OR2_X2 U408 ( .A1(n557), .A2(n345), .ZN(n384) );
  AND2_X1 U409 ( .A1(n386), .A2(n387), .ZN(n385) );
  INV_X1 U410 ( .A(G469), .ZN(n391) );
  NOR2_X1 U411 ( .A1(G902), .A2(n688), .ZN(n430) );
  XNOR2_X1 U412 ( .A(G107), .B(G110), .ZN(n425) );
  XNOR2_X1 U413 ( .A(n457), .B(n456), .ZN(n708) );
  XOR2_X1 U414 ( .A(KEYINPUT16), .B(KEYINPUT71), .Z(n455) );
  XOR2_X1 U415 ( .A(KEYINPUT23), .B(G119), .Z(n412) );
  XNOR2_X1 U416 ( .A(G128), .B(G110), .ZN(n411) );
  XNOR2_X1 U417 ( .A(n451), .B(n410), .ZN(n717) );
  XNOR2_X1 U418 ( .A(G140), .B(KEYINPUT10), .ZN(n410) );
  XNOR2_X1 U419 ( .A(G137), .B(KEYINPUT91), .ZN(n416) );
  XOR2_X1 U420 ( .A(KEYINPUT80), .B(KEYINPUT24), .Z(n417) );
  XNOR2_X1 U421 ( .A(n397), .B(n415), .ZN(n493) );
  XNOR2_X1 U422 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n415) );
  XNOR2_X1 U423 ( .A(G122), .B(G104), .ZN(n477) );
  INV_X1 U424 ( .A(n717), .ZN(n481) );
  XNOR2_X1 U425 ( .A(n472), .B(n471), .ZN(n474) );
  AND2_X1 U426 ( .A1(n360), .A2(n349), .ZN(n358) );
  XNOR2_X1 U427 ( .A(n420), .B(KEYINPUT25), .ZN(n401) );
  XNOR2_X1 U428 ( .A(n487), .B(n486), .ZN(n517) );
  NOR2_X1 U429 ( .A1(G953), .A2(G237), .ZN(n475) );
  NAND2_X1 U430 ( .A1(G237), .A2(G234), .ZN(n442) );
  INV_X1 U431 ( .A(G237), .ZN(n462) );
  INV_X1 U432 ( .A(KEYINPUT72), .ZN(n362) );
  NAND2_X1 U433 ( .A1(n583), .A2(n390), .ZN(n363) );
  INV_X1 U434 ( .A(KEYINPUT45), .ZN(n395) );
  XOR2_X1 U435 ( .A(KEYINPUT9), .B(G107), .Z(n489) );
  XNOR2_X1 U436 ( .A(n439), .B(n429), .ZN(n688) );
  XNOR2_X1 U437 ( .A(n708), .B(n459), .ZN(n460) );
  INV_X1 U438 ( .A(n458), .ZN(n459) );
  NAND2_X1 U439 ( .A1(n370), .A2(n369), .ZN(n368) );
  AND2_X1 U440 ( .A1(n374), .A2(n372), .ZN(n371) );
  AND2_X1 U441 ( .A1(n646), .A2(n373), .ZN(n369) );
  XNOR2_X1 U442 ( .A(n546), .B(KEYINPUT105), .ZN(n547) );
  XNOR2_X1 U443 ( .A(n388), .B(KEYINPUT22), .ZN(n504) );
  INV_X1 U444 ( .A(n583), .ZN(n657) );
  XNOR2_X1 U445 ( .A(n413), .B(n418), .ZN(n365) );
  XNOR2_X1 U446 ( .A(n367), .B(n717), .ZN(n366) );
  XNOR2_X1 U447 ( .A(n483), .B(n482), .ZN(n604) );
  XNOR2_X1 U448 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U449 ( .A(G143), .B(G131), .ZN(n473) );
  BUF_X1 U450 ( .A(n687), .Z(n694) );
  NAND2_X1 U451 ( .A1(n361), .A2(n346), .ZN(n498) );
  NAND2_X1 U452 ( .A1(n358), .A2(n355), .ZN(n361) );
  NAND2_X1 U453 ( .A1(n357), .A2(n356), .ZN(n355) );
  NOR2_X1 U454 ( .A1(n557), .A2(n556), .ZN(n628) );
  OR2_X1 U455 ( .A1(n466), .A2(KEYINPUT0), .ZN(n345) );
  NOR2_X1 U456 ( .A1(n517), .A2(n514), .ZN(n346) );
  XOR2_X1 U457 ( .A(n451), .B(n450), .Z(n347) );
  AND2_X1 U458 ( .A1(n464), .A2(G210), .ZN(n348) );
  OR2_X1 U459 ( .A1(n467), .A2(n359), .ZN(n349) );
  AND2_X1 U460 ( .A1(n523), .A2(n617), .ZN(n350) );
  XOR2_X1 U461 ( .A(KEYINPUT82), .B(KEYINPUT48), .Z(n351) );
  AND2_X1 U462 ( .A1(n590), .A2(n588), .ZN(n352) );
  AND2_X1 U463 ( .A1(n590), .A2(KEYINPUT2), .ZN(n353) );
  XNOR2_X2 U464 ( .A(n538), .B(KEYINPUT40), .ZN(n603) );
  NAND2_X1 U465 ( .A1(n577), .A2(n354), .ZN(n578) );
  AND2_X1 U466 ( .A1(n575), .A2(n576), .ZN(n354) );
  NOR2_X1 U467 ( .A1(n511), .A2(n468), .ZN(n356) );
  INV_X1 U468 ( .A(n677), .ZN(n357) );
  INV_X1 U469 ( .A(n468), .ZN(n359) );
  NAND2_X1 U470 ( .A1(n677), .A2(n468), .ZN(n360) );
  NOR2_X2 U471 ( .A1(n723), .A2(n700), .ZN(n639) );
  XNOR2_X2 U472 ( .A(n642), .B(KEYINPUT81), .ZN(n723) );
  AND2_X2 U473 ( .A1(n364), .A2(n406), .ZN(n642) );
  XNOR2_X1 U474 ( .A(n578), .B(n351), .ZN(n364) );
  INV_X1 U475 ( .A(n559), .ZN(n370) );
  NAND2_X1 U476 ( .A1(n559), .A2(KEYINPUT39), .ZN(n374) );
  NAND2_X1 U477 ( .A1(n579), .A2(n632), .ZN(n538) );
  NAND2_X1 U478 ( .A1(n535), .A2(n645), .ZN(n566) );
  XNOR2_X1 U479 ( .A(n379), .B(n378), .ZN(n389) );
  NAND2_X1 U480 ( .A1(n382), .A2(n380), .ZN(n379) );
  XNOR2_X1 U481 ( .A(n381), .B(KEYINPUT85), .ZN(n380) );
  INV_X1 U482 ( .A(n730), .ZN(n382) );
  NAND2_X1 U483 ( .A1(n385), .A2(n384), .ZN(n511) );
  NAND2_X1 U484 ( .A1(n383), .A2(n385), .ZN(n388) );
  NAND2_X1 U485 ( .A1(n557), .A2(KEYINPUT0), .ZN(n386) );
  NAND2_X1 U486 ( .A1(n466), .A2(KEYINPUT0), .ZN(n387) );
  XNOR2_X2 U487 ( .A(n441), .B(n440), .ZN(n545) );
  NAND2_X1 U488 ( .A1(n389), .A2(n350), .ZN(n396) );
  XNOR2_X2 U489 ( .A(n498), .B(KEYINPUT35), .ZN(n730) );
  XNOR2_X2 U490 ( .A(n393), .B(n392), .ZN(n677) );
  XNOR2_X1 U491 ( .A(n394), .B(G119), .ZN(G21) );
  XNOR2_X2 U492 ( .A(n503), .B(KEYINPUT32), .ZN(n394) );
  XNOR2_X2 U493 ( .A(n566), .B(n465), .ZN(n557) );
  XNOR2_X2 U494 ( .A(n396), .B(n395), .ZN(n700) );
  NAND2_X1 U495 ( .A1(n447), .A2(G234), .ZN(n397) );
  XNOR2_X2 U496 ( .A(n414), .B(G953), .ZN(n447) );
  NAND2_X1 U497 ( .A1(n398), .A2(n642), .ZN(n681) );
  INV_X1 U498 ( .A(n700), .ZN(n398) );
  NAND2_X1 U499 ( .A1(n529), .A2(n541), .ZN(n400) );
  XNOR2_X2 U500 ( .A(n402), .B(n401), .ZN(n660) );
  XNOR2_X2 U501 ( .A(n403), .B(G146), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n403), .B(n718), .ZN(n721) );
  XNOR2_X2 U503 ( .A(n491), .B(n424), .ZN(n403) );
  NAND2_X1 U504 ( .A1(n687), .A2(G478), .ZN(n599) );
  NAND2_X2 U505 ( .A1(n404), .A2(n405), .ZN(n687) );
  NAND2_X1 U506 ( .A1(n639), .A2(n352), .ZN(n404) );
  NAND2_X1 U507 ( .A1(n681), .A2(n353), .ZN(n405) );
  XNOR2_X2 U508 ( .A(n453), .B(G134), .ZN(n491) );
  AND2_X1 U509 ( .A1(n602), .A2(n587), .ZN(n406) );
  INV_X1 U510 ( .A(G113), .ZN(n469) );
  XNOR2_X1 U511 ( .A(n470), .B(n469), .ZN(n472) );
  XNOR2_X1 U512 ( .A(KEYINPUT103), .B(n500), .ZN(n501) );
  XNOR2_X1 U513 ( .A(n455), .B(G122), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n485), .B(n484), .ZN(n486) );
  OR2_X1 U515 ( .A1(n447), .A2(G952), .ZN(n612) );
  XOR2_X1 U516 ( .A(KEYINPUT70), .B(KEYINPUT34), .Z(n468) );
  XOR2_X1 U517 ( .A(KEYINPUT21), .B(KEYINPUT92), .Z(n409) );
  XNOR2_X1 U518 ( .A(KEYINPUT15), .B(G902), .ZN(n589) );
  NAND2_X1 U519 ( .A1(G234), .A2(n589), .ZN(n407) );
  XNOR2_X1 U520 ( .A(KEYINPUT20), .B(n407), .ZN(n419) );
  NAND2_X1 U521 ( .A1(n419), .A2(G221), .ZN(n408) );
  XNOR2_X1 U522 ( .A(n409), .B(n408), .ZN(n659) );
  XNOR2_X1 U523 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U524 ( .A(n417), .B(n416), .ZN(n418) );
  NAND2_X1 U525 ( .A1(n419), .A2(G217), .ZN(n420) );
  NAND2_X1 U526 ( .A1(n659), .A2(n660), .ZN(n656) );
  XNOR2_X2 U527 ( .A(KEYINPUT76), .B(G143), .ZN(n422) );
  INV_X1 U528 ( .A(G128), .ZN(n421) );
  XNOR2_X2 U529 ( .A(n422), .B(n421), .ZN(n453) );
  XNOR2_X1 U530 ( .A(n452), .B(n423), .ZN(n424) );
  XNOR2_X1 U531 ( .A(n425), .B(G104), .ZN(n709) );
  XNOR2_X1 U532 ( .A(n709), .B(n435), .ZN(n458) );
  XOR2_X1 U533 ( .A(G140), .B(KEYINPUT90), .Z(n427) );
  NAND2_X1 U534 ( .A1(G227), .A2(n447), .ZN(n426) );
  XNOR2_X1 U535 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U536 ( .A(n458), .B(n428), .ZN(n429) );
  NAND2_X1 U537 ( .A1(n475), .A2(G210), .ZN(n434) );
  XNOR2_X1 U538 ( .A(KEYINPUT73), .B(KEYINPUT5), .ZN(n433) );
  XNOR2_X1 U539 ( .A(n434), .B(n433), .ZN(n436) );
  XNOR2_X1 U540 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U541 ( .A(n457), .B(n437), .ZN(n438) );
  XNOR2_X1 U542 ( .A(n439), .B(n438), .ZN(n609) );
  XNOR2_X1 U543 ( .A(G472), .B(KEYINPUT93), .ZN(n440) );
  XOR2_X1 U544 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n443) );
  XNOR2_X1 U545 ( .A(n443), .B(n442), .ZN(n444) );
  NAND2_X1 U546 ( .A1(G952), .A2(n444), .ZN(n674) );
  NOR2_X1 U547 ( .A1(G953), .A2(n674), .ZN(n527) );
  NAND2_X1 U548 ( .A1(n444), .A2(G902), .ZN(n445) );
  XOR2_X1 U549 ( .A(n445), .B(KEYINPUT89), .Z(n524) );
  XOR2_X1 U550 ( .A(KEYINPUT88), .B(G898), .Z(n704) );
  NAND2_X1 U551 ( .A1(G953), .A2(n704), .ZN(n713) );
  NOR2_X1 U552 ( .A1(n524), .A2(n713), .ZN(n446) );
  NOR2_X1 U553 ( .A1(n527), .A2(n446), .ZN(n466) );
  INV_X1 U554 ( .A(KEYINPUT19), .ZN(n465) );
  NAND2_X1 U555 ( .A1(G224), .A2(n447), .ZN(n448) );
  XNOR2_X1 U556 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U557 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U558 ( .A(n347), .B(n454), .ZN(n461) );
  INV_X1 U559 ( .A(G902), .ZN(n463) );
  NAND2_X1 U560 ( .A1(n463), .A2(n462), .ZN(n464) );
  NAND2_X1 U561 ( .A1(n464), .A2(G214), .ZN(n645) );
  INV_X1 U562 ( .A(n511), .ZN(n467) );
  XNOR2_X1 U563 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n470) );
  XOR2_X1 U564 ( .A(KEYINPUT96), .B(KEYINPUT99), .Z(n471) );
  XNOR2_X1 U565 ( .A(n474), .B(n473), .ZN(n483) );
  NAND2_X1 U566 ( .A1(n475), .A2(G214), .ZN(n476) );
  XNOR2_X1 U567 ( .A(n477), .B(n476), .ZN(n479) );
  XOR2_X1 U568 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n478) );
  XNOR2_X1 U569 ( .A(n479), .B(n478), .ZN(n480) );
  NOR2_X1 U570 ( .A1(G902), .A2(n604), .ZN(n487) );
  XNOR2_X1 U571 ( .A(KEYINPUT13), .B(KEYINPUT100), .ZN(n485) );
  INV_X1 U572 ( .A(G475), .ZN(n484) );
  XNOR2_X1 U573 ( .A(G116), .B(G122), .ZN(n488) );
  XNOR2_X1 U574 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U575 ( .A(n490), .B(KEYINPUT101), .Z(n492) );
  XNOR2_X1 U576 ( .A(n491), .B(n492), .ZN(n496) );
  NAND2_X1 U577 ( .A1(n493), .A2(G217), .ZN(n494) );
  XNOR2_X1 U578 ( .A(n494), .B(KEYINPUT7), .ZN(n495) );
  XNOR2_X1 U579 ( .A(n496), .B(n495), .ZN(n598) );
  NOR2_X1 U580 ( .A1(n598), .A2(G902), .ZN(n497) );
  XNOR2_X1 U581 ( .A(G478), .B(n497), .ZN(n514) );
  NAND2_X1 U582 ( .A1(n517), .A2(n514), .ZN(n648) );
  INV_X1 U583 ( .A(n648), .ZN(n499) );
  NAND2_X1 U584 ( .A1(n659), .A2(n499), .ZN(n500) );
  NOR2_X1 U585 ( .A1(n504), .A2(n562), .ZN(n520) );
  NOR2_X1 U586 ( .A1(n660), .A2(n657), .ZN(n502) );
  NAND2_X1 U587 ( .A1(n520), .A2(n502), .ZN(n503) );
  NOR2_X1 U588 ( .A1(n504), .A2(n583), .ZN(n506) );
  INV_X1 U589 ( .A(n545), .ZN(n662) );
  INV_X1 U590 ( .A(n660), .ZN(n542) );
  AND2_X1 U591 ( .A1(n545), .A2(n542), .ZN(n505) );
  NAND2_X1 U592 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U593 ( .A(n507), .B(KEYINPUT104), .ZN(n732) );
  NAND2_X1 U594 ( .A1(n508), .A2(n662), .ZN(n667) );
  NOR2_X1 U595 ( .A1(n511), .A2(n667), .ZN(n510) );
  XOR2_X1 U596 ( .A(KEYINPUT31), .B(KEYINPUT94), .Z(n509) );
  XNOR2_X1 U597 ( .A(n510), .B(n509), .ZN(n635) );
  NAND2_X1 U598 ( .A1(n529), .A2(n467), .ZN(n512) );
  NOR2_X1 U599 ( .A1(n512), .A2(n662), .ZN(n620) );
  NOR2_X1 U600 ( .A1(n635), .A2(n620), .ZN(n513) );
  XNOR2_X1 U601 ( .A(n513), .B(KEYINPUT95), .ZN(n519) );
  INV_X1 U602 ( .A(n514), .ZN(n516) );
  NAND2_X1 U603 ( .A1(n517), .A2(n516), .ZN(n515) );
  XOR2_X1 U604 ( .A(n515), .B(KEYINPUT102), .Z(n634) );
  INV_X1 U605 ( .A(n634), .ZN(n518) );
  OR2_X1 U606 ( .A1(n517), .A2(n516), .ZN(n537) );
  NAND2_X1 U607 ( .A1(n518), .A2(n537), .ZN(n649) );
  NAND2_X1 U608 ( .A1(n519), .A2(n649), .ZN(n523) );
  XOR2_X1 U609 ( .A(n520), .B(KEYINPUT84), .Z(n521) );
  NOR2_X1 U610 ( .A1(n542), .A2(n521), .ZN(n522) );
  NAND2_X1 U611 ( .A1(n657), .A2(n522), .ZN(n617) );
  OR2_X1 U612 ( .A1(n447), .A2(n524), .ZN(n525) );
  NOR2_X1 U613 ( .A1(G900), .A2(n525), .ZN(n526) );
  NOR2_X1 U614 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U615 ( .A(KEYINPUT77), .B(n528), .ZN(n541) );
  INV_X1 U616 ( .A(n645), .ZN(n530) );
  OR2_X1 U617 ( .A1(n545), .A2(n530), .ZN(n532) );
  INV_X1 U618 ( .A(KEYINPUT30), .ZN(n531) );
  XNOR2_X1 U619 ( .A(n532), .B(n531), .ZN(n533) );
  INV_X1 U620 ( .A(KEYINPUT38), .ZN(n536) );
  XNOR2_X1 U621 ( .A(n585), .B(n536), .ZN(n646) );
  INV_X1 U622 ( .A(n537), .ZN(n632) );
  NAND2_X1 U623 ( .A1(n646), .A2(n645), .ZN(n650) );
  NOR2_X1 U624 ( .A1(n648), .A2(n650), .ZN(n540) );
  XNOR2_X1 U625 ( .A(KEYINPUT41), .B(KEYINPUT106), .ZN(n539) );
  XNOR2_X1 U626 ( .A(n540), .B(n539), .ZN(n676) );
  AND2_X1 U627 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U628 ( .A1(n543), .A2(n659), .ZN(n544) );
  NOR2_X1 U629 ( .A1(n564), .A2(n545), .ZN(n548) );
  XNOR2_X1 U630 ( .A(n548), .B(n547), .ZN(n550) );
  NAND2_X1 U631 ( .A1(n550), .A2(n549), .ZN(n556) );
  INV_X1 U632 ( .A(KEYINPUT107), .ZN(n551) );
  XNOR2_X1 U633 ( .A(n551), .B(KEYINPUT42), .ZN(n552) );
  XNOR2_X1 U634 ( .A(n553), .B(n552), .ZN(n731) );
  NAND2_X1 U635 ( .A1(n603), .A2(n731), .ZN(n555) );
  XNOR2_X1 U636 ( .A(KEYINPUT83), .B(KEYINPUT46), .ZN(n554) );
  XNOR2_X1 U637 ( .A(n555), .B(n554), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n628), .A2(n649), .ZN(n571) );
  NAND2_X1 U639 ( .A1(n571), .A2(KEYINPUT47), .ZN(n560) );
  NAND2_X1 U640 ( .A1(n585), .A2(n346), .ZN(n558) );
  OR2_X1 U641 ( .A1(n559), .A2(n558), .ZN(n627) );
  NAND2_X1 U642 ( .A1(n560), .A2(n627), .ZN(n561) );
  XNOR2_X1 U643 ( .A(n561), .B(KEYINPUT79), .ZN(n576) );
  INV_X1 U644 ( .A(n562), .ZN(n563) );
  NOR2_X1 U645 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U646 ( .A1(n632), .A2(n565), .ZN(n580) );
  XNOR2_X1 U647 ( .A(KEYINPUT36), .B(n567), .ZN(n568) );
  INV_X1 U648 ( .A(KEYINPUT108), .ZN(n569) );
  INV_X1 U649 ( .A(n571), .ZN(n573) );
  INV_X1 U650 ( .A(KEYINPUT47), .ZN(n572) );
  NAND2_X1 U651 ( .A1(n573), .A2(n572), .ZN(n574) );
  AND2_X1 U652 ( .A1(n727), .A2(n574), .ZN(n575) );
  NAND2_X1 U653 ( .A1(n579), .A2(n634), .ZN(n602) );
  INV_X1 U654 ( .A(n580), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n581), .A2(n645), .ZN(n582) );
  NOR2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U657 ( .A(n584), .B(KEYINPUT43), .ZN(n586) );
  NOR2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n638) );
  INV_X1 U659 ( .A(n638), .ZN(n587) );
  INV_X1 U660 ( .A(KEYINPUT2), .ZN(n588) );
  INV_X1 U661 ( .A(n589), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n687), .A2(G210), .ZN(n595) );
  XNOR2_X1 U663 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n593) );
  XNOR2_X1 U664 ( .A(n591), .B(KEYINPUT118), .ZN(n592) );
  XNOR2_X1 U665 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U666 ( .A(n595), .B(n594), .ZN(n596) );
  INV_X1 U667 ( .A(n612), .ZN(n699) );
  NOR2_X2 U668 ( .A1(n596), .A2(n699), .ZN(n597) );
  XNOR2_X1 U669 ( .A(n597), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U670 ( .A(n599), .B(n598), .ZN(n600) );
  NOR2_X2 U671 ( .A1(n600), .A2(n699), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n601), .B(KEYINPUT120), .ZN(G63) );
  XNOR2_X1 U673 ( .A(n602), .B(G134), .ZN(G36) );
  XNOR2_X1 U674 ( .A(n603), .B(G131), .ZN(G33) );
  NAND2_X1 U675 ( .A1(n687), .A2(G475), .ZN(n606) );
  XOR2_X1 U676 ( .A(n604), .B(KEYINPUT59), .Z(n605) );
  XNOR2_X1 U677 ( .A(n606), .B(n605), .ZN(n607) );
  NOR2_X2 U678 ( .A1(n607), .A2(n699), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n608), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U680 ( .A1(n687), .A2(G472), .ZN(n611) );
  XOR2_X1 U681 ( .A(KEYINPUT62), .B(n609), .Z(n610) );
  XNOR2_X1 U682 ( .A(n611), .B(n610), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n613), .A2(n612), .ZN(n615) );
  XNOR2_X1 U684 ( .A(KEYINPUT86), .B(KEYINPUT63), .ZN(n614) );
  XNOR2_X1 U685 ( .A(n615), .B(n614), .ZN(G57) );
  XOR2_X1 U686 ( .A(G101), .B(KEYINPUT109), .Z(n616) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(G3) );
  NAND2_X1 U688 ( .A1(n620), .A2(n632), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n618), .B(KEYINPUT110), .ZN(n619) );
  XNOR2_X1 U690 ( .A(G104), .B(n619), .ZN(G6) );
  XOR2_X1 U691 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n622) );
  NAND2_X1 U692 ( .A1(n620), .A2(n634), .ZN(n621) );
  XNOR2_X1 U693 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U694 ( .A(G107), .B(n623), .ZN(G9) );
  XOR2_X1 U695 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n625) );
  NAND2_X1 U696 ( .A1(n628), .A2(n634), .ZN(n624) );
  XNOR2_X1 U697 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U698 ( .A(G128), .B(n626), .ZN(G30) );
  XNOR2_X1 U699 ( .A(G143), .B(n627), .ZN(G45) );
  XOR2_X1 U700 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n630) );
  NAND2_X1 U701 ( .A1(n628), .A2(n632), .ZN(n629) );
  XNOR2_X1 U702 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U703 ( .A(G146), .B(n631), .ZN(G48) );
  NAND2_X1 U704 ( .A1(n635), .A2(n632), .ZN(n633) );
  XNOR2_X1 U705 ( .A(n633), .B(G113), .ZN(G15) );
  XOR2_X1 U706 ( .A(G116), .B(KEYINPUT115), .Z(n637) );
  NAND2_X1 U707 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n637), .B(n636), .ZN(G18) );
  XOR2_X1 U709 ( .A(G140), .B(n638), .Z(G42) );
  INV_X1 U710 ( .A(n639), .ZN(n641) );
  OR2_X1 U711 ( .A1(KEYINPUT2), .A2(KEYINPUT78), .ZN(n640) );
  NAND2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U713 ( .A1(n642), .A2(KEYINPUT2), .ZN(n643) );
  NAND2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n685) );
  NOR2_X1 U715 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U716 ( .A1(n648), .A2(n647), .ZN(n653) );
  INV_X1 U717 ( .A(n649), .ZN(n651) );
  NOR2_X1 U718 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U719 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U720 ( .A(KEYINPUT117), .B(n654), .Z(n655) );
  NOR2_X1 U721 ( .A1(n677), .A2(n655), .ZN(n671) );
  NAND2_X1 U722 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U723 ( .A(n658), .B(KEYINPUT50), .ZN(n665) );
  NOR2_X1 U724 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U725 ( .A(KEYINPUT49), .B(n661), .Z(n663) );
  NOR2_X1 U726 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U727 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U728 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U729 ( .A(KEYINPUT51), .B(n668), .ZN(n669) );
  NOR2_X1 U730 ( .A1(n676), .A2(n669), .ZN(n670) );
  NOR2_X1 U731 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U732 ( .A(n672), .B(KEYINPUT52), .ZN(n673) );
  NOR2_X1 U733 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U734 ( .A1(G953), .A2(n675), .ZN(n679) );
  OR2_X1 U735 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U736 ( .A1(n679), .A2(n678), .ZN(n683) );
  AND2_X1 U737 ( .A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(n680) );
  AND2_X1 U738 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U739 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U740 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U741 ( .A(KEYINPUT53), .B(n686), .Z(G75) );
  NAND2_X1 U742 ( .A1(n694), .A2(G469), .ZN(n692) );
  XNOR2_X1 U743 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n690) );
  XNOR2_X1 U744 ( .A(n688), .B(KEYINPUT57), .ZN(n689) );
  XNOR2_X1 U745 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U746 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U747 ( .A1(n699), .A2(n693), .ZN(G54) );
  NAND2_X1 U748 ( .A1(n694), .A2(G217), .ZN(n697) );
  XOR2_X1 U749 ( .A(n695), .B(KEYINPUT121), .Z(n696) );
  XNOR2_X1 U750 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U751 ( .A1(n699), .A2(n698), .ZN(G66) );
  NOR2_X1 U752 ( .A1(n700), .A2(G953), .ZN(n701) );
  XOR2_X1 U753 ( .A(KEYINPUT123), .B(n701), .Z(n707) );
  NAND2_X1 U754 ( .A1(G953), .A2(G224), .ZN(n702) );
  XOR2_X1 U755 ( .A(KEYINPUT61), .B(n702), .Z(n703) );
  NOR2_X1 U756 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U757 ( .A(KEYINPUT122), .B(n705), .ZN(n706) );
  NOR2_X1 U758 ( .A1(n707), .A2(n706), .ZN(n716) );
  XOR2_X1 U759 ( .A(KEYINPUT125), .B(n708), .Z(n711) );
  XNOR2_X1 U760 ( .A(G101), .B(n709), .ZN(n710) );
  XNOR2_X1 U761 ( .A(n711), .B(n710), .ZN(n712) );
  NAND2_X1 U762 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U763 ( .A(n714), .B(KEYINPUT124), .ZN(n715) );
  XNOR2_X1 U764 ( .A(n716), .B(n715), .ZN(G69) );
  XNOR2_X1 U765 ( .A(n717), .B(KEYINPUT126), .ZN(n718) );
  XOR2_X1 U766 ( .A(G227), .B(n721), .Z(n719) );
  NAND2_X1 U767 ( .A1(n719), .A2(G900), .ZN(n720) );
  NAND2_X1 U768 ( .A1(G953), .A2(n720), .ZN(n726) );
  XNOR2_X1 U769 ( .A(n721), .B(KEYINPUT127), .ZN(n722) );
  XNOR2_X1 U770 ( .A(n723), .B(n722), .ZN(n724) );
  NAND2_X1 U771 ( .A1(n724), .A2(n447), .ZN(n725) );
  NAND2_X1 U772 ( .A1(n726), .A2(n725), .ZN(G72) );
  XOR2_X1 U773 ( .A(KEYINPUT37), .B(KEYINPUT116), .Z(n729) );
  XNOR2_X1 U774 ( .A(G125), .B(n727), .ZN(n728) );
  XNOR2_X1 U775 ( .A(n729), .B(n728), .ZN(G27) );
  XOR2_X1 U776 ( .A(n730), .B(G122), .Z(G24) );
  XNOR2_X1 U777 ( .A(G137), .B(n731), .ZN(G39) );
  XOR2_X1 U778 ( .A(n732), .B(G110), .Z(n733) );
  XNOR2_X1 U779 ( .A(KEYINPUT111), .B(n733), .ZN(G12) );
endmodule

