

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U556 ( .A(KEYINPUT66), .B(n550), .Z(G160) );
  XNOR2_X1 U557 ( .A(n542), .B(n541), .ZN(G164) );
  BUF_X1 U558 ( .A(n880), .Z(n524) );
  XNOR2_X1 U559 ( .A(n536), .B(KEYINPUT67), .ZN(n880) );
  NOR2_X1 U560 ( .A1(G1384), .A2(G164), .ZN(n784) );
  NOR2_X1 U561 ( .A1(n538), .A2(n526), .ZN(n539) );
  NOR2_X1 U562 ( .A1(n815), .A2(n528), .ZN(n525) );
  XOR2_X1 U563 ( .A(KEYINPUT88), .B(n537), .Z(n526) );
  XNOR2_X1 U564 ( .A(n566), .B(KEYINPUT13), .ZN(n527) );
  INV_X1 U565 ( .A(G2105), .ZN(n535) );
  AND2_X1 U566 ( .A1(n997), .A2(n826), .ZN(n528) );
  AND2_X1 U567 ( .A1(n796), .A2(n822), .ZN(n529) );
  NOR2_X1 U568 ( .A1(n718), .A2(n717), .ZN(n719) );
  INV_X1 U569 ( .A(KEYINPUT29), .ZN(n725) );
  NOR2_X1 U570 ( .A1(n738), .A2(n737), .ZN(n739) );
  AND2_X1 U571 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U572 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U573 ( .A1(n784), .A2(n691), .ZN(n743) );
  NOR2_X1 U574 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U575 ( .A1(n983), .A2(n771), .ZN(n772) );
  NOR2_X1 U576 ( .A1(n773), .A2(n772), .ZN(n782) );
  NOR2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  NOR2_X1 U578 ( .A1(G651), .A2(n552), .ZN(n657) );
  NOR2_X1 U579 ( .A1(G651), .A2(G543), .ZN(n658) );
  NOR2_X1 U580 ( .A1(n570), .A2(n569), .ZN(n571) );
  INV_X1 U581 ( .A(KEYINPUT90), .ZN(n542) );
  XOR2_X1 U582 ( .A(KEYINPUT68), .B(n530), .Z(n531) );
  XNOR2_X1 U583 ( .A(KEYINPUT17), .B(n531), .ZN(n622) );
  NAND2_X1 U584 ( .A1(G138), .A2(n622), .ZN(n532) );
  XOR2_X1 U585 ( .A(KEYINPUT89), .B(n532), .Z(n540) );
  NOR2_X1 U586 ( .A1(G2104), .A2(n535), .ZN(n884) );
  NAND2_X1 U587 ( .A1(G126), .A2(n884), .ZN(n534) );
  AND2_X1 U588 ( .A1(G2105), .A2(G2104), .ZN(n885) );
  NAND2_X1 U589 ( .A1(G114), .A2(n885), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U591 ( .A1(n535), .A2(G2104), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n880), .A2(G102), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n884), .A2(G125), .ZN(n549) );
  NAND2_X1 U595 ( .A1(G137), .A2(n622), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G113), .A2(n885), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n547) );
  NAND2_X1 U598 ( .A1(G101), .A2(n880), .ZN(n545) );
  XNOR2_X1 U599 ( .A(KEYINPUT23), .B(n545), .ZN(n546) );
  NOR2_X1 U600 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U601 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U602 ( .A(KEYINPUT0), .B(G543), .Z(n552) );
  NAND2_X1 U603 ( .A1(G52), .A2(n657), .ZN(n551) );
  XNOR2_X1 U604 ( .A(n551), .B(KEYINPUT71), .ZN(n562) );
  NAND2_X1 U605 ( .A1(G90), .A2(n658), .ZN(n555) );
  INV_X1 U606 ( .A(G651), .ZN(n557) );
  OR2_X1 U607 ( .A1(n557), .A2(n552), .ZN(n553) );
  XNOR2_X2 U608 ( .A(KEYINPUT69), .B(n553), .ZN(n654) );
  NAND2_X1 U609 ( .A1(G77), .A2(n654), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U611 ( .A(n556), .B(KEYINPUT9), .ZN(n560) );
  NOR2_X1 U612 ( .A1(G543), .A2(n557), .ZN(n558) );
  XOR2_X1 U613 ( .A(KEYINPUT1), .B(n558), .Z(n663) );
  NAND2_X1 U614 ( .A1(G64), .A2(n663), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U616 ( .A1(n562), .A2(n561), .ZN(G171) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U618 ( .A(G860), .ZN(n633) );
  NAND2_X1 U619 ( .A1(n658), .A2(G81), .ZN(n563) );
  XNOR2_X1 U620 ( .A(n563), .B(KEYINPUT12), .ZN(n565) );
  NAND2_X1 U621 ( .A1(G68), .A2(n654), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U623 ( .A1(G43), .A2(n657), .ZN(n567) );
  NAND2_X1 U624 ( .A1(n527), .A2(n567), .ZN(n570) );
  NAND2_X1 U625 ( .A1(n663), .A2(G56), .ZN(n568) );
  XOR2_X1 U626 ( .A(KEYINPUT14), .B(n568), .Z(n569) );
  XOR2_X1 U627 ( .A(KEYINPUT72), .B(n571), .Z(n981) );
  OR2_X1 U628 ( .A1(n633), .A2(n981), .ZN(G153) );
  INV_X1 U629 ( .A(G120), .ZN(G236) );
  INV_X1 U630 ( .A(G69), .ZN(G235) );
  INV_X1 U631 ( .A(G108), .ZN(G238) );
  NAND2_X1 U632 ( .A1(n657), .A2(G50), .ZN(n572) );
  XOR2_X1 U633 ( .A(KEYINPUT83), .B(n572), .Z(n574) );
  NAND2_X1 U634 ( .A1(n663), .A2(G62), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U636 ( .A(KEYINPUT84), .B(n575), .Z(n579) );
  NAND2_X1 U637 ( .A1(G88), .A2(n658), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G75), .A2(n654), .ZN(n576) );
  AND2_X1 U639 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n579), .A2(n578), .ZN(G303) );
  NAND2_X1 U641 ( .A1(n658), .A2(G89), .ZN(n580) );
  XNOR2_X1 U642 ( .A(n580), .B(KEYINPUT4), .ZN(n582) );
  NAND2_X1 U643 ( .A1(G76), .A2(n654), .ZN(n581) );
  NAND2_X1 U644 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U645 ( .A(n583), .B(KEYINPUT5), .ZN(n588) );
  NAND2_X1 U646 ( .A1(G51), .A2(n657), .ZN(n585) );
  NAND2_X1 U647 ( .A1(G63), .A2(n663), .ZN(n584) );
  NAND2_X1 U648 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U649 ( .A(KEYINPUT6), .B(n586), .Z(n587) );
  NAND2_X1 U650 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U651 ( .A(n589), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U652 ( .A(G168), .B(KEYINPUT8), .ZN(n590) );
  XNOR2_X1 U653 ( .A(n590), .B(KEYINPUT75), .ZN(G286) );
  NAND2_X1 U654 ( .A1(G7), .A2(G661), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U656 ( .A(G223), .ZN(n832) );
  NAND2_X1 U657 ( .A1(n832), .A2(G567), .ZN(n592) );
  XOR2_X1 U658 ( .A(KEYINPUT11), .B(n592), .Z(G234) );
  INV_X1 U659 ( .A(G171), .ZN(G301) );
  NAND2_X1 U660 ( .A1(G66), .A2(n663), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G54), .A2(n657), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G92), .A2(n658), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U664 ( .A1(G79), .A2(n654), .ZN(n595) );
  XNOR2_X1 U665 ( .A(KEYINPUT73), .B(n595), .ZN(n596) );
  NOR2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U668 ( .A(n600), .B(KEYINPUT15), .ZN(n601) );
  XNOR2_X1 U669 ( .A(KEYINPUT74), .B(n601), .ZN(n716) );
  INV_X1 U670 ( .A(n716), .ZN(n978) );
  NOR2_X1 U671 ( .A1(n978), .A2(G868), .ZN(n603) );
  INV_X1 U672 ( .A(G868), .ZN(n610) );
  NOR2_X1 U673 ( .A1(n610), .A2(G301), .ZN(n602) );
  NOR2_X1 U674 ( .A1(n603), .A2(n602), .ZN(G284) );
  NAND2_X1 U675 ( .A1(G91), .A2(n658), .ZN(n605) );
  NAND2_X1 U676 ( .A1(G78), .A2(n654), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U678 ( .A1(G53), .A2(n657), .ZN(n607) );
  NAND2_X1 U679 ( .A1(G65), .A2(n663), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n993) );
  INV_X1 U682 ( .A(n993), .ZN(G299) );
  NOR2_X1 U683 ( .A1(G286), .A2(n610), .ZN(n611) );
  XNOR2_X1 U684 ( .A(n611), .B(KEYINPUT76), .ZN(n613) );
  NOR2_X1 U685 ( .A1(G299), .A2(G868), .ZN(n612) );
  NOR2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U687 ( .A(KEYINPUT77), .B(n614), .Z(G297) );
  NAND2_X1 U688 ( .A1(n633), .A2(G559), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n615), .A2(n716), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n616), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U691 ( .A1(n981), .A2(G868), .ZN(n617) );
  XNOR2_X1 U692 ( .A(KEYINPUT78), .B(n617), .ZN(n620) );
  NAND2_X1 U693 ( .A1(G868), .A2(n716), .ZN(n618) );
  NOR2_X1 U694 ( .A1(G559), .A2(n618), .ZN(n619) );
  NOR2_X1 U695 ( .A1(n620), .A2(n619), .ZN(G282) );
  XOR2_X1 U696 ( .A(G2100), .B(KEYINPUT80), .Z(n631) );
  NAND2_X1 U697 ( .A1(G123), .A2(n884), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n621), .B(KEYINPUT18), .ZN(n629) );
  NAND2_X1 U699 ( .A1(G111), .A2(n885), .ZN(n624) );
  BUF_X1 U700 ( .A(n622), .Z(n881) );
  NAND2_X1 U701 ( .A1(G135), .A2(n881), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U703 ( .A1(G99), .A2(n524), .ZN(n625) );
  XNOR2_X1 U704 ( .A(KEYINPUT79), .B(n625), .ZN(n626) );
  NOR2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n927) );
  XOR2_X1 U707 ( .A(G2096), .B(n927), .Z(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(G156) );
  NAND2_X1 U709 ( .A1(n716), .A2(G559), .ZN(n632) );
  XOR2_X1 U710 ( .A(n981), .B(n632), .Z(n671) );
  NAND2_X1 U711 ( .A1(n633), .A2(n671), .ZN(n640) );
  NAND2_X1 U712 ( .A1(G55), .A2(n657), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G67), .A2(n663), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G93), .A2(n658), .ZN(n637) );
  NAND2_X1 U716 ( .A1(G80), .A2(n654), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U718 ( .A1(n639), .A2(n638), .ZN(n673) );
  XOR2_X1 U719 ( .A(n640), .B(n673), .Z(G145) );
  NAND2_X1 U720 ( .A1(G87), .A2(n552), .ZN(n642) );
  NAND2_X1 U721 ( .A1(G74), .A2(G651), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U723 ( .A1(n663), .A2(n643), .ZN(n646) );
  NAND2_X1 U724 ( .A1(G49), .A2(n657), .ZN(n644) );
  XOR2_X1 U725 ( .A(KEYINPUT81), .B(n644), .Z(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(G288) );
  NAND2_X1 U727 ( .A1(G47), .A2(n657), .ZN(n648) );
  NAND2_X1 U728 ( .A1(G60), .A2(n663), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U730 ( .A1(G72), .A2(n654), .ZN(n649) );
  XOR2_X1 U731 ( .A(KEYINPUT70), .B(n649), .Z(n650) );
  NOR2_X1 U732 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U733 ( .A1(n658), .A2(G85), .ZN(n652) );
  NAND2_X1 U734 ( .A1(n653), .A2(n652), .ZN(G290) );
  XOR2_X1 U735 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n656) );
  NAND2_X1 U736 ( .A1(G73), .A2(n654), .ZN(n655) );
  XNOR2_X1 U737 ( .A(n656), .B(n655), .ZN(n662) );
  NAND2_X1 U738 ( .A1(G48), .A2(n657), .ZN(n660) );
  NAND2_X1 U739 ( .A1(G86), .A2(n658), .ZN(n659) );
  NAND2_X1 U740 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U741 ( .A1(n662), .A2(n661), .ZN(n665) );
  NAND2_X1 U742 ( .A1(n663), .A2(G61), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(G305) );
  XNOR2_X1 U744 ( .A(KEYINPUT19), .B(G288), .ZN(n670) );
  XNOR2_X1 U745 ( .A(n993), .B(n673), .ZN(n668) );
  XNOR2_X1 U746 ( .A(G290), .B(G303), .ZN(n666) );
  XNOR2_X1 U747 ( .A(n666), .B(G305), .ZN(n667) );
  XNOR2_X1 U748 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U749 ( .A(n670), .B(n669), .ZN(n907) );
  XNOR2_X1 U750 ( .A(n671), .B(n907), .ZN(n672) );
  NAND2_X1 U751 ( .A1(n672), .A2(G868), .ZN(n675) );
  OR2_X1 U752 ( .A1(G868), .A2(n673), .ZN(n674) );
  NAND2_X1 U753 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U755 ( .A(KEYINPUT20), .B(n676), .Z(n677) );
  NAND2_X1 U756 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U757 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U758 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XOR2_X1 U759 ( .A(KEYINPUT85), .B(G44), .Z(n680) );
  XNOR2_X1 U760 ( .A(KEYINPUT3), .B(n680), .ZN(G218) );
  NOR2_X1 U761 ( .A1(G235), .A2(G236), .ZN(n681) );
  XNOR2_X1 U762 ( .A(n681), .B(KEYINPUT87), .ZN(n682) );
  NOR2_X1 U763 ( .A1(G238), .A2(n682), .ZN(n683) );
  NAND2_X1 U764 ( .A1(G57), .A2(n683), .ZN(n836) );
  NAND2_X1 U765 ( .A1(G567), .A2(n836), .ZN(n689) );
  NAND2_X1 U766 ( .A1(G132), .A2(G82), .ZN(n684) );
  XNOR2_X1 U767 ( .A(n684), .B(KEYINPUT22), .ZN(n685) );
  XNOR2_X1 U768 ( .A(n685), .B(KEYINPUT86), .ZN(n686) );
  NOR2_X1 U769 ( .A1(G218), .A2(n686), .ZN(n687) );
  NAND2_X1 U770 ( .A1(G96), .A2(n687), .ZN(n837) );
  NAND2_X1 U771 ( .A1(G2106), .A2(n837), .ZN(n688) );
  NAND2_X1 U772 ( .A1(n689), .A2(n688), .ZN(n838) );
  NAND2_X1 U773 ( .A1(G483), .A2(G661), .ZN(n690) );
  NOR2_X1 U774 ( .A1(n838), .A2(n690), .ZN(n835) );
  NAND2_X1 U775 ( .A1(n835), .A2(G36), .ZN(G176) );
  NAND2_X1 U776 ( .A1(G40), .A2(G160), .ZN(n783) );
  INV_X1 U777 ( .A(n783), .ZN(n691) );
  NAND2_X1 U778 ( .A1(G8), .A2(n743), .ZN(n779) );
  NOR2_X1 U779 ( .A1(G1981), .A2(G305), .ZN(n692) );
  XOR2_X1 U780 ( .A(n692), .B(KEYINPUT96), .Z(n693) );
  XNOR2_X1 U781 ( .A(KEYINPUT24), .B(n693), .ZN(n694) );
  NOR2_X1 U782 ( .A1(n779), .A2(n694), .ZN(n773) );
  XOR2_X1 U783 ( .A(G1981), .B(KEYINPUT101), .Z(n695) );
  XNOR2_X1 U784 ( .A(G305), .B(n695), .ZN(n983) );
  INV_X1 U785 ( .A(KEYINPUT33), .ZN(n699) );
  NOR2_X1 U786 ( .A1(G1976), .A2(G288), .ZN(n762) );
  INV_X1 U787 ( .A(n762), .ZN(n696) );
  NOR2_X1 U788 ( .A1(KEYINPUT100), .A2(n696), .ZN(n697) );
  NOR2_X1 U789 ( .A1(n779), .A2(n697), .ZN(n698) );
  NOR2_X1 U790 ( .A1(n699), .A2(n698), .ZN(n770) );
  NAND2_X1 U791 ( .A1(n762), .A2(KEYINPUT33), .ZN(n700) );
  NAND2_X1 U792 ( .A1(KEYINPUT100), .A2(n700), .ZN(n768) );
  INV_X1 U793 ( .A(n743), .ZN(n728) );
  NAND2_X1 U794 ( .A1(n728), .A2(G2072), .ZN(n701) );
  XNOR2_X1 U795 ( .A(KEYINPUT27), .B(n701), .ZN(n704) );
  NAND2_X1 U796 ( .A1(G1956), .A2(n743), .ZN(n702) );
  XNOR2_X1 U797 ( .A(KEYINPUT99), .B(n702), .ZN(n703) );
  NOR2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n721) );
  NAND2_X1 U799 ( .A1(n721), .A2(n993), .ZN(n720) );
  INV_X1 U800 ( .A(G1996), .ZN(n953) );
  NOR2_X1 U801 ( .A1(n743), .A2(n953), .ZN(n706) );
  XOR2_X1 U802 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n705) );
  XNOR2_X1 U803 ( .A(n706), .B(n705), .ZN(n708) );
  NAND2_X1 U804 ( .A1(n743), .A2(G1341), .ZN(n707) );
  NAND2_X1 U805 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U806 ( .A1(n709), .A2(n981), .ZN(n710) );
  XNOR2_X1 U807 ( .A(n710), .B(KEYINPUT65), .ZN(n714) );
  AND2_X1 U808 ( .A1(n743), .A2(G1348), .ZN(n712) );
  AND2_X1 U809 ( .A1(n728), .A2(G2067), .ZN(n711) );
  NOR2_X1 U810 ( .A1(n712), .A2(n711), .ZN(n715) );
  NOR2_X1 U811 ( .A1(n716), .A2(n715), .ZN(n713) );
  NOR2_X1 U812 ( .A1(n714), .A2(n713), .ZN(n718) );
  AND2_X1 U813 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U814 ( .A1(n720), .A2(n719), .ZN(n724) );
  NOR2_X1 U815 ( .A1(n721), .A2(n993), .ZN(n722) );
  XOR2_X1 U816 ( .A(n722), .B(KEYINPUT28), .Z(n723) );
  NAND2_X1 U817 ( .A1(n724), .A2(n723), .ZN(n726) );
  XNOR2_X1 U818 ( .A(n726), .B(n725), .ZN(n732) );
  XNOR2_X1 U819 ( .A(G2078), .B(KEYINPUT25), .ZN(n954) );
  NAND2_X1 U820 ( .A1(n728), .A2(n954), .ZN(n727) );
  XNOR2_X1 U821 ( .A(n727), .B(KEYINPUT98), .ZN(n730) );
  OR2_X1 U822 ( .A1(G1961), .A2(n728), .ZN(n729) );
  NAND2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n736) );
  NAND2_X1 U824 ( .A1(n736), .A2(G171), .ZN(n731) );
  NAND2_X1 U825 ( .A1(n732), .A2(n731), .ZN(n741) );
  NOR2_X1 U826 ( .A1(G1966), .A2(n779), .ZN(n755) );
  NOR2_X1 U827 ( .A1(G2084), .A2(n743), .ZN(n753) );
  NOR2_X1 U828 ( .A1(n755), .A2(n753), .ZN(n733) );
  NAND2_X1 U829 ( .A1(G8), .A2(n733), .ZN(n734) );
  XNOR2_X1 U830 ( .A(KEYINPUT30), .B(n734), .ZN(n735) );
  NOR2_X1 U831 ( .A1(G168), .A2(n735), .ZN(n738) );
  NOR2_X1 U832 ( .A1(G171), .A2(n736), .ZN(n737) );
  XOR2_X1 U833 ( .A(KEYINPUT31), .B(n739), .Z(n740) );
  NAND2_X1 U834 ( .A1(n741), .A2(n740), .ZN(n752) );
  AND2_X1 U835 ( .A1(G286), .A2(G8), .ZN(n742) );
  NAND2_X1 U836 ( .A1(n752), .A2(n742), .ZN(n750) );
  INV_X1 U837 ( .A(G8), .ZN(n748) );
  NOR2_X1 U838 ( .A1(G1971), .A2(n779), .ZN(n745) );
  NOR2_X1 U839 ( .A1(G2090), .A2(n743), .ZN(n744) );
  NOR2_X1 U840 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U841 ( .A1(n746), .A2(G303), .ZN(n747) );
  OR2_X1 U842 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U843 ( .A(n751), .B(KEYINPUT32), .ZN(n775) );
  NAND2_X1 U844 ( .A1(G8), .A2(n753), .ZN(n754) );
  XNOR2_X1 U845 ( .A(KEYINPUT97), .B(n754), .ZN(n756) );
  NOR2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U847 ( .A1(n752), .A2(n757), .ZN(n774) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n988) );
  INV_X1 U849 ( .A(n779), .ZN(n758) );
  NAND2_X1 U850 ( .A1(n988), .A2(n758), .ZN(n763) );
  INV_X1 U851 ( .A(n763), .ZN(n759) );
  AND2_X1 U852 ( .A1(n774), .A2(n759), .ZN(n760) );
  NAND2_X1 U853 ( .A1(n775), .A2(n760), .ZN(n766) );
  NOR2_X1 U854 ( .A1(G1971), .A2(G303), .ZN(n761) );
  NOR2_X1 U855 ( .A1(n762), .A2(n761), .ZN(n989) );
  NOR2_X1 U856 ( .A1(n763), .A2(n989), .ZN(n764) );
  NOR2_X1 U857 ( .A1(n764), .A2(KEYINPUT33), .ZN(n765) );
  AND2_X1 U858 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U859 ( .A1(n775), .A2(n774), .ZN(n778) );
  NOR2_X1 U860 ( .A1(G2090), .A2(G303), .ZN(n776) );
  NAND2_X1 U861 ( .A1(G8), .A2(n776), .ZN(n777) );
  NAND2_X1 U862 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U863 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U864 ( .A1(n782), .A2(n781), .ZN(n796) );
  NOR2_X1 U865 ( .A1(n784), .A2(n783), .ZN(n826) );
  NAND2_X1 U866 ( .A1(n524), .A2(G104), .ZN(n785) );
  XOR2_X1 U867 ( .A(KEYINPUT91), .B(n785), .Z(n787) );
  NAND2_X1 U868 ( .A1(G140), .A2(n881), .ZN(n786) );
  NAND2_X1 U869 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U870 ( .A(KEYINPUT34), .B(n788), .ZN(n793) );
  NAND2_X1 U871 ( .A1(G128), .A2(n884), .ZN(n790) );
  NAND2_X1 U872 ( .A1(G116), .A2(n885), .ZN(n789) );
  NAND2_X1 U873 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U874 ( .A(n791), .B(KEYINPUT35), .Z(n792) );
  NOR2_X1 U875 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U876 ( .A(KEYINPUT36), .B(n794), .Z(n795) );
  XOR2_X1 U877 ( .A(KEYINPUT92), .B(n795), .Z(n901) );
  XNOR2_X1 U878 ( .A(G2067), .B(KEYINPUT37), .ZN(n824) );
  NOR2_X1 U879 ( .A1(n901), .A2(n824), .ZN(n945) );
  NAND2_X1 U880 ( .A1(n826), .A2(n945), .ZN(n822) );
  NAND2_X1 U881 ( .A1(n524), .A2(G95), .ZN(n798) );
  NAND2_X1 U882 ( .A1(G131), .A2(n881), .ZN(n797) );
  NAND2_X1 U883 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U884 ( .A(KEYINPUT93), .B(n799), .ZN(n803) );
  NAND2_X1 U885 ( .A1(G119), .A2(n884), .ZN(n801) );
  NAND2_X1 U886 ( .A1(G107), .A2(n885), .ZN(n800) );
  AND2_X1 U887 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U888 ( .A1(n803), .A2(n802), .ZN(n896) );
  AND2_X1 U889 ( .A1(n896), .A2(G1991), .ZN(n813) );
  XOR2_X1 U890 ( .A(KEYINPUT94), .B(KEYINPUT38), .Z(n805) );
  NAND2_X1 U891 ( .A1(G105), .A2(n524), .ZN(n804) );
  XNOR2_X1 U892 ( .A(n805), .B(n804), .ZN(n809) );
  NAND2_X1 U893 ( .A1(G117), .A2(n885), .ZN(n807) );
  NAND2_X1 U894 ( .A1(G141), .A2(n881), .ZN(n806) );
  NAND2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U896 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U897 ( .A1(n884), .A2(G129), .ZN(n810) );
  NAND2_X1 U898 ( .A1(n811), .A2(n810), .ZN(n891) );
  AND2_X1 U899 ( .A1(n891), .A2(G1996), .ZN(n812) );
  NOR2_X1 U900 ( .A1(n813), .A2(n812), .ZN(n932) );
  INV_X1 U901 ( .A(n826), .ZN(n814) );
  NOR2_X1 U902 ( .A1(n932), .A2(n814), .ZN(n819) );
  XOR2_X1 U903 ( .A(KEYINPUT95), .B(n819), .Z(n815) );
  XNOR2_X1 U904 ( .A(G1986), .B(G290), .ZN(n997) );
  NAND2_X1 U905 ( .A1(n529), .A2(n525), .ZN(n829) );
  NOR2_X1 U906 ( .A1(n891), .A2(G1996), .ZN(n816) );
  XNOR2_X1 U907 ( .A(n816), .B(KEYINPUT102), .ZN(n938) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U909 ( .A1(G1991), .A2(n896), .ZN(n930) );
  NOR2_X1 U910 ( .A1(n817), .A2(n930), .ZN(n818) );
  NOR2_X1 U911 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U912 ( .A1(n938), .A2(n820), .ZN(n821) );
  XNOR2_X1 U913 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U914 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n901), .A2(n824), .ZN(n944) );
  NAND2_X1 U916 ( .A1(n825), .A2(n944), .ZN(n827) );
  NAND2_X1 U917 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U918 ( .A1(n829), .A2(n828), .ZN(n831) );
  XOR2_X1 U919 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n830) );
  XNOR2_X1 U920 ( .A(n831), .B(n830), .ZN(G329) );
  INV_X1 U921 ( .A(G303), .ZN(G166) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U924 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U926 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U928 ( .A(G132), .ZN(G219) );
  INV_X1 U929 ( .A(G82), .ZN(G220) );
  NOR2_X1 U930 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  XOR2_X1 U932 ( .A(KEYINPUT104), .B(n838), .Z(G319) );
  XOR2_X1 U933 ( .A(G1981), .B(G1956), .Z(n840) );
  XNOR2_X1 U934 ( .A(G1986), .B(G1966), .ZN(n839) );
  XNOR2_X1 U935 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U936 ( .A(G1976), .B(G1971), .Z(n842) );
  XNOR2_X1 U937 ( .A(G1996), .B(G1991), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U939 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U940 ( .A(KEYINPUT107), .B(G2474), .ZN(n845) );
  XNOR2_X1 U941 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U942 ( .A(KEYINPUT41), .B(n847), .ZN(n848) );
  XOR2_X1 U943 ( .A(n848), .B(G1961), .Z(G229) );
  XOR2_X1 U944 ( .A(KEYINPUT106), .B(G2678), .Z(n850) );
  XNOR2_X1 U945 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U947 ( .A(KEYINPUT42), .B(G2090), .Z(n852) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U950 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U951 ( .A(G2100), .B(G2096), .ZN(n855) );
  XNOR2_X1 U952 ( .A(n856), .B(n855), .ZN(n858) );
  XOR2_X1 U953 ( .A(G2078), .B(G2084), .Z(n857) );
  XNOR2_X1 U954 ( .A(n858), .B(n857), .ZN(G227) );
  NAND2_X1 U955 ( .A1(G112), .A2(n885), .ZN(n860) );
  NAND2_X1 U956 ( .A1(G100), .A2(n524), .ZN(n859) );
  NAND2_X1 U957 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U958 ( .A(KEYINPUT108), .B(n861), .ZN(n864) );
  NAND2_X1 U959 ( .A1(n884), .A2(G124), .ZN(n862) );
  XOR2_X1 U960 ( .A(KEYINPUT44), .B(n862), .Z(n863) );
  NOR2_X1 U961 ( .A1(n864), .A2(n863), .ZN(n866) );
  NAND2_X1 U962 ( .A1(G136), .A2(n881), .ZN(n865) );
  NAND2_X1 U963 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U964 ( .A(KEYINPUT109), .B(n867), .ZN(G162) );
  NAND2_X1 U965 ( .A1(G142), .A2(n881), .ZN(n868) );
  XOR2_X1 U966 ( .A(KEYINPUT111), .B(n868), .Z(n870) );
  NAND2_X1 U967 ( .A1(n524), .A2(G106), .ZN(n869) );
  NAND2_X1 U968 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U969 ( .A(n871), .B(KEYINPUT45), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G118), .A2(n885), .ZN(n872) );
  NAND2_X1 U971 ( .A1(n873), .A2(n872), .ZN(n876) );
  NAND2_X1 U972 ( .A1(n884), .A2(G130), .ZN(n874) );
  XOR2_X1 U973 ( .A(KEYINPUT110), .B(n874), .Z(n875) );
  NOR2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n895) );
  XOR2_X1 U975 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n878) );
  XNOR2_X1 U976 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U978 ( .A(n927), .B(n879), .ZN(n893) );
  NAND2_X1 U979 ( .A1(n524), .A2(G103), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G139), .A2(n881), .ZN(n882) );
  NAND2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n890) );
  NAND2_X1 U982 ( .A1(G127), .A2(n884), .ZN(n887) );
  NAND2_X1 U983 ( .A1(G115), .A2(n885), .ZN(n886) );
  NAND2_X1 U984 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U985 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U986 ( .A1(n890), .A2(n889), .ZN(n933) );
  XOR2_X1 U987 ( .A(n891), .B(n933), .Z(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n898) );
  XOR2_X1 U990 ( .A(G160), .B(n896), .Z(n897) );
  XNOR2_X1 U991 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U992 ( .A(G162), .B(n899), .Z(n900) );
  XNOR2_X1 U993 ( .A(G164), .B(n900), .ZN(n902) );
  XNOR2_X1 U994 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U995 ( .A1(G37), .A2(n903), .ZN(n904) );
  XNOR2_X1 U996 ( .A(KEYINPUT114), .B(n904), .ZN(G395) );
  XOR2_X1 U997 ( .A(KEYINPUT115), .B(n981), .Z(n906) );
  XNOR2_X1 U998 ( .A(G171), .B(n978), .ZN(n905) );
  XNOR2_X1 U999 ( .A(n906), .B(n905), .ZN(n909) );
  XOR2_X1 U1000 ( .A(G286), .B(n907), .Z(n908) );
  XNOR2_X1 U1001 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n910), .ZN(n911) );
  XNOR2_X1 U1003 ( .A(KEYINPUT116), .B(n911), .ZN(G397) );
  XOR2_X1 U1004 ( .A(G2451), .B(G2430), .Z(n913) );
  XNOR2_X1 U1005 ( .A(G2438), .B(G2443), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n913), .B(n912), .ZN(n919) );
  XOR2_X1 U1007 ( .A(G2435), .B(G2454), .Z(n915) );
  XNOR2_X1 U1008 ( .A(G1348), .B(G1341), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n917) );
  XOR2_X1 U1010 ( .A(G2446), .B(G2427), .Z(n916) );
  XNOR2_X1 U1011 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1012 ( .A(n919), .B(n918), .Z(n920) );
  NAND2_X1 U1013 ( .A1(G14), .A2(n920), .ZN(n926) );
  NAND2_X1 U1014 ( .A1(n926), .A2(G319), .ZN(n923) );
  NOR2_X1 U1015 ( .A1(G229), .A2(G227), .ZN(n921) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(n921), .ZN(n922) );
  NOR2_X1 U1017 ( .A1(n923), .A2(n922), .ZN(n925) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n924) );
  NAND2_X1 U1019 ( .A1(n925), .A2(n924), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(G96), .ZN(G221) );
  INV_X1 U1022 ( .A(G57), .ZN(G237) );
  INV_X1 U1023 ( .A(n926), .ZN(G401) );
  XNOR2_X1 U1024 ( .A(G160), .B(G2084), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n943) );
  XOR2_X1 U1028 ( .A(G2072), .B(n933), .Z(n935) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(KEYINPUT50), .B(n936), .ZN(n941) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1034 ( .A(KEYINPUT51), .B(n939), .Z(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n948) );
  INV_X1 U1037 ( .A(n944), .ZN(n946) );
  NOR2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1039 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1040 ( .A(KEYINPUT117), .B(n949), .ZN(n950) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n950), .ZN(n951) );
  XOR2_X1 U1042 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n974) );
  NAND2_X1 U1043 ( .A1(n951), .A2(n974), .ZN(n952) );
  NAND2_X1 U1044 ( .A1(n952), .A2(G29), .ZN(n1034) );
  XNOR2_X1 U1045 ( .A(G2090), .B(G35), .ZN(n969) );
  XNOR2_X1 U1046 ( .A(G32), .B(n953), .ZN(n961) );
  XOR2_X1 U1047 ( .A(n954), .B(G27), .Z(n959) );
  XNOR2_X1 U1048 ( .A(G2067), .B(G26), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(G2072), .B(G33), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(KEYINPUT121), .B(n957), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n966) );
  XNOR2_X1 U1054 ( .A(G1991), .B(G25), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n962), .B(KEYINPUT119), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(G28), .A2(n963), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(KEYINPUT120), .B(n964), .ZN(n965) );
  NOR2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(KEYINPUT53), .B(n967), .ZN(n968) );
  NOR2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n972) );
  XOR2_X1 U1061 ( .A(G2084), .B(KEYINPUT54), .Z(n970) );
  XNOR2_X1 U1062 ( .A(G34), .B(n970), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(n974), .B(n973), .ZN(n976) );
  INV_X1 U1065 ( .A(G29), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1067 ( .A1(G11), .A2(n977), .ZN(n1032) );
  XNOR2_X1 U1068 ( .A(G16), .B(KEYINPUT56), .ZN(n1004) );
  XNOR2_X1 U1069 ( .A(G301), .B(G1961), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(n978), .B(G1348), .ZN(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n1002) );
  XOR2_X1 U1072 ( .A(n981), .B(G1341), .Z(n987) );
  XOR2_X1 U1073 ( .A(G168), .B(G1966), .Z(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1075 ( .A(KEYINPUT57), .B(n984), .Z(n985) );
  XNOR2_X1 U1076 ( .A(KEYINPUT122), .B(n985), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n1000) );
  AND2_X1 U1078 ( .A1(G303), .A2(G1971), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1081 ( .A(KEYINPUT123), .B(n992), .Z(n995) );
  XNOR2_X1 U1082 ( .A(n993), .B(G1956), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1085 ( .A(KEYINPUT124), .B(n998), .Z(n999) );
  NOR2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1087 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1088 ( .A1(n1004), .A2(n1003), .ZN(n1030) );
  INV_X1 U1089 ( .A(G16), .ZN(n1028) );
  XOR2_X1 U1090 ( .A(G5), .B(G1961), .Z(n1023) );
  XNOR2_X1 U1091 ( .A(KEYINPUT126), .B(KEYINPUT60), .ZN(n1014) );
  XNOR2_X1 U1092 ( .A(KEYINPUT59), .B(G1348), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(n1005), .B(G4), .ZN(n1012) );
  XNOR2_X1 U1094 ( .A(G1956), .B(G20), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(G1341), .B(G19), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(G1981), .B(G6), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(KEYINPUT125), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(n1014), .B(n1013), .ZN(n1021) );
  XNOR2_X1 U1102 ( .A(G1971), .B(G22), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(G23), .B(G1976), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XOR2_X1 U1105 ( .A(G1986), .B(G24), .Z(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(KEYINPUT58), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1025) );
  XNOR2_X1 U1110 ( .A(G21), .B(G1966), .ZN(n1024) );
  NOR2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1112 ( .A(KEYINPUT61), .B(n1026), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1115 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1116 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1117 ( .A(n1035), .B(KEYINPUT62), .ZN(n1036) );
  XNOR2_X1 U1118 ( .A(KEYINPUT127), .B(n1036), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

