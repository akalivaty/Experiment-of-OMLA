//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT31), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT66), .A2(G146), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT66), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NOR3_X1   g005(.A1(new_n189), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n193));
  OAI21_X1  g007(.A(G128), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n189), .B2(new_n190), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n196), .B1(new_n191), .B2(G146), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT65), .A3(G143), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n198), .A2(G143), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n189), .A2(new_n190), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n194), .A2(new_n200), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT67), .B1(new_n207), .B2(G134), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G137), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT11), .B1(new_n210), .B2(G137), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT11), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n207), .A3(G134), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n212), .A2(new_n213), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n207), .A2(G134), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n210), .A2(G137), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n219), .B1(new_n222), .B2(new_n213), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n213), .B1(new_n220), .B2(new_n221), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT68), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n218), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT71), .B1(new_n206), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n198), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT66), .A2(G146), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(G143), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n201), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(new_n205), .ZN(new_n233));
  AOI21_X1  g047(.A(G143), .B1(new_n229), .B2(new_n230), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n197), .A2(new_n199), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n204), .B1(new_n231), .B2(KEYINPUT1), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n233), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT71), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n224), .B(new_n219), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n238), .A2(new_n239), .A3(new_n218), .A4(new_n240), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n231), .A2(KEYINPUT0), .A3(G128), .A4(new_n232), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT0), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n204), .A3(KEYINPUT64), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n245), .B1(KEYINPUT0), .B2(G128), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n244), .A2(new_n246), .B1(KEYINPUT0), .B2(G128), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n234), .B2(new_n235), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n212), .A2(new_n213), .A3(new_n217), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n213), .B1(new_n212), .B2(new_n217), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n242), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n227), .A2(new_n241), .A3(KEYINPUT30), .A4(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n249), .A2(new_n250), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n248), .A2(new_n242), .ZN(new_n254));
  OAI22_X1  g068(.A1(new_n253), .A2(new_n254), .B1(new_n206), .B2(new_n226), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(KEYINPUT2), .A2(G113), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT2), .ZN(new_n260));
  INV_X1    g074(.A(G113), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT69), .B1(KEYINPUT2), .B2(G113), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n258), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G119), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G116), .ZN(new_n266));
  INV_X1    g080(.A(G116), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G119), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT70), .B1(new_n264), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n263), .ZN(new_n272));
  NOR3_X1   g086(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n273));
  OAI22_X1  g087(.A1(new_n272), .A2(new_n273), .B1(new_n260), .B2(new_n261), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n269), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n274), .A2(KEYINPUT70), .A3(new_n269), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n252), .A2(new_n257), .A3(new_n279), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n227), .A2(new_n241), .A3(new_n278), .A4(new_n251), .ZN(new_n281));
  NOR2_X1   g095(.A1(G237), .A2(G953), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G210), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(KEYINPUT27), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(G101), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n284), .B(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n188), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n287), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n278), .B1(new_n255), .B2(new_n256), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n252), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n291), .A3(KEYINPUT31), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n238), .A2(new_n218), .A3(new_n240), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n278), .A3(new_n251), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT28), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n294), .A2(KEYINPUT72), .A3(new_n295), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n255), .A2(new_n279), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n281), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n298), .B(new_n299), .C1(new_n301), .C2(new_n295), .ZN(new_n302));
  INV_X1    g116(.A(new_n286), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n288), .A2(new_n292), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G472), .A2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n187), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n288), .A2(new_n292), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n298), .A2(new_n299), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n295), .B1(new_n281), .B2(new_n300), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n303), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n306), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT32), .ZN(new_n313));
  INV_X1    g127(.A(G902), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n227), .A2(new_n241), .A3(new_n251), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n279), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n281), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT28), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n294), .A2(KEYINPUT72), .A3(new_n295), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT72), .B1(new_n294), .B2(new_n295), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n303), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n318), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n315), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n278), .A2(new_n325), .B1(new_n290), .B2(new_n252), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n322), .B1(new_n326), .B2(new_n286), .ZN(new_n327));
  NOR4_X1   g141(.A1(new_n310), .A2(new_n319), .A3(new_n320), .A4(new_n303), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n314), .B(new_n324), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G472), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n307), .A2(new_n313), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT74), .B1(new_n265), .B2(G128), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT23), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n334));
  OAI211_X1 g148(.A(KEYINPUT74), .B(new_n334), .C1(new_n265), .C2(G128), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n265), .A2(G128), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT78), .B(G110), .ZN(new_n338));
  XNOR2_X1  g152(.A(G119), .B(G128), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT24), .B(G110), .Z(new_n340));
  OAI22_X1  g154(.A1(new_n337), .A2(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(G125), .B(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n202), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT79), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n202), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G140), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G125), .ZN(new_n349));
  INV_X1    g163(.A(G125), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G140), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n351), .A3(KEYINPUT16), .ZN(new_n352));
  OR3_X1    g166(.A1(new_n350), .A2(KEYINPUT16), .A3(G140), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(G146), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n341), .A2(new_n347), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G110), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n337), .B2(KEYINPUT75), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT75), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n333), .A2(new_n359), .A3(new_n335), .A4(new_n336), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n354), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(G146), .B1(new_n352), .B2(new_n353), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT76), .A4(G146), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n340), .A2(new_n339), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n361), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT77), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n361), .A2(new_n367), .A3(KEYINPUT77), .A4(new_n368), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n356), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT22), .B(G137), .ZN(new_n374));
  INV_X1    g188(.A(G221), .ZN(new_n375));
  INV_X1    g189(.A(G234), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n375), .A2(new_n376), .A3(G953), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n374), .B(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n373), .A2(new_n379), .ZN(new_n380));
  AOI211_X1 g194(.A(new_n356), .B(new_n378), .C1(new_n371), .C2(new_n372), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G217), .B1(new_n376), .B2(G902), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT73), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G902), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n371), .A2(new_n372), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n355), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n378), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n373), .A2(new_n379), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n314), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT25), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n382), .A2(KEYINPUT25), .A3(new_n314), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n388), .B1(new_n397), .B2(new_n385), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n331), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT9), .B(G234), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n375), .B1(new_n401), .B2(new_n314), .ZN(new_n402));
  INV_X1    g216(.A(G469), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(new_n314), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT80), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(KEYINPUT3), .ZN(new_n406));
  INV_X1    g220(.A(G104), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(G107), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(KEYINPUT3), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(G107), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT3), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT80), .ZN(new_n413));
  INV_X1    g227(.A(G107), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G104), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n411), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G101), .B1(new_n410), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n412), .A2(KEYINPUT80), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n413), .B1(new_n418), .B2(new_n415), .ZN(new_n419));
  INV_X1    g233(.A(G101), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n406), .A2(new_n408), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n419), .A2(new_n420), .A3(new_n411), .A4(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n417), .A2(KEYINPUT4), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT4), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n424), .B(G101), .C1(new_n410), .C2(new_n416), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n423), .A2(new_n242), .A3(new_n248), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n415), .A2(new_n411), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G101), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n238), .A3(KEYINPUT10), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n231), .A2(new_n232), .A3(new_n205), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n231), .A2(new_n232), .B1(G128), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n422), .B(new_n428), .C1(new_n431), .C2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT10), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n426), .A2(new_n430), .A3(new_n436), .A4(new_n253), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G140), .ZN(new_n438));
  INV_X1    g252(.A(G953), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n439), .A2(G227), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n438), .B(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n253), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n426), .A2(new_n430), .A3(new_n436), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT81), .B1(new_n429), .B2(new_n238), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT81), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n422), .A2(new_n428), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n206), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(new_n434), .A3(new_n450), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n451), .A2(KEYINPUT12), .A3(new_n444), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT12), .B1(new_n451), .B2(new_n444), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n437), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n446), .B1(new_n454), .B2(new_n441), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n404), .B1(new_n455), .B2(G469), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n451), .A2(new_n444), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT12), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n451), .A2(KEYINPUT12), .A3(new_n444), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n443), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n445), .A2(new_n444), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n442), .B1(new_n462), .B2(new_n437), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n403), .B(new_n314), .C1(new_n461), .C2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n402), .B1(new_n456), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G214), .B1(G237), .B2(G902), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n423), .A2(new_n276), .A3(new_n277), .A4(new_n425), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n264), .A2(new_n270), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT5), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n265), .A3(G116), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n471), .B(G113), .C1(new_n269), .C2(new_n470), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n429), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(G110), .B(G122), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n468), .A2(new_n473), .A3(new_n475), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(KEYINPUT6), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n474), .A2(new_n480), .A3(new_n476), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n238), .A2(new_n350), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n248), .A2(G125), .A3(new_n242), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G224), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(G953), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n484), .B(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n479), .A2(new_n481), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(KEYINPUT7), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n193), .B1(new_n202), .B2(G143), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n200), .B1(new_n492), .B2(new_n204), .ZN(new_n493));
  AOI21_X1  g307(.A(G125), .B1(new_n493), .B2(new_n233), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n248), .A2(G125), .A3(new_n242), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n475), .B(KEYINPUT8), .ZN(new_n497));
  AND4_X1   g311(.A1(new_n469), .A2(new_n422), .A3(new_n428), .A4(new_n472), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n422), .A2(new_n428), .B1(new_n469), .B2(new_n472), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n482), .A2(new_n483), .A3(new_n490), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n496), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT82), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n496), .A2(new_n500), .A3(new_n501), .A4(KEYINPUT82), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n478), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n489), .A2(new_n506), .A3(new_n314), .ZN(new_n507));
  OAI21_X1  g321(.A(G210), .B1(G237), .B2(G902), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n489), .A2(new_n506), .A3(new_n314), .A4(new_n508), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n467), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(G475), .A2(G902), .ZN(new_n513));
  INV_X1    g327(.A(G237), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n439), .A3(G214), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT83), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n515), .B1(new_n516), .B2(new_n191), .ZN(new_n517));
  AND2_X1   g331(.A1(KEYINPUT83), .A2(G143), .ZN(new_n518));
  NOR2_X1   g332(.A1(KEYINPUT83), .A2(G143), .ZN(new_n519));
  OAI211_X1 g333(.A(G214), .B(new_n282), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G131), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n517), .A2(new_n520), .A3(new_n213), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n364), .B1(new_n362), .B2(new_n354), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n213), .B1(new_n517), .B2(new_n520), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT17), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n525), .A2(new_n366), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n342), .A2(new_n198), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n347), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT18), .ZN(new_n533));
  AOI211_X1 g347(.A(new_n533), .B(new_n213), .C1(new_n517), .C2(new_n520), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n533), .A2(new_n213), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n521), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n532), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(G113), .B(G122), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n540), .A2(KEYINPUT85), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(KEYINPUT85), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT84), .B(G104), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n543), .B1(new_n541), .B2(new_n542), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n529), .A2(new_n539), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n524), .ZN(new_n548));
  XOR2_X1   g362(.A(new_n342), .B(KEYINPUT19), .Z(new_n549));
  INV_X1    g363(.A(new_n202), .ZN(new_n550));
  OAI221_X1 g364(.A(new_n354), .B1(new_n548), .B2(new_n527), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n546), .B1(new_n551), .B2(new_n539), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n513), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT20), .ZN(new_n554));
  INV_X1    g368(.A(new_n546), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n354), .B1(new_n549), .B2(new_n550), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n548), .A2(new_n527), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n530), .B1(new_n344), .B2(new_n346), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n559), .A2(new_n534), .A3(new_n537), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n555), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n529), .A2(new_n539), .A3(new_n546), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT20), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n513), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n554), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G478), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(KEYINPUT15), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n191), .A2(G128), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n204), .A2(G143), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n569), .A2(new_n570), .A3(new_n210), .ZN(new_n571));
  XOR2_X1   g385(.A(G116), .B(G122), .Z(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G107), .ZN(new_n573));
  XNOR2_X1  g387(.A(G116), .B(G122), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n414), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n571), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT13), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n569), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n570), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n569), .A2(new_n577), .ZN(new_n580));
  OAI21_X1  g394(.A(G134), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n267), .A2(KEYINPUT14), .A3(G122), .ZN(new_n583));
  OAI211_X1 g397(.A(G107), .B(new_n583), .C1(new_n572), .C2(KEYINPUT14), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n210), .B1(new_n569), .B2(new_n570), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n584), .B(new_n575), .C1(new_n571), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n401), .A2(G217), .A3(new_n439), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n588), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n582), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n314), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT88), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n568), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  AOI21_X1  g410(.A(G902), .B1(new_n589), .B2(new_n591), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT88), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n595), .B1(new_n599), .B2(new_n568), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT86), .B(G475), .Z(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n529), .A2(new_n539), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n555), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT87), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT87), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n603), .A2(new_n606), .A3(new_n555), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n547), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n602), .B1(new_n608), .B2(G902), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n439), .A2(G952), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n376), .B2(new_n514), .ZN(new_n611));
  AOI211_X1 g425(.A(new_n314), .B(new_n439), .C1(G234), .C2(G237), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT21), .B(G898), .Z(new_n614));
  OAI21_X1  g428(.A(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AND4_X1   g429(.A1(new_n566), .A2(new_n600), .A3(new_n609), .A4(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n465), .A2(new_n512), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n399), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT89), .B(G101), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G3));
  NOR3_X1   g434(.A1(new_n280), .A2(new_n188), .A3(new_n287), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT31), .B1(new_n289), .B2(new_n291), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n311), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(KEYINPUT90), .A2(G472), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n314), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n624), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n626), .B1(new_n304), .B2(G902), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n465), .A2(new_n398), .A3(new_n625), .A4(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n512), .A2(new_n615), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n609), .A2(new_n566), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n588), .B2(KEYINPUT91), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n589), .B2(new_n591), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n589), .A2(new_n591), .A3(new_n633), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n567), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n567), .A2(new_n314), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n593), .B2(G478), .ZN(new_n640));
  OAI21_X1  g454(.A(KEYINPUT92), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n636), .ZN(new_n642));
  OAI21_X1  g456(.A(G478), .B1(new_n642), .B2(new_n634), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT92), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n638), .B1(new_n597), .B2(new_n567), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n631), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n630), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n629), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  AOI21_X1  g466(.A(new_n606), .B1(new_n603), .B2(new_n555), .ZN(new_n653));
  AOI211_X1 g467(.A(KEYINPUT87), .B(new_n546), .C1(new_n529), .C2(new_n539), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n562), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AOI211_X1 g469(.A(KEYINPUT94), .B(new_n601), .C1(new_n655), .C2(new_n314), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n554), .A2(KEYINPUT93), .A3(new_n565), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT93), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n553), .A2(new_n659), .A3(KEYINPUT20), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n599), .A2(new_n568), .ZN(new_n662));
  INV_X1    g476(.A(new_n595), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n609), .A2(KEYINPUT94), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n657), .A2(new_n661), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n630), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n629), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT35), .B(G107), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  NAND2_X1  g484(.A1(new_n627), .A2(new_n625), .ZN(new_n671));
  AOI211_X1 g485(.A(KEYINPUT95), .B(new_n356), .C1(new_n371), .C2(new_n372), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n390), .A2(KEYINPUT95), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n378), .A2(KEYINPUT36), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT95), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n373), .A2(new_n677), .ZN(new_n678));
  OAI22_X1  g492(.A1(new_n678), .A2(new_n672), .B1(KEYINPUT36), .B2(new_n378), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n387), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n397), .B2(new_n385), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT96), .B1(new_n671), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT25), .B1(new_n382), .B2(new_n314), .ZN(new_n683));
  NOR4_X1   g497(.A1(new_n380), .A2(new_n381), .A3(new_n394), .A4(G902), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n385), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n680), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT96), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n687), .A2(new_n688), .A3(new_n625), .A4(new_n627), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n617), .B1(new_n682), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT37), .B(G110), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G12));
  INV_X1    g506(.A(new_n402), .ZN(new_n693));
  INV_X1    g507(.A(new_n443), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n462), .ZN(new_n695));
  INV_X1    g509(.A(new_n437), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n459), .B2(new_n460), .ZN(new_n697));
  OAI211_X1 g511(.A(G469), .B(new_n695), .C1(new_n697), .C2(new_n442), .ZN(new_n698));
  INV_X1    g512(.A(new_n404), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n464), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n512), .A2(new_n693), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n601), .B1(new_n655), .B2(new_n314), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT94), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n660), .B(new_n658), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(G900), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n612), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n611), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NOR4_X1   g522(.A1(new_n704), .A2(new_n600), .A3(new_n656), .A4(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n701), .A2(new_n709), .A3(new_n331), .A4(new_n687), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G128), .ZN(G30));
  XNOR2_X1  g525(.A(new_n707), .B(KEYINPUT39), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n465), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n713), .B(KEYINPUT40), .Z(new_n714));
  OR2_X1    g528(.A1(new_n714), .A2(KEYINPUT98), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(KEYINPUT98), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n510), .A2(new_n511), .ZN(new_n717));
  XOR2_X1   g531(.A(new_n717), .B(KEYINPUT38), .Z(new_n718));
  OAI21_X1  g532(.A(new_n314), .B1(new_n317), .B2(new_n286), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n303), .B1(new_n291), .B2(new_n281), .ZN(new_n720));
  OAI21_X1  g534(.A(G472), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT97), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n307), .A3(new_n313), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n600), .B1(new_n609), .B2(new_n566), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n466), .ZN(new_n727));
  NOR4_X1   g541(.A1(new_n718), .A2(new_n725), .A3(new_n687), .A4(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n715), .A2(new_n716), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G143), .ZN(G45));
  NAND3_X1  g544(.A1(new_n631), .A2(new_n647), .A3(new_n707), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n701), .A2(new_n331), .A3(new_n687), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G146), .ZN(G48));
  NAND2_X1  g548(.A1(new_n459), .A2(new_n460), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n463), .B1(new_n735), .B2(new_n694), .ZN(new_n736));
  OAI21_X1  g550(.A(G469), .B1(new_n736), .B2(G902), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n693), .A3(new_n464), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT99), .ZN(new_n739));
  INV_X1    g553(.A(new_n388), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n685), .A2(new_n740), .ZN(new_n741));
  AOI211_X1 g555(.A(new_n187), .B(new_n306), .C1(new_n308), .C2(new_n311), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT32), .B1(new_n623), .B2(new_n305), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n741), .B1(new_n744), .B2(new_n330), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(new_n649), .ZN(new_n747));
  XOR2_X1   g561(.A(KEYINPUT41), .B(G113), .Z(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G15));
  AND2_X1   g563(.A1(new_n746), .A2(new_n667), .ZN(new_n750));
  XOR2_X1   g564(.A(KEYINPUT100), .B(G116), .Z(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(G18));
  AOI21_X1  g566(.A(new_n681), .B1(new_n744), .B2(new_n330), .ZN(new_n753));
  INV_X1    g567(.A(new_n464), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n694), .B1(new_n452), .B2(new_n453), .ZN(new_n755));
  INV_X1    g569(.A(new_n463), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n403), .B1(new_n757), .B2(new_n314), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n616), .A2(new_n759), .A3(new_n512), .A4(new_n693), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT101), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n753), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n331), .A2(new_n687), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT101), .B1(new_n764), .B2(new_n760), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G119), .ZN(G21));
  AOI21_X1  g581(.A(new_n295), .B1(new_n316), .B2(new_n281), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT102), .B1(new_n309), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n303), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n309), .A2(new_n768), .A3(KEYINPUT102), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n308), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n623), .A2(new_n314), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n772), .A2(new_n305), .B1(new_n773), .B2(G472), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(new_n398), .ZN(new_n775));
  INV_X1    g589(.A(new_n726), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n630), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n739), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G122), .ZN(G24));
  NAND2_X1  g593(.A1(new_n717), .A2(new_n466), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n738), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n781), .A2(new_n774), .A3(new_n687), .A4(new_n732), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G125), .ZN(G27));
  NAND2_X1  g597(.A1(new_n700), .A2(KEYINPUT103), .ZN(new_n784));
  AND4_X1   g598(.A1(new_n466), .A2(new_n510), .A3(new_n511), .A4(new_n693), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT103), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n456), .A2(new_n786), .A3(new_n464), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT104), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT104), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n784), .A2(new_n785), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT105), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(new_n312), .B2(KEYINPUT32), .ZN(new_n794));
  OAI211_X1 g608(.A(KEYINPUT105), .B(new_n187), .C1(new_n304), .C2(new_n306), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n794), .A2(new_n795), .A3(new_n313), .A4(new_n330), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT42), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n731), .A2(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n796), .A2(new_n398), .A3(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n792), .A2(KEYINPUT106), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT106), .B1(new_n792), .B2(new_n799), .ZN(new_n801));
  AOI211_X1 g615(.A(new_n731), .B(new_n399), .C1(new_n789), .C2(new_n791), .ZN(new_n802));
  OAI22_X1  g616(.A1(new_n800), .A2(new_n801), .B1(new_n802), .B2(KEYINPUT42), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G131), .ZN(G33));
  NAND3_X1  g618(.A1(new_n792), .A2(new_n745), .A3(new_n709), .ZN(new_n805));
  XOR2_X1   g619(.A(KEYINPUT107), .B(G134), .Z(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(G36));
  NAND3_X1  g621(.A1(new_n647), .A2(new_n566), .A3(new_n609), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT43), .ZN(new_n809));
  INV_X1    g623(.A(new_n671), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n809), .A2(new_n810), .A3(new_n681), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(KEYINPUT44), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(KEYINPUT44), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n717), .A2(new_n467), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT109), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT109), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n813), .A2(new_n817), .A3(new_n814), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n812), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(G469), .B1(new_n455), .B2(KEYINPUT45), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT45), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n821), .B(new_n446), .C1(new_n454), .C2(new_n441), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT108), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n823), .B1(new_n820), .B2(new_n822), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n699), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT46), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n826), .A2(KEYINPUT46), .A3(new_n699), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n464), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n693), .A3(new_n712), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n819), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(KEYINPUT110), .B(G137), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n834), .B(new_n835), .ZN(G39));
  INV_X1    g650(.A(new_n814), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n331), .A2(new_n837), .A3(new_n398), .A4(new_n731), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n831), .A2(KEYINPUT47), .A3(new_n693), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT47), .B1(new_n831), .B2(new_n693), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(G140), .ZN(G42));
  NOR4_X1   g657(.A1(new_n741), .A2(new_n808), .A3(new_n467), .A4(new_n402), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n759), .B(KEYINPUT49), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n844), .A2(new_n845), .A3(new_n725), .A4(new_n718), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n739), .B(new_n745), .C1(new_n649), .C2(new_n667), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n762), .B1(new_n753), .B2(new_n761), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n764), .A2(KEYINPUT101), .A3(new_n760), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n848), .B(new_n778), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT111), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT111), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n766), .A2(new_n853), .A3(new_n778), .A4(new_n848), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n792), .A2(new_n799), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT106), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n792), .A2(new_n799), .A3(KEYINPUT106), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n792), .A2(new_n745), .A3(new_n732), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n797), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n784), .A2(new_n787), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n708), .A2(new_n402), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n512), .A2(new_n726), .A3(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n863), .A2(new_n681), .A3(new_n724), .A4(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n710), .A3(new_n733), .A4(new_n782), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n710), .A2(new_n782), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(KEYINPUT52), .A3(new_n733), .A4(new_n866), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n860), .A2(new_n862), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n664), .A2(new_n566), .A3(new_n609), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n648), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n512), .A3(new_n615), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n399), .A2(new_n617), .B1(new_n628), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n600), .A2(new_n707), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n704), .A2(new_n877), .A3(new_n656), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n878), .A2(new_n465), .A3(new_n814), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n764), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n876), .A2(new_n690), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n774), .A2(new_n687), .A3(new_n732), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n789), .B2(new_n791), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n881), .A2(new_n805), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n710), .A2(new_n782), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT52), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n855), .A2(new_n872), .A3(new_n886), .A4(new_n890), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n883), .A2(new_n876), .A3(new_n690), .A4(new_n880), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n852), .A2(new_n892), .A3(new_n805), .A4(new_n854), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n871), .A2(new_n869), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n803), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n889), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n847), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n888), .A2(KEYINPUT53), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n851), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n885), .A2(KEYINPUT113), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT113), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n892), .A2(new_n901), .A3(new_n805), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n872), .A2(new_n899), .A3(new_n900), .A4(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n896), .A2(KEYINPUT112), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT112), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n906), .B(new_n889), .C1(new_n893), .C2(new_n895), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n904), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n897), .B1(new_n908), .B2(new_n847), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT51), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n809), .A2(new_n611), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n775), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n837), .ZN(new_n913));
  INV_X1    g727(.A(new_n841), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n839), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n754), .A2(new_n758), .A3(new_n693), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT114), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n718), .A2(new_n467), .A3(new_n693), .A4(new_n759), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n912), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT50), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n837), .A2(new_n738), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n741), .A2(new_n611), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n923), .A2(new_n725), .A3(new_n924), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n925), .A2(new_n631), .A3(new_n647), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n911), .A2(new_n923), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n774), .A2(new_n687), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n929), .A2(KEYINPUT115), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(KEYINPUT115), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n919), .A2(new_n922), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n917), .A2(new_n918), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n910), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n917), .A2(KEYINPUT51), .A3(new_n932), .A4(new_n922), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n796), .A2(new_n398), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n927), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT117), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n940), .A2(KEYINPUT48), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT48), .B1(new_n940), .B2(new_n941), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n911), .A2(new_n781), .A3(new_n775), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n944), .B(new_n610), .C1(new_n648), .C2(new_n925), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT116), .Z(new_n946));
  NOR3_X1   g760(.A1(new_n942), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  AND4_X1   g761(.A1(new_n909), .A2(new_n935), .A3(new_n936), .A4(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(G952), .A2(G953), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n846), .B1(new_n948), .B2(new_n949), .ZN(G75));
  NAND3_X1  g764(.A1(new_n855), .A2(new_n872), .A3(new_n886), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n906), .B1(new_n951), .B2(new_n889), .ZN(new_n952));
  INV_X1    g766(.A(new_n907), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n903), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n954), .A2(KEYINPUT118), .A3(G210), .A4(G902), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n479), .A2(new_n481), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(new_n488), .Z(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT55), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT56), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n955), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n905), .A2(new_n907), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n314), .B1(new_n962), .B2(new_n903), .ZN(new_n963));
  AOI21_X1  g777(.A(KEYINPUT118), .B1(new_n963), .B2(G210), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n439), .A2(G952), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT119), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT56), .B1(new_n963), .B2(G210), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n958), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n965), .A2(new_n969), .ZN(G51));
  XNOR2_X1  g784(.A(new_n404), .B(KEYINPUT57), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n908), .A2(new_n847), .ZN(new_n972));
  AOI211_X1 g786(.A(KEYINPUT54), .B(new_n904), .C1(new_n905), .C2(new_n907), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n757), .B(KEYINPUT120), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n963), .A2(new_n825), .A3(new_n824), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n966), .B1(new_n976), .B2(new_n977), .ZN(G54));
  NAND2_X1  g792(.A1(KEYINPUT58), .A2(G475), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n963), .A2(new_n563), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n563), .B1(new_n963), .B2(new_n980), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n981), .A2(new_n982), .A3(new_n966), .ZN(G60));
  XNOR2_X1  g797(.A(new_n638), .B(KEYINPUT59), .ZN(new_n984));
  OAI22_X1  g798(.A1(new_n909), .A2(new_n984), .B1(new_n634), .B2(new_n642), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n642), .A2(new_n634), .A3(new_n984), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n972), .B2(new_n973), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n985), .A2(new_n967), .A3(new_n987), .ZN(G63));
  NAND2_X1  g802(.A1(G217), .A2(G902), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT60), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n676), .ZN(new_n992));
  INV_X1    g806(.A(new_n679), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n954), .B(new_n991), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n383), .B1(new_n908), .B2(new_n990), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n994), .A2(new_n967), .A3(new_n995), .ZN(new_n996));
  XNOR2_X1  g810(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n994), .A2(new_n967), .A3(new_n995), .A4(new_n997), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(G66));
  AOI21_X1  g815(.A(new_n439), .B1(new_n614), .B2(G224), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n876), .A2(new_n690), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n855), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1002), .B1(new_n1004), .B2(new_n439), .ZN(new_n1005));
  INV_X1    g819(.A(G898), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n956), .B1(new_n1006), .B2(G953), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1005), .B(new_n1007), .ZN(G69));
  NAND2_X1  g822(.A1(new_n252), .A2(new_n257), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT122), .Z(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(new_n549), .Z(new_n1011));
  NAND2_X1  g825(.A1(new_n834), .A2(new_n842), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n833), .A2(new_n512), .A3(new_n726), .A4(new_n937), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n870), .A2(new_n733), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n1014), .A2(new_n805), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1013), .A2(new_n803), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n439), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT126), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n705), .A2(G953), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT125), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1017), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1018), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1011), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(G227), .A2(G900), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(G953), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1011), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT123), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n837), .B1(new_n1029), .B2(new_n874), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n1030), .B(new_n745), .C1(new_n1029), .C2(new_n874), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1031), .A2(new_n713), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1032), .B(KEYINPUT124), .ZN(new_n1033));
  AND3_X1   g847(.A1(new_n729), .A2(KEYINPUT62), .A3(new_n1014), .ZN(new_n1034));
  AOI21_X1  g848(.A(KEYINPUT62), .B1(new_n729), .B2(new_n1014), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n1036), .A2(new_n1012), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1028), .B1(new_n1037), .B2(G953), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1025), .A2(new_n1027), .A3(new_n1038), .ZN(new_n1039));
  AND3_X1   g853(.A1(new_n1013), .A2(new_n803), .A3(new_n1015), .ZN(new_n1040));
  AOI22_X1  g854(.A1(new_n915), .A2(new_n838), .B1(new_n819), .B2(new_n833), .ZN(new_n1041));
  AOI21_X1  g855(.A(G953), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g856(.A(KEYINPUT126), .B1(new_n1042), .B2(new_n1020), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(new_n1022), .ZN(new_n1044));
  OAI211_X1 g858(.A(G953), .B(new_n1026), .C1(new_n1044), .C2(new_n1028), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1039), .A2(new_n1045), .ZN(G72));
  INV_X1    g860(.A(new_n1004), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1037), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g862(.A1(G472), .A2(G902), .ZN(new_n1049));
  XOR2_X1   g863(.A(new_n1049), .B(KEYINPUT63), .Z(new_n1050));
  NAND2_X1  g864(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n891), .A2(new_n896), .ZN(new_n1052));
  INV_X1    g866(.A(new_n1050), .ZN(new_n1053));
  OR2_X1    g867(.A1(new_n326), .A2(new_n286), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n289), .A2(new_n291), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI22_X1  g870(.A1(new_n1051), .A2(new_n720), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g871(.A(new_n966), .ZN(new_n1058));
  NOR2_X1   g872(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n1053), .B1(new_n1059), .B2(new_n1047), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n326), .A2(new_n303), .ZN(new_n1061));
  OAI21_X1  g875(.A(new_n1058), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g876(.A(KEYINPUT127), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g878(.A(KEYINPUT127), .B(new_n1058), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1065));
  AND3_X1   g879(.A1(new_n1057), .A2(new_n1064), .A3(new_n1065), .ZN(G57));
endmodule


