//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1052, new_n1053;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G228gat), .A2(G233gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT72), .B(G211gat), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT22), .B1(new_n209), .B2(G218gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(G197gat), .B(G204gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n208), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G218gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT72), .ZN(new_n215));
  INV_X1    g014(.A(G211gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n207), .B(new_n211), .C1(new_n219), .C2(KEYINPUT22), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n213), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT29), .ZN(new_n222));
  AND2_X1   g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT75), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G141gat), .ZN(new_n226));
  INV_X1    g025(.A(G148gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n229));
  NAND2_X1  g028(.A1(G141gat), .A2(G148gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n225), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G155gat), .B(G162gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G155gat), .ZN(new_n237));
  INV_X1    g036(.A(G162gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n232), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(new_n237), .B2(new_n238), .ZN(new_n240));
  XNOR2_X1  g039(.A(G141gat), .B(G148gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n236), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n221), .A2(new_n222), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT83), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT2), .B1(new_n241), .B2(KEYINPUT75), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n234), .B1(new_n247), .B2(new_n231), .ZN(new_n248));
  INV_X1    g047(.A(new_n243), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT3), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n245), .A2(new_n246), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n246), .B1(new_n245), .B2(new_n250), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT84), .ZN(new_n254));
  AOI221_X4 g053(.A(KEYINPUT3), .B1(new_n240), .B2(new_n242), .C1(new_n233), .C2(new_n235), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(KEYINPUT29), .ZN(new_n256));
  OAI211_X1 g055(.A(KEYINPUT84), .B(new_n222), .C1(new_n244), .C2(KEYINPUT3), .ZN(new_n257));
  INV_X1    g056(.A(new_n220), .ZN(new_n258));
  AND2_X1   g057(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n260));
  OAI21_X1  g059(.A(G218gat), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT22), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n207), .B1(new_n263), .B2(new_n211), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n256), .A2(new_n257), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n206), .B1(new_n253), .B2(new_n266), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n233), .A2(new_n235), .B1(new_n242), .B2(new_n240), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT3), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT29), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT82), .B1(new_n270), .B2(new_n221), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n272), .B(new_n265), .C1(new_n255), .C2(KEYINPUT29), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n206), .A3(new_n273), .ZN(new_n274));
  AOI221_X4 g073(.A(KEYINPUT76), .B1(new_n240), .B2(new_n242), .C1(new_n233), .C2(new_n235), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT76), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n276), .B1(new_n236), .B2(new_n243), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT29), .B1(new_n264), .B2(KEYINPUT80), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT80), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n213), .A2(new_n281), .A3(new_n220), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT81), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n280), .A2(new_n282), .A3(KEYINPUT81), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n269), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n274), .B1(new_n279), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n205), .B1(new_n267), .B2(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n271), .A2(new_n206), .A3(new_n273), .ZN(new_n290));
  INV_X1    g089(.A(new_n286), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT81), .B1(new_n280), .B2(new_n282), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT3), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n290), .B1(new_n293), .B2(new_n278), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n222), .B1(new_n248), .B2(new_n249), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n250), .B1(new_n295), .B2(new_n265), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT83), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n245), .A2(new_n246), .A3(new_n250), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n266), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n206), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n294), .A2(new_n301), .A3(G22gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n289), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT79), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n204), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n204), .ZN(new_n306));
  AOI211_X1 g105(.A(KEYINPUT79), .B(new_n306), .C1(new_n289), .C2(new_n302), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT65), .ZN(new_n309));
  NOR2_X1   g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT66), .B1(new_n310), .B2(KEYINPUT23), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT66), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n312), .B(new_n313), .C1(G169gat), .C2(G176gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(G183gat), .B(G190gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n311), .B(new_n314), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G169gat), .ZN(new_n318));
  INV_X1    g117(.A(G176gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT23), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(G183gat), .A3(G190gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n309), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT25), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT25), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n309), .B(new_n326), .C1(new_n317), .C2(new_n323), .ZN(new_n327));
  INV_X1    g126(.A(G183gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT27), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT27), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G183gat), .ZN(new_n331));
  INV_X1    g130(.A(G190gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT28), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT26), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n310), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n322), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n328), .B2(new_n332), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT28), .B1(new_n333), .B2(new_n334), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n325), .A2(new_n327), .B1(new_n335), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G134gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT68), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT68), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G134gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n347), .A3(G127gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n348), .B1(G127gat), .B2(new_n344), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT1), .ZN(new_n350));
  INV_X1    g149(.A(G120gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G113gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n351), .A2(G113gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT69), .B(G113gat), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n352), .B1(new_n357), .B2(new_n351), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n350), .B1(new_n344), .B2(G127gat), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n359), .B1(G127gat), .B2(new_n344), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n342), .A2(new_n335), .ZN(new_n364));
  INV_X1    g163(.A(new_n327), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n332), .A2(G183gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n328), .A2(G190gat), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT24), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n366), .A2(new_n369), .A3(new_n311), .A4(new_n314), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n326), .B1(new_n370), .B2(new_n309), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n364), .B1(new_n365), .B2(new_n371), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n349), .A2(new_n355), .B1(new_n358), .B2(new_n360), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G227gat), .A2(G233gat), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n375), .B(KEYINPUT64), .Z(new_n376));
  NAND3_X1  g175(.A1(new_n363), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT32), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT70), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT70), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n377), .A2(new_n380), .A3(KEYINPUT32), .ZN(new_n381));
  XNOR2_X1  g180(.A(G15gat), .B(G43gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(G71gat), .B(G99gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT33), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n384), .B1(new_n377), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n379), .A2(new_n381), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT34), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n363), .A2(new_n374), .ZN(new_n389));
  INV_X1    g188(.A(new_n376), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI211_X1 g190(.A(KEYINPUT34), .B(new_n376), .C1(new_n363), .C2(new_n374), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n377), .B(KEYINPUT32), .C1(new_n385), .C2(new_n384), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n387), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n393), .B1(new_n387), .B2(new_n394), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT5), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n373), .B(new_n268), .ZN(new_n400));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n399), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n362), .B1(new_n268), .B2(new_n269), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n404), .A2(new_n255), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(new_n244), .B2(new_n362), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n408), .A3(new_n401), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n279), .A2(new_n407), .A3(new_n362), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n403), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n407), .B1(new_n373), .B2(new_n268), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT76), .B1(new_n248), .B2(new_n249), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n236), .A2(new_n276), .A3(new_n243), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n413), .A2(new_n407), .A3(new_n373), .A4(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n412), .B1(new_n415), .B2(KEYINPUT77), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT77), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n278), .A2(new_n417), .A3(new_n407), .A4(new_n373), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n399), .B(new_n401), .C1(new_n404), .C2(new_n255), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT78), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n423));
  AOI211_X1 g222(.A(new_n423), .B(new_n420), .C1(new_n416), .C2(new_n418), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n411), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G1gat), .B(G29gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT0), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(G57gat), .ZN(new_n428));
  INV_X1    g227(.A(G85gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n430), .B(new_n411), .C1(new_n422), .C2(new_n424), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n425), .A2(KEYINPUT6), .A3(new_n431), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G226gat), .A2(G233gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(new_n343), .B2(KEYINPUT29), .ZN(new_n439));
  INV_X1    g238(.A(new_n438), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n372), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n221), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(G92gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT74), .B(G64gat), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n444), .B(new_n445), .Z(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n440), .B1(new_n372), .B2(new_n222), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT73), .B1(new_n343), .B2(new_n438), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT73), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n372), .A2(new_n450), .A3(new_n440), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n448), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n442), .B(new_n447), .C1(new_n452), .C2(new_n221), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT30), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n452), .A2(new_n221), .ZN(new_n456));
  INV_X1    g255(.A(new_n442), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n446), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n343), .A2(KEYINPUT73), .A3(new_n438), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n450), .B1(new_n372), .B2(new_n440), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n439), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n265), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n462), .A2(KEYINPUT30), .A3(new_n442), .A4(new_n447), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n455), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n308), .A2(new_n398), .A3(new_n437), .A4(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT35), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n294), .A2(new_n301), .A3(G22gat), .ZN(new_n470));
  AOI21_X1  g269(.A(G22gat), .B1(new_n294), .B2(new_n301), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n304), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n306), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n303), .A2(new_n304), .A3(new_n204), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n435), .A2(new_n436), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT37), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n477), .B(new_n442), .C1(new_n452), .C2(new_n221), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n446), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT38), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n449), .A2(new_n451), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n265), .B1(new_n481), .B2(new_n439), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n439), .A2(new_n265), .A3(new_n441), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT37), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n480), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n453), .B1(new_n479), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n478), .A2(new_n446), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n477), .B1(new_n462), .B2(new_n442), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n486), .B1(KEYINPUT38), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT40), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n405), .B1(new_n416), .B2(new_n418), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n494), .A2(KEYINPUT39), .A3(new_n401), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n495), .A2(KEYINPUT87), .A3(new_n431), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT87), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n419), .A2(new_n406), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT39), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(new_n402), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n500), .B2(new_n430), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT39), .B1(new_n400), .B2(new_n402), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n498), .B2(new_n402), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n493), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n493), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(new_n496), .B2(new_n501), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT88), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n464), .A2(new_n432), .ZN(new_n510));
  OAI211_X1 g309(.A(KEYINPUT88), .B(new_n506), .C1(new_n496), .C2(new_n501), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n505), .A2(new_n509), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n492), .A2(KEYINPUT89), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT89), .B1(new_n492), .B2(new_n512), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT85), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n305), .B2(new_n307), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n473), .A2(KEYINPUT85), .A3(new_n474), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n420), .B1(new_n416), .B2(new_n418), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT78), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n430), .B1(new_n521), .B2(new_n411), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n434), .A2(new_n433), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n436), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n465), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n519), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT71), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n530), .B(new_n531), .C1(new_n396), .C2(new_n397), .ZN(new_n532));
  INV_X1    g331(.A(new_n397), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n533), .A2(new_n528), .A3(new_n529), .A4(new_n395), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT86), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n527), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n517), .A2(new_n518), .B1(new_n437), .B2(new_n465), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT86), .B1(new_n539), .B2(new_n535), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n469), .B1(new_n515), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT97), .B(G183gat), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G71gat), .A2(G78gat), .ZN(new_n545));
  OR2_X1    g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT9), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G57gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(G64gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT95), .ZN(new_n551));
  INV_X1    g350(.A(G64gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(G57gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT96), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n548), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n550), .A2(new_n553), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n545), .B(new_n546), .C1(new_n556), .C2(new_n547), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(KEYINPUT21), .ZN(new_n560));
  XNOR2_X1  g359(.A(G127gat), .B(G155gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(new_n216), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n216), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n566));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n566), .B(new_n567), .Z(new_n568));
  NAND3_X1  g367(.A1(new_n564), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n568), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n562), .A2(new_n216), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n570), .B1(new_n571), .B2(new_n563), .ZN(new_n572));
  XNOR2_X1  g371(.A(G15gat), .B(G22gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT93), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT16), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n575), .B1(new_n576), .B2(G1gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n573), .B(KEYINPUT93), .ZN(new_n578));
  INV_X1    g377(.A(G1gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(G8gat), .ZN(new_n582));
  INV_X1    g381(.A(G8gat), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n577), .A2(new_n583), .A3(new_n580), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n585), .B1(KEYINPUT21), .B2(new_n559), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n572), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n587), .B1(new_n569), .B2(new_n572), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n544), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n569), .A2(new_n572), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n586), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(new_n543), .A3(new_n588), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n596), .B(KEYINPUT98), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n598), .A2(KEYINPUT41), .ZN(new_n599));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT7), .ZN(new_n604));
  OAI211_X1 g403(.A(G85gat), .B(G92gat), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT100), .B(G92gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n608), .A2(new_n429), .B1(KEYINPUT8), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G99gat), .B(G106gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n607), .A2(new_n612), .A3(new_n610), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G43gat), .B(G50gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT91), .B(G29gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(G36gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(G29gat), .A2(G36gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT14), .ZN(new_n624));
  OAI211_X1 g423(.A(KEYINPUT15), .B(new_n619), .C1(new_n622), .C2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n619), .A2(KEYINPUT15), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n619), .A2(KEYINPUT15), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .A4(new_n621), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n614), .A2(KEYINPUT101), .A3(new_n615), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n618), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n598), .A2(KEYINPUT41), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n625), .A2(new_n629), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT17), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(KEYINPUT92), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT92), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(KEYINPUT17), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(KEYINPUT17), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n630), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n618), .A2(new_n631), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(G190gat), .B1(new_n634), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n618), .A2(new_n631), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n637), .A2(new_n642), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n647), .A2(new_n332), .A3(new_n632), .A4(new_n633), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n644), .A2(G218gat), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(G218gat), .B1(new_n644), .B2(new_n648), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n602), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT103), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n653), .B(new_n602), .C1(new_n649), .C2(new_n650), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n644), .A2(new_n648), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n214), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n644), .A2(new_n648), .A3(G218gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(new_n601), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n656), .A2(KEYINPUT102), .A3(new_n601), .A4(new_n657), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n652), .A2(new_n654), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n595), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n642), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n640), .B1(new_n630), .B2(new_n641), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n582), .B(new_n584), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G229gat), .A2(G233gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n585), .A2(new_n630), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT18), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n582), .A2(new_n635), .A3(new_n584), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n667), .B(KEYINPUT13), .Z(new_n673));
  AOI22_X1  g472(.A1(new_n669), .A2(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(G169gat), .B(G197gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G113gat), .B(G141gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT12), .Z(new_n680));
  NAND4_X1  g479(.A1(new_n666), .A2(KEYINPUT18), .A3(new_n667), .A4(new_n668), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n674), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT94), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT94), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n674), .A2(new_n684), .A3(new_n680), .A4(new_n681), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n674), .A2(new_n681), .ZN(new_n686));
  INV_X1    g485(.A(new_n680), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n683), .A2(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(G120gat), .B(G148gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(G176gat), .ZN(new_n690));
  INV_X1    g489(.A(G204gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n558), .B(KEYINPUT104), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n694), .A2(new_n616), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n616), .B1(new_n696), .B2(new_n558), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(G230gat), .ZN(new_n699));
  INV_X1    g498(.A(G233gat), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT10), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n704), .B(new_n697), .C1(new_n694), .C2(new_n616), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n618), .A2(KEYINPUT10), .A3(new_n559), .A4(new_n631), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n701), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n693), .B1(new_n703), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n706), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n702), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n710), .B(new_n692), .C1(new_n702), .C2(new_n698), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n663), .A2(new_n688), .A3(new_n712), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n542), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n476), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g515(.A(KEYINPUT16), .B(G8gat), .Z(new_n717));
  NAND3_X1  g516(.A1(new_n714), .A2(new_n464), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n714), .ZN(new_n721));
  OAI21_X1  g520(.A(G8gat), .B1(new_n721), .B2(new_n465), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n719), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n720), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1325gat));
  INV_X1    g525(.A(new_n398), .ZN(new_n727));
  OR3_X1    g526(.A1(new_n721), .A2(G15gat), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G15gat), .B1(new_n721), .B2(new_n536), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1326gat));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n519), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT43), .B(G22gat), .Z(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT106), .Z(new_n733));
  XNOR2_X1  g532(.A(new_n731), .B(new_n733), .ZN(G1327gat));
  NAND2_X1  g533(.A1(new_n652), .A2(new_n654), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n660), .A2(new_n661), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n542), .A2(new_n737), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n595), .A2(new_n688), .A3(new_n712), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n437), .A2(new_n620), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT45), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n738), .A2(KEYINPUT44), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n305), .A2(new_n307), .A3(new_n516), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT85), .B1(new_n473), .B2(new_n474), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n526), .B(KEYINPUT107), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT107), .B1(new_n519), .B2(new_n526), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n536), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n469), .B1(new_n515), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n735), .A2(new_n736), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n735), .B2(new_n736), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n752), .A2(new_n753), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n740), .B1(new_n745), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n620), .B1(new_n760), .B2(new_n437), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n761), .ZN(G1328gat));
  OAI21_X1  g561(.A(G36gat), .B1(new_n760), .B2(new_n465), .ZN(new_n763));
  NOR4_X1   g562(.A1(new_n738), .A2(G36gat), .A3(new_n465), .A4(new_n740), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT46), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1329gat));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n753), .B1(new_n542), .B2(new_n737), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n527), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n535), .B1(new_n770), .B2(new_n748), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT89), .ZN(new_n772));
  AND4_X1   g571(.A1(new_n505), .A2(new_n509), .A3(new_n510), .A4(new_n511), .ZN(new_n773));
  OAI21_X1  g572(.A(KEYINPUT38), .B1(new_n479), .B2(new_n488), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n774), .B(new_n453), .C1(new_n479), .C2(new_n485), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n308), .B1(new_n775), .B2(new_n437), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n772), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n492), .A2(KEYINPUT89), .A3(new_n512), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n468), .B1(new_n771), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n757), .A2(new_n753), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n535), .B(new_n739), .C1(new_n768), .C2(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n783), .A2(G43gat), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n727), .A2(G43gat), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n741), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n767), .B(KEYINPUT47), .C1(new_n784), .C2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n783), .A2(G43gat), .B1(new_n741), .B2(new_n785), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(KEYINPUT109), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n787), .A2(new_n790), .ZN(G1330gat));
  INV_X1    g590(.A(G50gat), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n759), .B2(new_n519), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n741), .A2(new_n792), .A3(new_n519), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(KEYINPUT110), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(KEYINPUT48), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(KEYINPUT48), .A2(G50gat), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n759), .B2(new_n475), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n795), .A2(KEYINPUT48), .B1(new_n798), .B2(new_n800), .ZN(G1331gat));
  NAND2_X1  g600(.A1(new_n683), .A2(new_n685), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n686), .A2(new_n687), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n712), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n663), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n752), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(new_n437), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(new_n549), .ZN(G1332gat));
  NOR2_X1   g608(.A1(new_n807), .A2(new_n465), .ZN(new_n810));
  NOR2_X1   g609(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n811));
  AND2_X1   g610(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n810), .B2(new_n811), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT111), .ZN(G1333gat));
  NOR3_X1   g614(.A1(new_n807), .A2(G71gat), .A3(new_n727), .ZN(new_n816));
  INV_X1    g615(.A(new_n807), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n535), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n816), .B1(G71gat), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n519), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g621(.A1(new_n595), .A2(new_n804), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n662), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT51), .B1(new_n780), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n752), .A2(new_n828), .A3(new_n825), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n827), .A2(new_n712), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n830), .A2(new_n429), .A3(new_n476), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n824), .A2(new_n805), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n833), .B1(new_n768), .B2(new_n782), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n834), .B2(new_n437), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G85gat), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n834), .A2(new_n832), .A3(new_n437), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n831), .B1(new_n836), .B2(new_n837), .ZN(G1336gat));
  INV_X1    g637(.A(G92gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n830), .A2(new_n839), .A3(new_n464), .ZN(new_n840));
  INV_X1    g639(.A(new_n608), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n841), .B1(new_n834), .B2(new_n465), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT52), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n840), .A2(new_n842), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(G1337gat));
  XOR2_X1   g647(.A(KEYINPUT114), .B(G99gat), .Z(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n834), .B2(new_n536), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n727), .A2(new_n849), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n830), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(G1338gat));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n519), .B(new_n833), .C1(new_n768), .C2(new_n782), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(G106gat), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n752), .A2(new_n825), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n805), .B1(new_n857), .B2(KEYINPUT51), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n308), .A2(G106gat), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n858), .A2(KEYINPUT115), .A3(new_n829), .A4(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n854), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n827), .A2(new_n829), .A3(new_n712), .A4(new_n859), .ZN(new_n862));
  NAND2_X1  g661(.A1(KEYINPUT115), .A2(KEYINPUT53), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n475), .B(new_n833), .C1(new_n768), .C2(new_n782), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n854), .A2(G106gat), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT116), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n865), .A2(new_n866), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n862), .A3(new_n863), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n871));
  INV_X1    g670(.A(new_n862), .ZN(new_n872));
  AOI22_X1  g671(.A1(new_n872), .A2(KEYINPUT115), .B1(new_n855), .B2(G106gat), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n870), .B(new_n871), .C1(new_n873), .C2(new_n854), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n868), .A2(new_n874), .ZN(G1339gat));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n876));
  INV_X1    g675(.A(new_n595), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n737), .A2(KEYINPUT108), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n662), .A2(new_n754), .ZN(new_n879));
  INV_X1    g678(.A(new_n679), .ZN(new_n880));
  INV_X1    g679(.A(new_n673), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n668), .A2(new_n671), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT117), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n666), .A2(new_n668), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(G229gat), .A3(G233gat), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n683), .A2(new_n685), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n705), .A2(new_n706), .A3(new_n701), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n710), .A2(KEYINPUT54), .A3(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n692), .B1(new_n707), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n889), .A2(KEYINPUT55), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT55), .B1(new_n889), .B2(new_n891), .ZN(new_n893));
  INV_X1    g692(.A(new_n711), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n887), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n878), .A2(new_n879), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n892), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(new_n893), .A3(new_n894), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n899), .A2(new_n804), .B1(new_n887), .B2(new_n712), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n900), .B1(new_n878), .B2(new_n879), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n877), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n663), .A2(new_n804), .A3(new_n712), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n876), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n878), .A2(new_n879), .A3(new_n896), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n886), .A2(new_n880), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n802), .A2(new_n712), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n895), .A2(new_n892), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(new_n688), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n755), .B2(new_n756), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n595), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n912), .A2(KEYINPUT118), .A3(new_n903), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n905), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n437), .A2(new_n464), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n519), .A2(new_n727), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n914), .A2(KEYINPUT119), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n902), .A2(new_n904), .A3(new_n876), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT118), .B1(new_n912), .B2(new_n903), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n918), .A2(new_n919), .A3(new_n915), .A4(new_n916), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n917), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n804), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G113gat), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n727), .A2(new_n475), .A3(new_n464), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n914), .A2(new_n476), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n688), .A2(new_n357), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT120), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n925), .A2(new_n930), .ZN(G1340gat));
  AOI21_X1  g730(.A(G120gat), .B1(new_n927), .B2(new_n712), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n805), .A2(new_n351), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n923), .B2(new_n933), .ZN(G1341gat));
  NAND2_X1  g733(.A1(new_n923), .A2(new_n595), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G127gat), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n905), .A2(new_n913), .A3(new_n437), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n926), .ZN(new_n938));
  OR3_X1    g737(.A1(new_n938), .A2(G127gat), .A3(new_n877), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(G1342gat));
  INV_X1    g739(.A(KEYINPUT56), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n345), .A2(new_n347), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n737), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n941), .B1(new_n927), .B2(new_n944), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n938), .A2(KEYINPUT56), .A3(new_n943), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n917), .A2(new_n737), .A3(new_n922), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT121), .A3(G134gat), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT121), .B1(new_n948), .B2(G134gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G1343gat));
  INV_X1    g750(.A(KEYINPUT57), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n918), .A2(new_n919), .A3(new_n952), .A4(new_n475), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n536), .A2(new_n915), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n910), .A2(new_n662), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n595), .B1(new_n906), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n519), .B1(new_n956), .B2(new_n903), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n954), .B1(new_n957), .B2(KEYINPUT57), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n953), .A2(new_n804), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G141gat), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n937), .A2(new_n475), .A3(new_n465), .A4(new_n536), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n804), .A2(new_n226), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT58), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT58), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n960), .B(new_n965), .C1(new_n961), .C2(new_n962), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1344gat));
  NAND3_X1  g766(.A1(new_n953), .A2(new_n712), .A3(new_n958), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT122), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n227), .A2(KEYINPUT59), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n969), .B1(new_n968), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT59), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n896), .A2(new_n737), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n595), .B1(new_n955), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n519), .B1(new_n976), .B2(new_n903), .ZN(new_n977));
  AND3_X1   g776(.A1(new_n977), .A2(KEYINPUT123), .A3(new_n952), .ZN(new_n978));
  AOI21_X1  g777(.A(KEYINPUT123), .B1(new_n977), .B2(new_n952), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT57), .A4(new_n475), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(new_n954), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n982), .A2(new_n712), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n974), .B1(new_n984), .B2(G148gat), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n712), .A2(new_n227), .ZN(new_n986));
  OAI22_X1  g785(.A1(new_n973), .A2(new_n985), .B1(new_n961), .B2(new_n986), .ZN(G1345gat));
  NOR3_X1   g786(.A1(new_n961), .A2(G155gat), .A3(new_n877), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n953), .A2(new_n958), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n237), .B1(new_n989), .B2(new_n595), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n988), .A2(new_n990), .ZN(G1346gat));
  NAND2_X1  g790(.A1(new_n989), .A2(new_n757), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT124), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n989), .A2(KEYINPUT124), .A3(new_n757), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n994), .A2(G162gat), .A3(new_n995), .ZN(new_n996));
  OR3_X1    g795(.A1(new_n961), .A2(G162gat), .A3(new_n662), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n996), .A2(new_n997), .ZN(G1347gat));
  NOR2_X1   g797(.A1(new_n476), .A2(new_n465), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n914), .A2(new_n916), .A3(new_n999), .ZN(new_n1000));
  NOR3_X1   g799(.A1(new_n1000), .A2(new_n318), .A3(new_n688), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n905), .A2(new_n913), .A3(new_n476), .ZN(new_n1002));
  NOR3_X1   g801(.A1(new_n727), .A2(new_n475), .A3(new_n465), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g803(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1005), .A2(new_n804), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1001), .B1(new_n1006), .B2(new_n318), .ZN(G1348gat));
  OAI21_X1  g806(.A(G176gat), .B1(new_n1000), .B2(new_n805), .ZN(new_n1008));
  INV_X1    g807(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n712), .A2(new_n319), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n1004), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g810(.A(KEYINPUT125), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g811(.A(KEYINPUT125), .ZN(new_n1013));
  OAI211_X1 g812(.A(new_n1008), .B(new_n1013), .C1(new_n1004), .C2(new_n1010), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1012), .A2(new_n1014), .ZN(G1349gat));
  OAI21_X1  g814(.A(G183gat), .B1(new_n1000), .B2(new_n877), .ZN(new_n1016));
  INV_X1    g815(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n595), .A2(new_n329), .A3(new_n331), .ZN(new_n1018));
  NOR2_X1   g817(.A1(new_n1004), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g818(.A(KEYINPUT60), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g819(.A(KEYINPUT60), .ZN(new_n1021));
  OAI211_X1 g820(.A(new_n1016), .B(new_n1021), .C1(new_n1004), .C2(new_n1018), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1020), .A2(new_n1022), .ZN(G1350gat));
  NAND3_X1  g822(.A1(new_n1005), .A2(new_n332), .A3(new_n757), .ZN(new_n1024));
  INV_X1    g823(.A(KEYINPUT61), .ZN(new_n1025));
  OR2_X1    g824(.A1(new_n1000), .A2(new_n662), .ZN(new_n1026));
  AOI21_X1  g825(.A(new_n1025), .B1(new_n1026), .B2(G190gat), .ZN(new_n1027));
  OAI211_X1 g826(.A(new_n1025), .B(G190gat), .C1(new_n1000), .C2(new_n662), .ZN(new_n1028));
  INV_X1    g827(.A(new_n1028), .ZN(new_n1029));
  OAI21_X1  g828(.A(new_n1024), .B1(new_n1027), .B2(new_n1029), .ZN(G1351gat));
  NOR3_X1   g829(.A1(new_n535), .A2(new_n308), .A3(new_n465), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n1002), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g831(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g832(.A(G197gat), .B1(new_n1033), .B2(new_n804), .ZN(new_n1034));
  NAND2_X1  g833(.A1(new_n536), .A2(new_n999), .ZN(new_n1035));
  XNOR2_X1  g834(.A(new_n1035), .B(KEYINPUT126), .ZN(new_n1036));
  AND3_X1   g835(.A1(new_n1036), .A2(G197gat), .A3(new_n804), .ZN(new_n1037));
  AOI21_X1  g836(.A(new_n1034), .B1(new_n982), .B2(new_n1037), .ZN(G1352gat));
  NOR2_X1   g837(.A1(new_n805), .A2(G204gat), .ZN(new_n1039));
  INV_X1    g838(.A(new_n1039), .ZN(new_n1040));
  OR3_X1    g839(.A1(new_n1032), .A2(KEYINPUT62), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g840(.A(KEYINPUT62), .B1(new_n1032), .B2(new_n1040), .ZN(new_n1042));
  AND3_X1   g841(.A1(new_n982), .A2(new_n712), .A3(new_n1036), .ZN(new_n1043));
  OAI211_X1 g842(.A(new_n1041), .B(new_n1042), .C1(new_n691), .C2(new_n1043), .ZN(G1353gat));
  NOR2_X1   g843(.A1(new_n1035), .A2(new_n877), .ZN(new_n1045));
  AOI21_X1  g844(.A(new_n216), .B1(new_n982), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g845(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n1047));
  NAND2_X1  g846(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OR3_X1    g847(.A1(new_n1032), .A2(new_n209), .A3(new_n877), .ZN(new_n1049));
  XNOR2_X1  g848(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1050));
  OAI211_X1 g849(.A(new_n1048), .B(new_n1049), .C1(new_n1046), .C2(new_n1050), .ZN(G1354gat));
  AOI21_X1  g850(.A(G218gat), .B1(new_n1033), .B2(new_n757), .ZN(new_n1052));
  AND3_X1   g851(.A1(new_n1036), .A2(G218gat), .A3(new_n737), .ZN(new_n1053));
  AOI21_X1  g852(.A(new_n1052), .B1(new_n982), .B2(new_n1053), .ZN(G1355gat));
endmodule


