//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n553, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT65), .B1(new_n465), .B2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(new_n462), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G101), .ZN(new_n470));
  OAI22_X1  g045(.A1(new_n463), .A2(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n461), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n462), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT66), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n478), .A2(new_n462), .ZN(new_n482));
  MUX2_X1   g057(.A(G100), .B(G112), .S(G2105), .Z(new_n483));
  AOI22_X1  g058(.A1(new_n482), .A2(G124), .B1(G2104), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n481), .A2(new_n484), .ZN(G162));
  NAND2_X1  g060(.A1(G114), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G102), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2104), .ZN(new_n489));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n476), .C2(new_n477), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT67), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n462), .C1(new_n476), .C2(new_n477), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n461), .A2(new_n495), .A3(G138), .A4(new_n462), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n489), .A2(new_n490), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n492), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  OR3_X1    g080(.A1(new_n504), .A2(KEYINPUT68), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT68), .B1(new_n504), .B2(new_n505), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n510), .A2(new_n512), .B1(new_n509), .B2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(new_n502), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n506), .A2(new_n507), .B1(new_n515), .B2(G88), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n513), .A2(KEYINPUT70), .A3(G62), .ZN(new_n517));
  INV_X1    g092(.A(G75), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(new_n511), .ZN(new_n519));
  AOI21_X1  g094(.A(KEYINPUT70), .B1(new_n513), .B2(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(G651), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n516), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  OR2_X1    g098(.A1(new_n513), .A2(KEYINPUT71), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n513), .A2(KEYINPUT71), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n515), .A2(G89), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n503), .A2(G51), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n527), .A2(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n524), .A2(G64), .A3(new_n525), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n503), .A2(G52), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n541), .B2(new_n514), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n504), .A2(new_n544), .B1(new_n514), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n548), .B2(new_n536), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT72), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n503), .A2(G53), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(new_n513), .ZN(new_n562));
  XNOR2_X1  g137(.A(KEYINPUT74), .B(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n559), .A2(new_n560), .B1(G651), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n514), .B(KEYINPUT73), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G299));
  OR2_X1    g143(.A1(new_n539), .A2(new_n542), .ZN(G301));
  OAI21_X1  g144(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(G87), .ZN(new_n571));
  INV_X1    g146(.A(G49), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n570), .B(new_n571), .C1(new_n572), .C2(new_n504), .ZN(G288));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n514), .B(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G86), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n566), .A2(KEYINPUT75), .A3(G86), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n562), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G48), .B2(new_n503), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n578), .A2(new_n579), .A3(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n515), .A2(G85), .B1(G47), .B2(new_n503), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT77), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n526), .A2(G60), .ZN(new_n587));
  INV_X1    g162(.A(G72), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n588), .B2(new_n511), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n536), .B1(new_n589), .B2(new_n590), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n586), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G290));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n503), .A2(G54), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n536), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n576), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n566), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n595), .A2(new_n604), .B1(new_n605), .B2(KEYINPUT78), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(KEYINPUT78), .B2(new_n605), .ZN(G284));
  OAI21_X1  g182(.A(new_n606), .B1(KEYINPUT78), .B2(new_n605), .ZN(G321));
  MUX2_X1   g183(.A(G286), .B(G299), .S(new_n595), .Z(G280));
  XNOR2_X1  g184(.A(G280), .B(KEYINPUT79), .ZN(G297));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n603), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n549), .A2(new_n595), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n603), .A2(new_n611), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT80), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n613), .B1(new_n615), .B2(new_n595), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g192(.A(new_n469), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n461), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  INV_X1    g196(.A(G2100), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  MUX2_X1   g199(.A(G99), .B(G111), .S(G2105), .Z(new_n625));
  AOI22_X1  g200(.A1(new_n482), .A2(G123), .B1(G2104), .B2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G135), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n463), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND3_X1  g204(.A1(new_n623), .A2(new_n624), .A3(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2430), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT81), .B(KEYINPUT14), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g213(.A(KEYINPUT82), .B1(new_n634), .B2(new_n635), .ZN(new_n639));
  OAI22_X1  g214(.A1(new_n638), .A2(new_n639), .B1(new_n632), .B2(new_n633), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2443), .B(G2446), .Z(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  OAI21_X1  g223(.A(KEYINPUT83), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT83), .ZN(new_n650));
  INV_X1    g225(.A(new_n648), .ZN(new_n651));
  NAND4_X1  g226(.A1(new_n645), .A2(new_n646), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(G14), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n647), .B2(new_n648), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n653), .A2(new_n655), .ZN(G401));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2084), .B(G2090), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n657), .B2(new_n658), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT84), .B(KEYINPUT17), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n658), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n663), .B1(new_n665), .B2(new_n657), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n657), .A2(new_n660), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n662), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2096), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2100), .ZN(G227));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n674), .A2(new_n677), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  AOI211_X1 g257(.A(new_n679), .B(new_n682), .C1(new_n674), .C2(new_n678), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XOR2_X1   g259(.A(new_n683), .B(new_n684), .Z(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n685), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NOR2_X1   g266(.A1(G168), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n691), .B2(G21), .ZN(new_n693));
  INV_X1    g268(.A(G1966), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT95), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(G5), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G171), .B2(new_n691), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G1961), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT31), .B(G11), .Z(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT30), .B(G28), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI221_X1 g280(.A(new_n705), .B1(new_n703), .B2(new_n628), .C1(new_n693), .C2(new_n694), .ZN(new_n706));
  NOR3_X1   g281(.A1(new_n696), .A2(new_n701), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT96), .ZN(new_n708));
  NOR2_X1   g283(.A1(G29), .A2(G33), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT93), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n479), .A2(G139), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT94), .Z(new_n712));
  AOI22_X1  g287(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n713), .A2(new_n462), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT25), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n710), .B1(new_n719), .B2(new_n703), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G2072), .Z(new_n721));
  NAND2_X1  g296(.A1(G164), .A2(G29), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G27), .B2(G29), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT97), .B(G2078), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n721), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n723), .B2(new_n724), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n700), .B2(new_n699), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT87), .B(G16), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(G19), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n550), .B2(new_n729), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1341), .ZN(new_n732));
  MUX2_X1   g307(.A(G104), .B(G116), .S(G2105), .Z(new_n733));
  AOI22_X1  g308(.A1(new_n482), .A2(G128), .B1(G2104), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G140), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n463), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G29), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n703), .A2(G26), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT28), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G2067), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n703), .A2(G32), .ZN(new_n743));
  AOI22_X1  g318(.A1(G129), .A2(new_n482), .B1(new_n479), .B2(G141), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT26), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n618), .B2(G105), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n743), .B1(new_n748), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT27), .B(G1996), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n471), .A2(new_n474), .A3(new_n703), .ZN(new_n753));
  NOR2_X1   g328(.A1(KEYINPUT24), .A2(G34), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(KEYINPUT24), .A2(G34), .ZN(new_n756));
  AOI21_X1  g331(.A(G29), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n751), .B1(new_n752), .B2(new_n759), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n749), .A2(new_n750), .B1(new_n758), .B2(G2084), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n742), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G29), .A2(G35), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G162), .B2(G29), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT29), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n762), .B1(new_n765), .B2(G2090), .ZN(new_n766));
  NOR2_X1   g341(.A1(G4), .A2(G16), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n603), .B2(G16), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n766), .B1(G1348), .B2(new_n768), .C1(G2090), .C2(new_n765), .ZN(new_n769));
  AOI211_X1 g344(.A(new_n732), .B(new_n769), .C1(G1348), .C2(new_n768), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n728), .A2(G20), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT23), .Z(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G299), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1956), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n727), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n708), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(G305), .A2(new_n691), .ZN(new_n778));
  OR2_X1    g353(.A1(G6), .A2(G16), .ZN(new_n779));
  AND3_X1   g354(.A1(new_n778), .A2(KEYINPUT89), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(KEYINPUT89), .B1(new_n778), .B2(new_n779), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT32), .B(G1981), .Z(new_n784));
  OR2_X1    g359(.A1(G16), .A2(G23), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G288), .B2(new_n691), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT90), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT33), .B(G1976), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n791), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n788), .B2(new_n789), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n783), .A2(new_n784), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n729), .A2(G22), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G166), .B2(new_n729), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1971), .ZN(new_n798));
  INV_X1    g373(.A(new_n784), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n798), .B1(new_n782), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT88), .B(KEYINPUT34), .Z(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT91), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n783), .A2(new_n784), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n792), .A2(new_n794), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n806), .A2(new_n807), .A3(new_n800), .A4(new_n802), .ZN(new_n808));
  NOR2_X1   g383(.A1(G25), .A2(G29), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n479), .A2(G131), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n482), .A2(G119), .ZN(new_n811));
  MUX2_X1   g386(.A(G95), .B(G107), .S(G2105), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G2104), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n809), .B1(new_n815), .B2(G29), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n729), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G24), .B2(new_n729), .ZN(new_n820));
  INV_X1    g395(.A(G1986), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n804), .A2(new_n805), .A3(new_n808), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n808), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n802), .B1(new_n795), .B2(new_n800), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT91), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n829));
  OR3_X1    g404(.A1(new_n825), .A2(new_n826), .A3(KEYINPUT36), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT92), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n828), .A2(new_n831), .A3(KEYINPUT36), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n777), .B1(new_n833), .B2(new_n834), .ZN(G311));
  INV_X1    g410(.A(new_n834), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n828), .A2(KEYINPUT36), .B1(new_n830), .B2(new_n831), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n776), .B1(new_n836), .B2(new_n837), .ZN(G150));
  NAND2_X1  g413(.A1(new_n526), .A2(G67), .ZN(new_n839));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n536), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n503), .A2(G55), .ZN(new_n842));
  INV_X1    g417(.A(G93), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(new_n514), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n549), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n550), .A2(new_n845), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n603), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n854));
  AOI21_X1  g429(.A(G860), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT99), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n846), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(G145));
  XNOR2_X1  g435(.A(new_n748), .B(new_n736), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n491), .B1(new_n494), .B2(new_n496), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n864), .B2(new_n718), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n620), .B(new_n814), .ZN(new_n866));
  MUX2_X1   g441(.A(G106), .B(G118), .S(G2105), .Z(new_n867));
  AOI22_X1  g442(.A1(new_n482), .A2(G130), .B1(G2104), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G142), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n868), .B1(new_n869), .B2(new_n463), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n866), .B(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n719), .A2(KEYINPUT101), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n865), .A2(new_n871), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n628), .B(G160), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(KEYINPUT100), .Z(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(G162), .Z(new_n879));
  AOI21_X1  g454(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(new_n880));
  OR3_X1    g455(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n879), .B1(new_n876), .B2(new_n880), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g460(.A1(new_n846), .A2(G868), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n615), .B(KEYINPUT102), .ZN(new_n887));
  INV_X1    g462(.A(new_n849), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n603), .A2(G299), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT104), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n603), .A2(G299), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT103), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT41), .B1(new_n891), .B2(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n889), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n891), .A2(new_n894), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n900), .B1(new_n889), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G288), .B(KEYINPUT106), .ZN(new_n904));
  NAND2_X1  g479(.A1(G290), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g480(.A(G288), .B(KEYINPUT106), .Z(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n593), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(G166), .B(G305), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n905), .A2(new_n907), .A3(new_n909), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT42), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n903), .B(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n886), .B1(new_n915), .B2(G868), .ZN(G295));
  AOI21_X1  g491(.A(new_n886), .B1(new_n915), .B2(G868), .ZN(G331));
  NAND2_X1  g492(.A1(G301), .A2(KEYINPUT107), .ZN(new_n918));
  OR3_X1    g493(.A1(new_n539), .A2(KEYINPUT107), .A3(new_n542), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(G286), .A3(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n919), .A2(G286), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n849), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n847), .A2(new_n920), .A3(new_n921), .A4(new_n848), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n897), .A2(new_n925), .A3(new_n898), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(new_n927), .A3(new_n924), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n888), .A2(KEYINPUT108), .A3(new_n920), .A4(new_n921), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n901), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n913), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n911), .A2(new_n912), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n897), .A2(new_n898), .A3(new_n925), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n928), .A2(new_n929), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n932), .B(new_n933), .C1(new_n934), .C2(new_n901), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n931), .A2(new_n935), .A3(new_n936), .A4(new_n882), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT44), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n928), .B(new_n929), .C1(new_n901), .C2(new_n896), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n925), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n902), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT41), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n932), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n935), .A2(new_n882), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT109), .B1(new_n939), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n935), .A2(new_n882), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n901), .B1(new_n940), .B2(new_n925), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n940), .A2(new_n943), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n913), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n936), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n953), .A2(new_n938), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n936), .B1(new_n945), .B2(new_n946), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n949), .A2(KEYINPUT43), .A3(new_n931), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI22_X1  g533(.A1(new_n948), .A2(new_n955), .B1(KEYINPUT44), .B2(new_n958), .ZN(G397));
  AND2_X1   g534(.A1(new_n489), .A2(new_n490), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n497), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(KEYINPUT45), .ZN(new_n962));
  INV_X1    g537(.A(G40), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n471), .A2(new_n474), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(G1996), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT46), .Z(new_n967));
  XOR2_X1   g542(.A(new_n965), .B(KEYINPUT110), .Z(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n748), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n736), .B(G2067), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n972), .B(KEYINPUT47), .Z(new_n973));
  INV_X1    g548(.A(new_n966), .ZN(new_n974));
  INV_X1    g549(.A(G1996), .ZN(new_n975));
  OAI221_X1 g550(.A(new_n971), .B1(new_n748), .B2(new_n974), .C1(new_n969), .C2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n815), .A2(new_n817), .ZN(new_n977));
  OAI22_X1  g552(.A1(new_n976), .A2(new_n977), .B1(G2067), .B2(new_n736), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n978), .A2(new_n968), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n814), .B(new_n817), .Z(new_n980));
  AOI21_X1  g555(.A(new_n976), .B1(new_n980), .B2(new_n968), .ZN(new_n981));
  NOR3_X1   g556(.A1(G290), .A2(G1986), .A3(new_n965), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT124), .B(KEYINPUT48), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n982), .B(new_n983), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n973), .B(new_n979), .C1(new_n981), .C2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n862), .B2(G1384), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n497), .A2(new_n960), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(KEYINPUT111), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n990), .A3(new_n964), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(G305), .A2(G1981), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n583), .B1(new_n577), .B2(new_n514), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(G1981), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT113), .ZN(new_n1001));
  AOI211_X1 g576(.A(new_n993), .B(new_n992), .C1(new_n998), .C2(new_n999), .ZN(new_n1002));
  AOI211_X1 g577(.A(G1976), .B(G288), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n995), .B(KEYINPUT114), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n994), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1006));
  INV_X1    g581(.A(G1976), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n994), .B1(new_n1007), .B2(G288), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT112), .B(G1976), .ZN(new_n1009));
  AOI211_X1 g584(.A(KEYINPUT52), .B(new_n1008), .C1(G288), .C2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(KEYINPUT52), .B2(new_n1008), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1006), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G303), .A2(G8), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT55), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT50), .B1(new_n987), .B2(new_n990), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n500), .A2(new_n989), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n964), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n961), .A2(KEYINPUT45), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n964), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT45), .B1(new_n500), .B2(new_n989), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI22_X1  g599(.A1(new_n1020), .A2(G2090), .B1(G1971), .B2(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1025), .A2(G8), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1015), .A2(new_n1026), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1012), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n752), .B(new_n964), .C1(new_n1016), .C2(new_n1019), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G125), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n478), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n473), .ZN(new_n1033));
  OAI21_X1  g608(.A(G2105), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n618), .A2(G101), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n479), .A2(G137), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1034), .A2(new_n1035), .A3(G40), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n987), .A2(new_n990), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT45), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT116), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n500), .A2(new_n1043), .A3(KEYINPUT45), .A4(new_n989), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1966), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(G8), .B1(new_n1030), .B2(new_n1046), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1047), .A2(G286), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1015), .A2(new_n1026), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1012), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT63), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1005), .B(new_n1028), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1037), .B1(KEYINPUT45), .B2(new_n961), .ZN(new_n1053));
  INV_X1    g628(.A(G2078), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n500), .A2(new_n989), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1053), .B(new_n1054), .C1(KEYINPUT45), .C2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1056), .A2(KEYINPUT122), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT122), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT121), .B(G1961), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1020), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1040), .A2(new_n1045), .A3(KEYINPUT53), .A4(new_n1054), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(G171), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n1030), .B2(new_n1046), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT111), .B1(new_n988), .B2(new_n989), .ZN(new_n1070));
  AOI211_X1 g645(.A(new_n986), .B(G1384), .C1(new_n497), .C2(new_n960), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1039), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n964), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n694), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(KEYINPUT118), .A3(new_n1029), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1068), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g651(.A(KEYINPUT51), .B(G8), .C1(new_n1076), .C2(G286), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT119), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n993), .B1(new_n1068), .B2(new_n1075), .ZN(new_n1080));
  NOR2_X1   g655(.A1(G168), .A2(new_n993), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1079), .B(KEYINPUT51), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1047), .A2(KEYINPUT120), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1047), .A2(KEYINPUT120), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1081), .A2(KEYINPUT51), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1078), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1080), .A2(G286), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1087), .A2(KEYINPUT62), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT62), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1066), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1048), .A2(KEYINPUT63), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT56), .B(G2072), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1024), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n987), .A2(new_n990), .A3(KEYINPUT50), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1037), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1094), .B1(G1956), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(KEYINPUT57), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n565), .A2(new_n567), .A3(new_n1100), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n565), .B2(new_n567), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1098), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1106), .B(new_n1094), .C1(G1956), .C2(new_n1097), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1022), .A2(G1996), .A3(new_n1023), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT58), .B(G1341), .Z(new_n1112));
  AND2_X1   g687(.A1(new_n991), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n550), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT59), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n550), .B(new_n1116), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n991), .A2(G2067), .ZN(new_n1118));
  INV_X1    g693(.A(G1348), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n1020), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n604), .A2(KEYINPUT60), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1115), .A2(new_n1117), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1105), .A2(new_n1107), .A3(KEYINPUT61), .ZN(new_n1123));
  AOI211_X1 g698(.A(new_n1118), .B(new_n603), .C1(new_n1020), .C2(new_n1119), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1020), .A2(new_n1119), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1118), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n604), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT60), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1110), .A2(new_n1122), .A3(new_n1123), .A4(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1107), .A2(new_n1127), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1130), .A2(new_n1105), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  OR3_X1    g707(.A1(new_n1060), .A2(G171), .A3(new_n1064), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1060), .ZN(new_n1134));
  NOR4_X1   g709(.A1(new_n1022), .A2(new_n962), .A3(new_n1057), .A4(G2078), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n1020), .B2(new_n1061), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(KEYINPUT54), .B(new_n1133), .C1(new_n1137), .C2(G301), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1132), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1136), .B(G301), .C1(new_n1059), .C2(new_n1058), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1065), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g719(.A(KEYINPUT123), .B(KEYINPUT54), .C1(new_n1065), .C2(new_n1141), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1139), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1092), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1091), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1006), .A2(KEYINPUT115), .A3(new_n1011), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT115), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1012), .A2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1024), .A2(G1971), .ZN(new_n1154));
  INV_X1    g729(.A(G2090), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1154), .B1(new_n1155), .B2(new_n1097), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1014), .B1(new_n1156), .B2(new_n993), .ZN(new_n1157));
  AND4_X1   g732(.A1(new_n1151), .A2(new_n1153), .A3(new_n1157), .A4(new_n1027), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1052), .B1(new_n1150), .B2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n593), .B(G1986), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n981), .B1(new_n965), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n985), .B1(new_n1159), .B2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n1164));
  OR2_X1    g738(.A1(G227), .A2(new_n459), .ZN(new_n1165));
  OAI21_X1  g739(.A(new_n1164), .B1(G401), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g740(.A(new_n1165), .B1(new_n653), .B2(new_n655), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n1167), .A2(KEYINPUT125), .ZN(new_n1168));
  NAND4_X1  g742(.A1(new_n1166), .A2(KEYINPUT126), .A3(new_n689), .A4(new_n1168), .ZN(new_n1169));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n1170));
  OAI21_X1  g744(.A(new_n689), .B1(new_n1167), .B2(KEYINPUT125), .ZN(new_n1171));
  AOI211_X1 g745(.A(new_n1164), .B(new_n1165), .C1(new_n653), .C2(new_n655), .ZN(new_n1172));
  OAI21_X1  g746(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g747(.A1(new_n1169), .A2(new_n1173), .A3(new_n884), .ZN(new_n1174));
  NOR2_X1   g748(.A1(new_n1174), .A2(new_n958), .ZN(G308));
  INV_X1    g749(.A(G308), .ZN(G225));
endmodule


