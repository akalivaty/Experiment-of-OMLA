//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT65), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  AND2_X1   g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G20), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT66), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n211), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT68), .B(G244), .Z(new_n221));
  AOI21_X1  g0021(.A(new_n220), .B1(G77), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT67), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT69), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n222), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(new_n207), .ZN(new_n228));
  AND2_X1   g0028(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n216), .A2(new_n229), .A3(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n202), .A2(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n218), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n242), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(KEYINPUT71), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT71), .A2(G1), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n251), .A2(G13), .A3(G20), .A4(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G116), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n251), .A2(G33), .A3(new_n252), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT72), .B1(new_n207), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G1), .A2(G13), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT72), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n261), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n255), .B1(new_n264), .B2(new_n254), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G283), .ZN(new_n266));
  INV_X1    g0066(.A(G20), .ZN(new_n267));
  INV_X1    g0067(.A(G97), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n266), .B(new_n267), .C1(G33), .C2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT85), .A2(KEYINPUT20), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(G20), .B2(new_n254), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n263), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT85), .A2(KEYINPUT20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n272), .A2(new_n274), .ZN(new_n276));
  AND3_X1   g0076(.A1(new_n265), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n212), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT77), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n258), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n282), .A2(G33), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  MUX2_X1   g0087(.A(G257), .B(G264), .S(G1698), .Z(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G303), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n279), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT5), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n251), .A2(new_n295), .A3(G45), .A4(new_n252), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT70), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n294), .ZN(new_n298));
  NAND2_X1  g0098(.A1(KEYINPUT70), .A2(G41), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT5), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(G270), .B(new_n279), .C1(new_n296), .C2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n252), .ZN(new_n302));
  NOR2_X1   g0102(.A1(KEYINPUT71), .A2(G1), .ZN(new_n303));
  INV_X1    g0103(.A(G45), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT5), .ZN(new_n306));
  INV_X1    g0106(.A(new_n299), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT70), .A2(G41), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G274), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(new_n212), .B2(new_n278), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n305), .A2(new_n309), .A3(new_n311), .A4(new_n295), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n301), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(G200), .B1(new_n293), .B2(new_n313), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n293), .A2(new_n313), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n277), .B(new_n314), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT21), .ZN(new_n318));
  OAI21_X1  g0118(.A(G169), .B1(new_n293), .B2(new_n313), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n318), .B1(new_n277), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n265), .A2(new_n276), .A3(new_n275), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n315), .A2(new_n321), .A3(KEYINPUT21), .A4(G169), .ZN(new_n322));
  INV_X1    g0122(.A(G179), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n293), .A2(new_n323), .A3(new_n313), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n321), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n317), .A2(new_n320), .A3(new_n322), .A4(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n328));
  NOR2_X1   g0128(.A1(G20), .A2(G33), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT8), .B(G58), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT73), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n258), .A2(G20), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n330), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n253), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n335), .A2(new_n263), .B1(new_n202), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n302), .A2(new_n303), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n263), .B1(G20), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n337), .B1(new_n202), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT9), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G1698), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n290), .A2(G222), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G77), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n290), .A2(G1698), .ZN(new_n347));
  INV_X1    g0147(.A(G223), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n345), .B1(new_n346), .B2(new_n290), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n260), .B1(G33), .B2(G41), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n298), .A2(new_n299), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n311), .B(new_n250), .C1(new_n352), .C2(G45), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n305), .A2(new_n350), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n251), .A2(G41), .A3(new_n252), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(G226), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n351), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n357), .A2(G200), .ZN(new_n358));
  NAND2_X1  g0158(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n357), .B2(new_n316), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n328), .B1(new_n343), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n341), .B(KEYINPUT9), .ZN(new_n364));
  INV_X1    g0164(.A(new_n328), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n357), .A2(G179), .ZN(new_n367));
  INV_X1    g0167(.A(G169), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n357), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n341), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n363), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n334), .A2(new_n346), .B1(new_n267), .B2(G68), .ZN(new_n372));
  INV_X1    g0172(.A(new_n329), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n373), .A2(new_n202), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n263), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT11), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n336), .A2(KEYINPUT12), .A3(new_n218), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT12), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n253), .B2(G68), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n340), .A2(new_n218), .B1(new_n376), .B2(new_n375), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n290), .A2(G232), .A3(G1698), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n290), .A2(G226), .A3(new_n344), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G97), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n350), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n251), .A2(G45), .A3(new_n252), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n391), .A2(new_n355), .A3(G238), .A4(new_n279), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n353), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT13), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n393), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT13), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n389), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT76), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT14), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(G169), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n394), .A2(G179), .A3(new_n397), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n400), .B1(new_n398), .B2(G169), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n384), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n398), .A2(G200), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n394), .A2(G190), .A3(new_n397), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n383), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n354), .A2(new_n221), .A3(new_n355), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n410), .A2(new_n353), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n290), .A2(G232), .A3(new_n344), .ZN(new_n412));
  INV_X1    g0212(.A(G107), .ZN(new_n413));
  OAI221_X1 g0213(.A(new_n412), .B1(new_n413), .B2(new_n290), .C1(new_n347), .C2(new_n219), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n350), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G200), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT74), .ZN(new_n418));
  INV_X1    g0218(.A(new_n331), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n329), .B1(G20), .B2(G77), .ZN(new_n420));
  XNOR2_X1  g0220(.A(KEYINPUT15), .B(G87), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n334), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n263), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n339), .A2(G77), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n336), .A2(new_n346), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n417), .A2(new_n418), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n411), .A2(new_n415), .A3(G190), .ZN(new_n428));
  INV_X1    g0228(.A(G200), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n411), .B2(new_n415), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT74), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n427), .A2(new_n428), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n416), .A2(new_n368), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n411), .A2(new_n415), .A3(new_n323), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(new_n431), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n371), .A2(new_n409), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G58), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(new_n218), .ZN(new_n440));
  OAI21_X1  g0240(.A(G20), .B1(new_n440), .B2(new_n201), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n329), .A2(G159), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n285), .A2(new_n286), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT78), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n284), .ZN(new_n447));
  NAND2_X1  g0247(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(G33), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n267), .B1(KEYINPUT79), .B2(KEYINPUT7), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(KEYINPUT79), .A2(KEYINPUT7), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G68), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n451), .B1(new_n445), .B2(new_n449), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(new_n453), .ZN(new_n457));
  OAI211_X1 g0257(.A(KEYINPUT16), .B(new_n444), .C1(new_n455), .C2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT16), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT7), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(G20), .ZN(new_n461));
  AOI21_X1  g0261(.A(G33), .B1(new_n447), .B2(new_n448), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n284), .A2(G33), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n461), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n460), .B1(new_n290), .B2(G20), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n218), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n459), .B1(new_n467), .B2(new_n443), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n458), .A2(new_n263), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n332), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n340), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n332), .A2(new_n253), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT18), .ZN(new_n475));
  NOR2_X1   g0275(.A1(G223), .A2(G1698), .ZN(new_n476));
  INV_X1    g0276(.A(G226), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(G1698), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n445), .A2(new_n478), .A3(new_n449), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G87), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n279), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n391), .A2(new_n355), .A3(G232), .A4(new_n279), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n353), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G179), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n368), .B2(new_n484), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n474), .A2(new_n475), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n475), .B1(new_n474), .B2(new_n486), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR4_X1   g0290(.A1(new_n481), .A2(new_n483), .A3(KEYINPUT80), .A4(G190), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n479), .A2(new_n480), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n350), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n482), .A2(new_n353), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n495), .A3(new_n316), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n429), .B1(new_n481), .B2(new_n483), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT80), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n469), .A2(new_n492), .A3(new_n473), .A4(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT17), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT81), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT80), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n484), .B2(new_n316), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n491), .B1(new_n504), .B2(new_n497), .ZN(new_n505));
  XNOR2_X1  g0305(.A(KEYINPUT81), .B(KEYINPUT17), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n505), .A2(new_n507), .A3(new_n469), .A4(new_n473), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n490), .A2(KEYINPUT82), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT82), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n502), .A2(new_n508), .ZN(new_n512));
  INV_X1    g0312(.A(new_n473), .ZN(new_n513));
  INV_X1    g0313(.A(new_n263), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n218), .B1(new_n456), .B2(new_n453), .ZN(new_n515));
  OAI211_X1 g0315(.A(KEYINPUT79), .B(KEYINPUT7), .C1(new_n287), .C2(G20), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n443), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n517), .B2(KEYINPUT16), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n513), .B1(new_n518), .B2(new_n468), .ZN(new_n519));
  INV_X1    g0319(.A(new_n486), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT18), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n487), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n511), .B1(new_n512), .B2(new_n522), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n438), .A2(new_n510), .A3(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(G264), .B(new_n279), .C1(new_n296), .C2(new_n300), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G294), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  MUX2_X1   g0327(.A(G250), .B(G257), .S(G1698), .Z(new_n528));
  AOI21_X1  g0328(.A(new_n527), .B1(new_n287), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n312), .B(new_n525), .C1(new_n529), .C2(new_n279), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G169), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT88), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n445), .A2(new_n528), .A3(new_n449), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n279), .B1(new_n533), .B2(new_n526), .ZN(new_n534));
  INV_X1    g0334(.A(new_n525), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(KEYINPUT88), .B(new_n525), .C1(new_n529), .C2(new_n279), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n536), .A2(new_n537), .A3(G179), .A4(new_n312), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n539), .A2(new_n463), .A3(new_n267), .A4(G87), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT22), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OR2_X1    g0342(.A1(KEYINPUT86), .A2(KEYINPUT23), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n413), .A2(G20), .ZN(new_n544));
  NAND2_X1  g0344(.A1(KEYINPUT86), .A2(KEYINPUT23), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT87), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G116), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n544), .A2(KEYINPUT23), .B1(G20), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT87), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n543), .A2(new_n544), .A3(new_n551), .A4(new_n545), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n542), .A2(new_n547), .A3(new_n550), .A4(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(G87), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n541), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n445), .A2(new_n449), .A3(new_n267), .A4(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT24), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n546), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n559), .A2(new_n551), .B1(new_n540), .B2(new_n541), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT24), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n549), .B1(new_n546), .B2(KEYINPUT87), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .A4(new_n556), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n263), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n336), .A2(KEYINPUT25), .A3(new_n413), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT25), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n253), .B2(G107), .ZN(new_n568));
  AOI22_X1  g0368(.A1(G107), .A2(new_n264), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n531), .A2(new_n538), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n565), .A2(new_n569), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n536), .A2(new_n537), .A3(new_n312), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n429), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n530), .A2(G190), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n570), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n413), .B1(new_n465), .B2(new_n466), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n329), .A2(G77), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT6), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n580), .A2(new_n268), .A3(G107), .ZN(new_n581));
  XNOR2_X1  g0381(.A(G97), .B(G107), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n579), .B1(new_n583), .B2(new_n267), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n263), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n253), .A2(G97), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n264), .B2(G97), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G244), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(G1698), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n445), .A2(new_n449), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT4), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(KEYINPUT4), .A2(G244), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n539), .A2(new_n463), .A3(new_n594), .A4(new_n344), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n539), .A2(new_n463), .A3(G250), .A4(G1698), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n595), .A2(new_n596), .A3(new_n266), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n279), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(G257), .B(new_n279), .C1(new_n296), .C2(new_n300), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n312), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n368), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n599), .A2(new_n312), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n595), .A2(new_n596), .A3(new_n266), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n592), .B2(new_n591), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n602), .B(new_n323), .C1(new_n279), .C2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n588), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n593), .A2(new_n597), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n350), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(G190), .A3(new_n602), .ZN(new_n609));
  OAI21_X1  g0409(.A(G200), .B1(new_n598), .B2(new_n600), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n609), .A2(new_n610), .A3(new_n585), .A4(new_n587), .ZN(new_n611));
  AND3_X1   g0411(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n212), .B1(new_n612), .B2(new_n261), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n613), .A2(new_n253), .A3(new_n259), .A4(new_n256), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT84), .B1(new_n614), .B2(new_n421), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n253), .A2(new_n256), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  INV_X1    g0417(.A(new_n421), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n514), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n618), .A2(new_n253), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n445), .A2(new_n449), .A3(new_n267), .A4(G68), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT19), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n333), .A2(new_n623), .A3(G97), .ZN(new_n624));
  NOR2_X1   g0424(.A1(G97), .A2(G107), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n625), .A2(new_n554), .B1(new_n387), .B2(new_n267), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n624), .B1(new_n626), .B2(new_n623), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n621), .B1(new_n628), .B2(new_n263), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n620), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(G238), .A2(G1698), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n589), .B2(G1698), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n445), .A2(new_n632), .A3(new_n449), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n548), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n350), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT83), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n391), .A2(new_n636), .A3(G250), .A4(new_n279), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n305), .A2(new_n311), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n391), .A2(G250), .A3(new_n279), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT83), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n635), .A2(new_n640), .A3(new_n323), .A4(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(new_n638), .A3(new_n637), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n279), .B1(new_n633), .B2(new_n548), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n368), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n630), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(G200), .B1(new_n644), .B2(new_n645), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n635), .A2(new_n640), .A3(G190), .A4(new_n642), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n514), .B1(new_n622), .B2(new_n627), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n257), .A2(new_n263), .A3(new_n554), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n650), .A2(new_n651), .A3(new_n621), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n648), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  AND4_X1   g0453(.A1(new_n606), .A2(new_n611), .A3(new_n647), .A4(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n327), .A2(new_n524), .A3(new_n577), .A4(new_n654), .ZN(G372));
  INV_X1    g0455(.A(new_n370), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n398), .A2(G169), .ZN(new_n657));
  INV_X1    g0457(.A(new_n400), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n659), .A2(new_n402), .A3(new_n401), .ZN(new_n660));
  INV_X1    g0460(.A(new_n436), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n660), .A2(new_n384), .B1(new_n408), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n490), .B1(new_n662), .B2(new_n512), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n363), .A2(new_n366), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n656), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n438), .A2(new_n510), .A3(new_n523), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n574), .B1(new_n572), .B2(new_n429), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n565), .A2(new_n569), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n606), .B(new_n611), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT89), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n641), .A2(KEYINPUT83), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n639), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n642), .A2(KEYINPUT89), .A3(new_n638), .A4(new_n637), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n645), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n630), .B(new_n643), .C1(new_n674), .C2(G169), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n649), .B(new_n652), .C1(new_n674), .C2(new_n429), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT90), .B1(new_n669), .B2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n576), .A2(new_n571), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT90), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n611), .A2(new_n606), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n679), .A2(new_n680), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n320), .A2(new_n322), .A3(new_n325), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(new_n570), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n678), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n600), .B1(new_n607), .B2(new_n350), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n687), .A2(new_n323), .B1(new_n585), .B2(new_n587), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n688), .A2(new_n647), .A3(new_n601), .A4(new_n653), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT26), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n588), .A2(new_n601), .A3(new_n605), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n675), .A2(new_n676), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n690), .A2(new_n693), .A3(new_n675), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n686), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n665), .B1(new_n666), .B2(new_n696), .ZN(G369));
  INV_X1    g0497(.A(G330), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n267), .A2(G13), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n338), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G213), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G343), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n277), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n684), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n326), .B2(new_n706), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT91), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT91), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n707), .B(new_n710), .C1(new_n326), .C2(new_n706), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n698), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n570), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n713), .B(new_n680), .C1(new_n571), .C2(new_n705), .ZN(new_n714));
  INV_X1    g0514(.A(new_n705), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n570), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n712), .A2(KEYINPUT92), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT92), .B1(new_n712), .B2(new_n717), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n713), .A2(new_n715), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n684), .A2(new_n705), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n723), .A2(KEYINPUT93), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(KEYINPUT93), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n722), .B1(new_n726), .B2(new_n717), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n721), .A2(new_n727), .ZN(G399));
  INV_X1    g0528(.A(new_n208), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n352), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR4_X1   g0531(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(G1), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(new_n215), .B2(new_n731), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT28), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n695), .A2(new_n705), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT29), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(KEYINPUT94), .A3(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT96), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT95), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n647), .A2(new_n653), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n740), .B(new_n692), .C1(new_n741), .C2(new_n606), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n675), .A2(new_n676), .A3(new_n691), .A4(KEYINPUT26), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n740), .B1(new_n689), .B2(new_n692), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n739), .B(new_n675), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n685), .A2(new_n680), .A3(new_n682), .A4(new_n679), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n692), .B1(new_n741), .B2(new_n606), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT95), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(new_n743), .A3(new_n742), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n739), .B1(new_n751), .B2(new_n675), .ZN(new_n752));
  OAI211_X1 g0552(.A(KEYINPUT29), .B(new_n705), .C1(new_n748), .C2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT94), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n715), .B1(new_n686), .B2(new_n694), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n754), .B1(new_n755), .B2(KEYINPUT29), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n738), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n577), .A2(new_n327), .A3(new_n654), .A4(new_n705), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT30), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n644), .A2(new_n645), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n687), .A2(new_n760), .A3(new_n536), .A4(new_n537), .ZN(new_n761));
  INV_X1    g0561(.A(new_n324), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n536), .A2(new_n537), .ZN(new_n764));
  NOR4_X1   g0564(.A1(new_n598), .A2(new_n644), .A3(new_n600), .A4(new_n645), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n764), .A2(new_n765), .A3(KEYINPUT30), .A4(new_n324), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n672), .A2(new_n673), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n635), .ZN(new_n768));
  AOI21_X1  g0568(.A(G179), .B1(new_n608), .B2(new_n602), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n768), .A2(new_n572), .A3(new_n315), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n763), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n715), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT31), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n771), .A2(KEYINPUT31), .A3(new_n715), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n758), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G330), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n757), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n735), .B1(new_n779), .B2(G1), .ZN(G364));
  AOI21_X1  g0580(.A(new_n250), .B1(new_n699), .B2(G45), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n730), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n712), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n709), .A2(new_n698), .A3(new_n711), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G13), .A2(G33), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G20), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n709), .A2(new_n711), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n290), .A2(new_n208), .ZN(new_n791));
  INV_X1    g0591(.A(G355), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(new_n792), .B1(G116), .B2(new_n208), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT97), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n247), .A2(new_n304), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n287), .A2(new_n729), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G45), .B2(new_n215), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n794), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n260), .B1(G20), .B2(new_n368), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n789), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n783), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(G20), .A2(G179), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT98), .Z(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G190), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n429), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(G200), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G50), .A2(new_n807), .B1(new_n808), .B2(G58), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n805), .A2(new_n316), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n429), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(G200), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G68), .A2(new_n811), .B1(new_n812), .B2(G77), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n316), .A2(G179), .A3(G200), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n267), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n291), .B1(new_n816), .B2(G97), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT32), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n267), .A2(G179), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n819), .A2(new_n316), .A3(new_n429), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n818), .B1(new_n821), .B2(G159), .ZN(new_n822));
  INV_X1    g0622(.A(G159), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n820), .A2(KEYINPUT32), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n819), .A2(G190), .A3(G200), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n554), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n819), .A2(new_n316), .A3(G200), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n413), .ZN(new_n828));
  NOR4_X1   g0628(.A1(new_n822), .A2(new_n824), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n809), .A2(new_n813), .A3(new_n817), .A4(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(KEYINPUT33), .B(G317), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G322), .A2(new_n808), .B1(new_n811), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n812), .A2(G311), .ZN(new_n833));
  INV_X1    g0633(.A(G329), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n291), .B1(new_n820), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(G283), .ZN(new_n836));
  INV_X1    g0636(.A(G303), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n836), .A2(new_n827), .B1(new_n825), .B2(new_n837), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n835), .B(new_n838), .C1(G294), .C2(new_n816), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n807), .A2(G326), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n832), .A2(new_n833), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n830), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n803), .B1(new_n800), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n790), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n786), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G396));
  INV_X1    g0646(.A(KEYINPUT100), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n436), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n434), .A2(KEYINPUT100), .A3(new_n435), .A4(new_n431), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n433), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n695), .A2(new_n705), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n715), .A2(new_n431), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n433), .A2(new_n848), .A3(new_n853), .A4(new_n849), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n661), .A2(new_n715), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n852), .B1(new_n755), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n783), .B1(new_n857), .B2(new_n777), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n777), .B2(new_n857), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n800), .A2(new_n787), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n783), .B1(G77), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT99), .ZN(new_n863));
  AOI22_X1  g0663(.A1(G143), .A2(new_n808), .B1(new_n812), .B2(G159), .ZN(new_n864));
  INV_X1    g0664(.A(G137), .ZN(new_n865));
  INV_X1    g0665(.A(new_n807), .ZN(new_n866));
  INV_X1    g0666(.A(G150), .ZN(new_n867));
  INV_X1    g0667(.A(new_n811), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n864), .B1(new_n865), .B2(new_n866), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT34), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n815), .A2(new_n439), .B1(new_n827), .B2(new_n218), .ZN(new_n871));
  INV_X1    g0671(.A(G132), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n287), .B1(new_n872), .B2(new_n820), .ZN(new_n873));
  INV_X1    g0673(.A(new_n825), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n871), .B(new_n873), .C1(G50), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n827), .A2(new_n554), .ZN(new_n877));
  INV_X1    g0677(.A(G311), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n291), .B1(new_n820), .B2(new_n878), .C1(new_n815), .C2(new_n268), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n877), .B(new_n879), .C1(G107), .C2(new_n874), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n812), .A2(G116), .ZN(new_n881));
  AOI22_X1  g0681(.A1(G294), .A2(new_n808), .B1(new_n807), .B2(G303), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n811), .A2(G283), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n880), .A2(new_n881), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n876), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n863), .B1(new_n885), .B2(new_n800), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n788), .B2(new_n856), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n859), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(G384));
  NOR2_X1   g0689(.A1(new_n214), .A2(new_n254), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n583), .B(KEYINPUT101), .Z(new_n891));
  INV_X1    g0691(.A(KEYINPUT35), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n892), .B2(new_n891), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT36), .ZN(new_n895));
  OR3_X1    g0695(.A1(new_n440), .A2(new_n215), .A3(new_n346), .ZN(new_n896));
  AOI211_X1 g0696(.A(G13), .B(new_n338), .C1(new_n896), .C2(new_n243), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n408), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n384), .B(new_n715), .C1(new_n660), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n384), .A2(new_n715), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n405), .A2(new_n408), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n848), .A2(new_n849), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n705), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n904), .B1(new_n852), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n444), .B1(new_n455), .B2(new_n457), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n459), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n513), .B1(new_n518), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(new_n703), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n512), .B2(new_n522), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n499), .B1(new_n910), .B2(new_n703), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n910), .A2(new_n520), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT37), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n474), .A2(new_n486), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n703), .B(KEYINPUT102), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n474), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT37), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n916), .A2(new_n918), .A3(new_n919), .A4(new_n499), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n912), .A2(KEYINPUT38), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n912), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n907), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  XOR2_X1   g0725(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n918), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n512), .B2(new_n522), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n916), .A2(new_n918), .A3(new_n499), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT37), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n920), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n927), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n925), .B1(new_n922), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n912), .A2(new_n921), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT38), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n912), .A2(KEYINPUT38), .A3(new_n921), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n937), .A2(KEYINPUT39), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n660), .A2(new_n384), .A3(new_n705), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n490), .A2(new_n917), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n924), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n524), .A2(new_n738), .A3(new_n753), .A4(new_n756), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n945), .A2(new_n665), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n944), .B(new_n946), .Z(new_n947));
  INV_X1    g0747(.A(KEYINPUT104), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n922), .B2(new_n933), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n931), .A2(new_n920), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n918), .B1(new_n490), .B2(new_n509), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n926), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(KEYINPUT104), .A3(new_n938), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n776), .A2(new_n903), .A3(new_n856), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n949), .A2(new_n953), .A3(KEYINPUT40), .A4(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT40), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n922), .A2(new_n923), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n854), .A2(new_n855), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n771), .A2(KEYINPUT31), .A3(new_n715), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT31), .B1(new_n771), .B2(new_n715), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n958), .B1(new_n961), .B2(new_n758), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n903), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n956), .B1(new_n957), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n955), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n524), .A2(new_n776), .ZN(new_n966));
  OAI21_X1  g0766(.A(G330), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n966), .B2(new_n965), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n947), .A2(new_n968), .B1(new_n338), .B2(new_n699), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n947), .A2(new_n968), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n898), .B1(new_n969), .B2(new_n970), .ZN(G367));
  OR3_X1    g0771(.A1(new_n719), .A2(KEYINPUT106), .A3(new_n720), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT106), .B1(new_n719), .B2(new_n720), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n715), .A2(new_n588), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n682), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n691), .A2(new_n715), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT45), .B1(new_n727), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n727), .A2(KEYINPUT45), .A3(new_n977), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT44), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n977), .B1(KEYINPUT105), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n727), .A2(new_n984), .B1(KEYINPUT105), .B2(new_n982), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n982), .A2(KEYINPUT105), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n724), .A2(new_n725), .B1(new_n714), .B2(new_n716), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n986), .B(new_n983), .C1(new_n987), .C2(new_n722), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n972), .A2(new_n973), .A3(new_n981), .A4(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n980), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n989), .B1(new_n991), .B2(new_n978), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT106), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n992), .A2(new_n993), .A3(new_n721), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n712), .A2(new_n717), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n712), .A2(new_n717), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(new_n726), .A3(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n726), .B1(new_n996), .B2(new_n997), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n778), .B1(new_n995), .B2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n730), .B(KEYINPUT41), .Z(new_n1003));
  OAI21_X1  g0803(.A(new_n781), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n987), .A2(new_n977), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT42), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n606), .B1(new_n975), .B2(new_n713), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1005), .A2(KEYINPUT42), .B1(new_n705), .B2(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n705), .A2(new_n652), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n679), .A2(new_n1009), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n675), .A2(new_n1009), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n1006), .A2(new_n1008), .B1(KEYINPUT43), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(KEYINPUT43), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1013), .B(new_n1014), .Z(new_n1015));
  INV_X1    g0815(.A(new_n977), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n721), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1015), .B(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1004), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n807), .A2(G143), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n812), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n808), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1020), .B1(new_n1021), .B2(new_n202), .C1(new_n867), .C2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n868), .A2(new_n823), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n290), .B1(new_n820), .B2(new_n865), .C1(new_n346), .C2(new_n827), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n815), .A2(new_n218), .B1(new_n825), .B2(new_n439), .ZN(new_n1026));
  NOR4_X1   g0826(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT108), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n812), .A2(G283), .B1(G107), .B2(new_n816), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT107), .Z(new_n1030));
  INV_X1    g0830(.A(G317), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n450), .B1(new_n1031), .B2(new_n820), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n825), .A2(new_n254), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT46), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n827), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1032), .B(new_n1034), .C1(G97), .C2(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n837), .A2(new_n1022), .B1(new_n866), .B2(new_n878), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G294), .B2(new_n811), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1030), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1028), .A2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT47), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n800), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1010), .A2(new_n789), .A3(new_n1011), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n796), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n801), .B1(new_n208), .B2(new_n421), .C1(new_n1044), .C2(new_n238), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1042), .A2(new_n783), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1019), .A2(new_n1046), .ZN(G387));
  OR2_X1    g0847(.A1(new_n999), .A2(new_n1000), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1048), .A2(new_n778), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1049), .A2(new_n731), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n779), .B2(new_n1001), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT109), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n1048), .B2(new_n781), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1001), .A2(KEYINPUT109), .A3(new_n782), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n714), .A2(new_n716), .A3(new_n789), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n791), .A2(new_n732), .B1(G107), .B2(new_n208), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n235), .A2(new_n304), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n732), .B(new_n304), .C1(new_n218), .C2(new_n346), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT50), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n331), .B2(G50), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n419), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1058), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1062), .A2(new_n1044), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1056), .B1(new_n1057), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n783), .B1(new_n1064), .B2(new_n802), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n808), .A2(G50), .B1(new_n618), .B2(new_n816), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT110), .Z(new_n1067));
  OAI22_X1  g0867(.A1(new_n346), .A2(new_n825), .B1(new_n827), .B2(new_n268), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n287), .B1(new_n867), .B2(new_n820), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n807), .C2(G159), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G68), .A2(new_n812), .B1(new_n811), .B2(new_n470), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1067), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n287), .B1(G326), .B2(new_n821), .ZN(new_n1073));
  INV_X1    g0873(.A(G294), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n815), .A2(new_n836), .B1(new_n825), .B2(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G311), .A2(new_n811), .B1(new_n807), .B2(G322), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n837), .B2(new_n1021), .C1(new_n1031), .C2(new_n1022), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT48), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT49), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1073), .B1(new_n254), .B2(new_n827), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1072), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1065), .B1(new_n1084), .B2(new_n800), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1053), .A2(new_n1054), .B1(new_n1055), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1051), .A2(new_n1086), .ZN(G393));
  AND2_X1   g0887(.A1(new_n990), .A2(new_n994), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(KEYINPUT111), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT111), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n781), .B1(new_n995), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1016), .A2(new_n789), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n242), .A2(new_n796), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1093), .B(new_n801), .C1(new_n268), .C2(new_n208), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n783), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT112), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n290), .B(new_n828), .C1(G322), .C2(new_n821), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n816), .A2(G116), .B1(new_n874), .B2(G283), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n837), .B2(new_n868), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G311), .A2(new_n808), .B1(new_n807), .B2(G317), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT52), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1100), .B(new_n1102), .C1(G294), .C2(new_n812), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1104), .A2(KEYINPUT114), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G150), .A2(new_n807), .B1(new_n808), .B2(G159), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT51), .Z(new_n1107));
  AOI21_X1  g0907(.A(new_n877), .B1(G77), .B2(new_n816), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n450), .B1(G143), .B2(new_n821), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1108), .B(new_n1109), .C1(new_n218), .C2(new_n825), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G50), .A2(new_n811), .B1(new_n812), .B2(new_n419), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1110), .B1(new_n1111), .B2(KEYINPUT113), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1107), .B(new_n1112), .C1(KEYINPUT113), .C2(new_n1111), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1104), .A2(KEYINPUT114), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1105), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1096), .B1(new_n1115), .B2(new_n800), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1089), .A2(new_n1091), .B1(new_n1092), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT115), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n995), .B2(new_n1049), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n779), .A2(new_n1001), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1120), .A2(new_n994), .A3(new_n990), .A4(KEYINPUT115), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT116), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n731), .B1(new_n995), .B2(new_n1049), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1123), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1117), .B1(new_n1125), .B2(new_n1126), .ZN(G390));
  AND4_X1   g0927(.A1(G330), .A2(new_n776), .A3(new_n903), .A4(new_n856), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n949), .A2(new_n953), .A3(new_n940), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n705), .B(new_n851), .C1(new_n748), .C2(new_n752), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n904), .B1(new_n1130), .B2(new_n906), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n715), .B(new_n850), .C1(new_n686), .C2(new_n694), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n906), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n903), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1135), .A2(new_n940), .B1(new_n934), .B2(new_n939), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1128), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT39), .B1(new_n952), .B2(new_n938), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n907), .A2(new_n941), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n962), .A2(G330), .A3(new_n903), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1140), .B(new_n1141), .C1(new_n1131), .C2(new_n1129), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n852), .A2(new_n906), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n903), .B1(new_n962), .B2(G330), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n1128), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT117), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n776), .A2(G330), .A3(new_n856), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n904), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1141), .A2(new_n1149), .A3(new_n1130), .A4(new_n906), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT117), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1151), .B(new_n1144), .C1(new_n1145), .C2(new_n1128), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1147), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n666), .A2(new_n777), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n945), .A2(new_n665), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1143), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1137), .A2(new_n1142), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n730), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1137), .A2(new_n1142), .A3(new_n782), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n787), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n783), .B1(new_n470), .B2(new_n861), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G128), .A2(new_n807), .B1(new_n811), .B2(G137), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT54), .B(G143), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1163), .B1(new_n872), .B2(new_n1022), .C1(new_n1021), .C2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n827), .A2(new_n202), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n291), .B(new_n1166), .C1(G125), .C2(new_n821), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n825), .A2(new_n867), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT53), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(new_n823), .C2(new_n815), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n290), .B(new_n826), .C1(G294), .C2(new_n821), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n816), .A2(G77), .B1(new_n1035), .B2(G68), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(new_n1021), .C2(new_n268), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G107), .A2(new_n811), .B1(new_n808), .B2(G116), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n836), .B2(new_n866), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1165), .A2(new_n1170), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1162), .B1(new_n1176), .B2(new_n800), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1161), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1159), .A2(new_n1160), .A3(new_n1178), .ZN(G378));
  NAND2_X1  g0979(.A1(new_n341), .A2(new_n704), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n371), .B(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1181), .B(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1183), .A2(new_n788), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n268), .A2(new_n868), .B1(new_n866), .B2(new_n254), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n618), .B2(new_n812), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n808), .A2(G107), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT118), .Z(new_n1188));
  NAND3_X1  g0988(.A1(new_n450), .A2(new_n298), .A3(new_n299), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n815), .A2(new_n218), .B1(new_n820), .B2(new_n836), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n825), .A2(new_n346), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n827), .A2(new_n439), .ZN(new_n1192));
  NOR4_X1   g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1186), .A2(new_n1188), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT58), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1189), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n816), .A2(G150), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n825), .B2(new_n1164), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G125), .A2(new_n807), .B1(new_n808), .B2(G128), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n865), .B2(new_n1021), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(G132), .C2(new_n811), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1035), .A2(G159), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n821), .C2(G124), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1198), .B1(new_n1195), .B2(new_n1194), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n800), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1211), .B(new_n783), .C1(G50), .C2(new_n861), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1184), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n955), .A2(G330), .A3(new_n964), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1183), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1183), .A2(G330), .A3(new_n964), .A4(new_n955), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n944), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT119), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1216), .A2(new_n944), .A3(new_n1217), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n944), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1220), .B1(new_n1223), .B2(new_n1219), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1213), .B1(new_n1224), .B2(new_n782), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1158), .A2(new_n1155), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT120), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1158), .A2(KEYINPUT120), .A3(new_n1155), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT57), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n944), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1231), .B1(new_n1234), .B2(new_n1218), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n731), .B1(new_n1230), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT57), .B1(new_n1230), .B2(new_n1224), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT121), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1158), .A2(KEYINPUT120), .A3(new_n1155), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT120), .B1(new_n1158), .B2(new_n1155), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1221), .A2(KEYINPUT119), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1234), .A2(new_n1218), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1243), .B1(new_n1244), .B2(KEYINPUT119), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1238), .B(new_n1231), .C1(new_n1242), .C2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1225), .B1(new_n1239), .B2(new_n1247), .ZN(G375));
  OR2_X1    g1048(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1003), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n1156), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n904), .A2(new_n787), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n783), .B1(G68), .B2(new_n861), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(G132), .A2(new_n807), .B1(new_n812), .B2(G150), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1254), .B1(new_n865), .B2(new_n1022), .C1(new_n868), .C2(new_n1164), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1192), .B1(G159), .B2(new_n874), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n450), .B1(G128), .B2(new_n821), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1256), .B(new_n1257), .C1(new_n202), .C2(new_n815), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n291), .B1(new_n820), .B2(new_n837), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G77), .B2(new_n1035), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n816), .A2(new_n618), .B1(new_n874), .B2(G97), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(new_n1021), .C2(new_n413), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G283), .A2(new_n808), .B1(new_n807), .B2(G294), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n254), .B2(new_n868), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n1255), .A2(new_n1258), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1253), .B1(new_n1265), .B2(new_n800), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1153), .A2(new_n782), .B1(new_n1252), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1251), .A2(new_n1267), .ZN(G381));
  INV_X1    g1068(.A(new_n1225), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1235), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n730), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1231), .B1(new_n1242), .B2(new_n1245), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1271), .B1(new_n1272), .B2(KEYINPUT121), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1269), .B1(new_n1273), .B2(new_n1246), .ZN(new_n1274));
  INV_X1    g1074(.A(G378), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1051), .A2(new_n1086), .A3(new_n845), .ZN(new_n1277));
  OR4_X1    g1077(.A1(G384), .A2(G387), .A3(G381), .A4(new_n1277), .ZN(new_n1278));
  OR3_X1    g1078(.A1(new_n1276), .A2(G390), .A3(new_n1278), .ZN(G407));
  OAI211_X1 g1079(.A(G407), .B(G213), .C1(G343), .C2(new_n1276), .ZN(G409));
  INV_X1    g1080(.A(new_n1277), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n845), .B1(new_n1051), .B2(new_n1086), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(G387), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(G390), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT115), .B1(new_n1088), .B2(new_n1120), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1121), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1124), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT116), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(G387), .A3(new_n1117), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1286), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1284), .B1(new_n1294), .B2(KEYINPUT124), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT124), .ZN(new_n1296));
  AOI211_X1 g1096(.A(new_n1296), .B(new_n1283), .C1(new_n1286), .C2(new_n1293), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1295), .A2(new_n1297), .A3(KEYINPUT126), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT126), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(G390), .A2(new_n1285), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G387), .B1(new_n1292), .B2(new_n1117), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT124), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1283), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1294), .A2(KEYINPUT124), .A3(new_n1284), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1299), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1298), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(G213), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1307), .A2(G343), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(G2897), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1156), .A2(KEYINPUT60), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1310), .A2(new_n1249), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n730), .B1(new_n1310), .B2(new_n1249), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1267), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n888), .ZN(new_n1314));
  OAI211_X1 g1114(.A(G384), .B(new_n1267), .C1(new_n1311), .C2(new_n1312), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT122), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1314), .A2(KEYINPUT122), .A3(new_n1315), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1309), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  AOI22_X1  g1120(.A1(new_n1316), .A2(new_n1317), .B1(G2897), .B2(new_n1308), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1230), .A2(new_n1224), .A3(new_n1250), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1213), .B1(new_n1244), .B2(new_n782), .ZN(new_n1324));
  AOI21_X1  g1124(.A(G378), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1325), .B1(new_n1274), .B2(G378), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1322), .B1(new_n1326), .B2(new_n1308), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT61), .ZN(new_n1328));
  OAI211_X1 g1128(.A(G378), .B(new_n1225), .C1(new_n1239), .C2(new_n1247), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1325), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1308), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1316), .ZN(new_n1333));
  XOR2_X1   g1133(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n1334));
  NAND4_X1  g1134(.A1(new_n1331), .A2(new_n1332), .A3(new_n1333), .A4(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1327), .A2(new_n1328), .A3(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1308), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1337), .B1(new_n1338), .B2(new_n1333), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1306), .B1(new_n1336), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT63), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1338), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1341), .B1(new_n1342), .B2(new_n1316), .ZN(new_n1343));
  OR3_X1    g1143(.A1(new_n1320), .A2(KEYINPUT123), .A3(new_n1321), .ZN(new_n1344));
  OAI21_X1  g1144(.A(KEYINPUT123), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1344), .A2(new_n1342), .A3(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1347), .A2(KEYINPUT61), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1338), .A2(KEYINPUT63), .A3(new_n1333), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1343), .A2(new_n1346), .A3(new_n1348), .A4(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1340), .A2(new_n1350), .ZN(G405));
  INV_X1    g1151(.A(KEYINPUT127), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1329), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1272), .A2(KEYINPUT121), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1354), .A2(new_n1246), .A3(new_n1236), .ZN(new_n1355));
  AOI21_X1  g1155(.A(G378), .B1(new_n1355), .B2(new_n1225), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1352), .B1(new_n1353), .B2(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(G375), .A2(new_n1275), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1358), .A2(KEYINPUT127), .A3(new_n1329), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1357), .A2(new_n1316), .A3(new_n1359), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1316), .B1(new_n1357), .B2(new_n1359), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1347), .B1(new_n1360), .B2(new_n1361), .ZN(new_n1362));
  NOR3_X1   g1162(.A1(new_n1353), .A2(new_n1356), .A3(new_n1352), .ZN(new_n1363));
  AOI21_X1  g1163(.A(KEYINPUT127), .B1(new_n1358), .B2(new_n1329), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1333), .B1(new_n1363), .B2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1347), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1357), .A2(new_n1316), .A3(new_n1359), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1365), .A2(new_n1366), .A3(new_n1367), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1362), .A2(new_n1368), .ZN(G402));
endmodule


