//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G119), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT74), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n191), .B1(G119), .B2(new_n188), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT24), .B(G110), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT75), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  OR2_X1    g009(.A1(new_n195), .A2(KEYINPUT76), .ZN(new_n196));
  XNOR2_X1  g010(.A(G125), .B(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT16), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  OR3_X1    g013(.A1(new_n199), .A2(KEYINPUT16), .A3(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(G146), .A3(new_n200), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT23), .B1(new_n188), .B2(G119), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT77), .A3(new_n189), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT77), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n207), .B1(new_n189), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G110), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n195), .A2(KEYINPUT76), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n196), .A2(new_n205), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT22), .B(G137), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n214), .B(KEYINPUT78), .ZN(new_n215));
  INV_X1    g029(.A(G953), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n216), .A2(G221), .A3(G234), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n215), .B(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT64), .B(G146), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n197), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n192), .A2(new_n194), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n210), .A2(G110), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n204), .B(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n213), .A2(new_n219), .A3(new_n225), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n218), .A2(KEYINPUT79), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n218), .A2(KEYINPUT79), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n213), .A2(new_n225), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n187), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT25), .ZN(new_n231));
  INV_X1    g045(.A(G217), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n232), .B1(G234), .B2(new_n187), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n234), .B(new_n187), .C1(new_n226), .C2(new_n229), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n231), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT80), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n231), .A2(KEYINPUT80), .A3(new_n233), .A4(new_n235), .ZN(new_n239));
  OR2_X1    g053(.A1(new_n226), .A2(new_n229), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n233), .A2(G902), .ZN(new_n241));
  XOR2_X1   g055(.A(new_n241), .B(KEYINPUT81), .Z(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n238), .A2(new_n239), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n244), .B(KEYINPUT82), .ZN(new_n245));
  INV_X1    g059(.A(G469), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n221), .A2(G143), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT1), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n202), .A2(G143), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n247), .A2(new_n248), .A3(G128), .A4(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n220), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(new_n249), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n202), .A2(G143), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n188), .B1(new_n255), .B2(KEYINPUT1), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n251), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT84), .ZN(new_n258));
  INV_X1    g072(.A(G104), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n258), .A2(KEYINPUT3), .B1(new_n259), .B2(G107), .ZN(new_n260));
  OAI22_X1  g074(.A1(new_n258), .A2(KEYINPUT3), .B1(new_n259), .B2(G107), .ZN(new_n261));
  INV_X1    g075(.A(G101), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT3), .ZN(new_n263));
  INV_X1    g077(.A(G107), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT84), .A4(G104), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n260), .A2(new_n261), .A3(new_n262), .A4(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT85), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n264), .A2(G104), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n259), .A2(G107), .ZN(new_n270));
  OAI21_X1  g084(.A(G101), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n257), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT86), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n266), .A2(new_n267), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n266), .A2(new_n267), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT86), .A3(new_n257), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT1), .B1(new_n220), .B2(new_n252), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n220), .A2(new_n252), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n280), .A2(G128), .B1(new_n281), .B2(new_n255), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n248), .A2(G128), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n253), .A2(new_n249), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n274), .A2(new_n279), .B1(new_n285), .B2(new_n277), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT12), .ZN(new_n287));
  INV_X1    g101(.A(G137), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n288), .A2(KEYINPUT65), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(KEYINPUT65), .ZN(new_n290));
  OAI211_X1 g104(.A(KEYINPUT11), .B(G134), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G131), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT11), .B1(new_n288), .B2(G134), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n288), .A2(G134), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n291), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n292), .B1(new_n291), .B2(new_n295), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n286), .A2(new_n287), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n287), .B1(new_n286), .B2(new_n299), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n274), .A2(new_n279), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT10), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n260), .A2(new_n261), .A3(new_n265), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G101), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n268), .A2(KEYINPUT4), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n281), .A2(new_n255), .ZN(new_n310));
  NAND2_X1  g124(.A1(KEYINPUT0), .A2(G128), .ZN(new_n311));
  OR2_X1    g125(.A1(KEYINPUT0), .A2(G128), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n247), .A2(KEYINPUT0), .A3(G128), .A4(new_n250), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n308), .A2(KEYINPUT4), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n309), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT87), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n277), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT87), .B1(new_n268), .B2(new_n271), .ZN(new_n320));
  OAI221_X1 g134(.A(KEYINPUT10), .B1(new_n282), .B2(new_n284), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n299), .B(KEYINPUT88), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n306), .A2(new_n317), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  XOR2_X1   g137(.A(G110), .B(G140), .Z(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT83), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n216), .A2(G227), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n325), .B(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n303), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n306), .A2(new_n317), .A3(new_n321), .ZN(new_n330));
  INV_X1    g144(.A(new_n299), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n327), .B1(new_n332), .B2(new_n323), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n246), .B(new_n187), .C1(new_n329), .C2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n323), .A3(new_n327), .ZN(new_n335));
  INV_X1    g149(.A(new_n330), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n301), .A2(new_n302), .B1(new_n336), .B2(new_n322), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n335), .B(G469), .C1(new_n337), .C2(new_n327), .ZN(new_n338));
  NAND2_X1  g152(.A1(G469), .A2(G902), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n334), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G221), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT9), .B(G234), .Z(new_n342));
  AOI21_X1  g156(.A(new_n341), .B1(new_n342), .B2(new_n187), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n245), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(KEYINPUT2), .A2(G113), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT66), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT2), .ZN(new_n351));
  INV_X1    g165(.A(G113), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n349), .A2(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G119), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G116), .ZN(new_n355));
  INV_X1    g169(.A(G116), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G119), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT67), .ZN(new_n359));
  XNOR2_X1  g173(.A(G116), .B(G119), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT67), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n353), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n349), .A2(new_n350), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n351), .A2(new_n352), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(new_n358), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT68), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n358), .A2(KEYINPUT67), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n360), .A2(new_n361), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT68), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n353), .A2(new_n360), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT65), .B(G137), .Z(new_n376));
  OAI21_X1  g190(.A(new_n294), .B1(new_n376), .B2(G134), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G131), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n296), .B(new_n378), .C1(new_n282), .C2(new_n284), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n313), .B(new_n314), .C1(new_n297), .C2(new_n298), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n375), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT28), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(G101), .ZN(new_n385));
  NOR2_X1   g199(.A1(G237), .A2(G953), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G210), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n385), .B(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n381), .A2(KEYINPUT69), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT69), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n375), .A2(new_n379), .A3(new_n380), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n371), .A2(new_n373), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n380), .A2(new_n379), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n389), .A2(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n383), .B(new_n388), .C1(new_n394), .C2(new_n382), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n389), .A2(new_n391), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT30), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n380), .A2(new_n379), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n380), .B2(new_n379), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n392), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n388), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n395), .A2(new_n396), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT71), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n375), .B1(new_n380), .B2(new_n379), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(KEYINPUT72), .ZN(new_n409));
  INV_X1    g223(.A(new_n397), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT28), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n411), .A2(KEYINPUT29), .A3(new_n383), .A4(new_n388), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n395), .A2(KEYINPUT71), .A3(new_n396), .A4(new_n404), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n407), .A2(new_n187), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G472), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT32), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n397), .A2(new_n401), .A3(new_n388), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT31), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n397), .A2(new_n401), .A3(KEYINPUT31), .A4(new_n388), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n383), .B1(new_n394), .B2(new_n382), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n403), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n421), .A2(new_n423), .A3(KEYINPUT70), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT70), .B1(new_n421), .B2(new_n423), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(G472), .A2(G902), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n416), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n427), .ZN(new_n429));
  NOR4_X1   g243(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT32), .A4(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n415), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT73), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT73), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n433), .B(new_n415), .C1(new_n428), .C2(new_n430), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n346), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT96), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n386), .A2(KEYINPUT91), .A3(new_n252), .A4(G214), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT91), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G143), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n252), .A2(KEYINPUT91), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G214), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n442), .A2(G237), .A3(G953), .ZN(new_n443));
  OAI211_X1 g257(.A(G131), .B(new_n437), .C1(new_n441), .C2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT18), .ZN(new_n445));
  OR2_X1    g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n386), .A2(G214), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n439), .A3(new_n440), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n437), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n445), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n222), .B1(new_n202), .B2(new_n197), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n292), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n446), .A2(new_n450), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT92), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n444), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n448), .A2(KEYINPUT92), .A3(G131), .A4(new_n437), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(KEYINPUT17), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT94), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT94), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n456), .A2(new_n460), .A3(KEYINPUT17), .A4(new_n457), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n205), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT95), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT95), .ZN(new_n465));
  AOI211_X1 g279(.A(new_n465), .B(new_n205), .C1(new_n459), .C2(new_n461), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n456), .A2(new_n457), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n452), .ZN(new_n469));
  OR2_X1    g283(.A1(new_n469), .A2(KEYINPUT17), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n454), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(G113), .B(G122), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(new_n259), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n436), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n462), .A2(new_n463), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n465), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n462), .A2(KEYINPUT95), .A3(new_n463), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n470), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n478), .A2(new_n436), .A3(new_n473), .A4(new_n453), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n473), .B1(new_n478), .B2(new_n453), .ZN(new_n482));
  OAI211_X1 g296(.A(KEYINPUT98), .B(new_n187), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT98), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n478), .A2(new_n473), .A3(new_n453), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT96), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n482), .B1(new_n486), .B2(new_n479), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n484), .B1(new_n487), .B2(G902), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n483), .A2(G475), .A3(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(G475), .A2(G902), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT97), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n486), .A2(new_n479), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n197), .B(KEYINPUT19), .Z(new_n493));
  OAI211_X1 g307(.A(new_n469), .B(new_n204), .C1(new_n220), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n453), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT93), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n473), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n494), .A2(KEYINPUT93), .A3(new_n453), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n491), .B1(new_n492), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n500), .ZN(new_n502));
  AOI211_X1 g316(.A(KEYINPUT97), .B(new_n502), .C1(new_n486), .C2(new_n479), .ZN(new_n503));
  OAI211_X1 g317(.A(KEYINPUT20), .B(new_n490), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n492), .A2(new_n500), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n490), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n489), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT99), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n356), .A2(G122), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT14), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT101), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n356), .A2(G122), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(new_n511), .B2(KEYINPUT14), .ZN(new_n515));
  OAI21_X1  g329(.A(G107), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n511), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n516), .B1(G107), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n252), .A2(G128), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT100), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n188), .A2(G143), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G134), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT13), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n523), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n522), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n517), .B(new_n264), .ZN(new_n528));
  OAI22_X1  g342(.A1(new_n518), .A2(new_n524), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n342), .A2(G217), .A3(new_n216), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n187), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(KEYINPUT102), .ZN(new_n533));
  INV_X1    g347(.A(G478), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(KEYINPUT15), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n532), .A2(new_n535), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n216), .A2(G952), .ZN(new_n540));
  NAND2_X1  g354(.A1(G234), .A2(G237), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  XOR2_X1   g357(.A(KEYINPUT21), .B(G898), .Z(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n541), .A2(G902), .A3(G953), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n543), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT99), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n489), .A2(new_n504), .A3(new_n550), .A4(new_n508), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n510), .A2(new_n539), .A3(new_n549), .A4(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(G214), .B1(G237), .B2(G902), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n315), .A2(G125), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(G125), .B2(new_n285), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n216), .A2(G224), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT6), .ZN(new_n559));
  XOR2_X1   g373(.A(G110), .B(G122), .Z(new_n560));
  XOR2_X1   g374(.A(new_n560), .B(KEYINPUT89), .Z(new_n561));
  AND3_X1   g375(.A1(new_n309), .A2(new_n392), .A3(new_n316), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n359), .A2(new_n362), .A3(KEYINPUT5), .ZN(new_n563));
  OAI21_X1  g377(.A(G113), .B1(new_n355), .B2(KEYINPUT5), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n367), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n277), .A2(new_n318), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n268), .A2(KEYINPUT87), .A3(new_n271), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n561), .B1(new_n562), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n566), .B1(new_n319), .B2(new_n320), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n309), .A2(new_n392), .A3(new_n316), .ZN(new_n573));
  INV_X1    g387(.A(new_n560), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n559), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n573), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT6), .B1(new_n577), .B2(new_n561), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n558), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT90), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(KEYINPUT90), .B(new_n558), .C1(new_n576), .C2(new_n578), .ZN(new_n582));
  AOI21_X1  g396(.A(G902), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n557), .A2(KEYINPUT7), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n556), .B(new_n584), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n360), .A2(KEYINPUT5), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n373), .B1(new_n586), .B2(new_n564), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n278), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n560), .B(KEYINPUT8), .Z(new_n589));
  OAI211_X1 g403(.A(new_n588), .B(new_n589), .C1(new_n278), .C2(new_n567), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n585), .A2(new_n575), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(G210), .B1(G237), .B2(G902), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n583), .A2(new_n593), .A3(new_n591), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n554), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n435), .A2(new_n552), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(new_n262), .ZN(G3));
  NAND2_X1  g414(.A1(new_n426), .A2(new_n427), .ZN(new_n601));
  INV_X1    g415(.A(G472), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n424), .A2(new_n425), .A3(G902), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n346), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n531), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT103), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT104), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n529), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(new_n530), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT33), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n534), .A2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n533), .A2(new_n534), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n583), .A2(new_n593), .A3(new_n591), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n593), .B1(new_n583), .B2(new_n591), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n553), .B(new_n549), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  AOI211_X1 g436(.A(new_n619), .B(new_n622), .C1(new_n510), .C2(new_n551), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n607), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT34), .B(G104), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  INV_X1    g440(.A(new_n622), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n501), .A2(new_n503), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n490), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n507), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n489), .A2(new_n504), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n627), .A2(new_n631), .A3(new_n538), .A4(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n606), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT35), .B(G107), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NOR3_X1   g450(.A1(new_n552), .A2(new_n598), .A3(new_n604), .ZN(new_n637));
  INV_X1    g451(.A(new_n345), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT36), .B1(new_n227), .B2(new_n228), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n213), .A2(new_n225), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n242), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n238), .A2(new_n239), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n637), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT105), .B(KEYINPUT37), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G110), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n644), .B(new_n646), .ZN(G12));
  NAND2_X1  g461(.A1(new_n432), .A2(new_n434), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n638), .A2(new_n597), .A3(new_n643), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n543), .B1(new_n547), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n631), .A2(new_n632), .A3(new_n538), .A4(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  AOI21_X1  g471(.A(new_n539), .B1(new_n510), .B2(new_n551), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n658), .A2(new_n553), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n660));
  INV_X1    g474(.A(new_n643), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n595), .A2(new_n596), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT38), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n428), .A2(new_n430), .ZN(new_n667));
  INV_X1    g481(.A(new_n417), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n403), .B1(new_n409), .B2(new_n410), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n671), .B1(new_n670), .B2(new_n669), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n187), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G472), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n662), .A2(new_n666), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n660), .B1(new_n659), .B2(new_n661), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n652), .B(KEYINPUT39), .Z(new_n678));
  NAND2_X1  g492(.A1(new_n638), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT40), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n676), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n252), .ZN(G45));
  NAND2_X1  g496(.A1(new_n510), .A2(new_n551), .ZN(new_n683));
  INV_X1    g497(.A(new_n619), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n684), .A3(new_n653), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n619), .B1(new_n510), .B2(new_n551), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(KEYINPUT109), .A3(new_n653), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n687), .A2(new_n650), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  INV_X1    g505(.A(KEYINPUT110), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n688), .A2(new_n627), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n332), .A2(new_n323), .ZN(new_n694));
  OAI22_X1  g508(.A1(new_n694), .A2(new_n327), .B1(new_n303), .B2(new_n328), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n246), .B1(new_n695), .B2(new_n187), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n344), .A3(new_n334), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n245), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n432), .A2(new_n699), .A3(new_n700), .A4(new_n434), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n692), .B1(new_n693), .B2(new_n701), .ZN(new_n702));
  AND4_X1   g516(.A1(new_n432), .A2(new_n699), .A3(new_n434), .A4(new_n700), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n623), .A3(KEYINPUT110), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT41), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G113), .ZN(G15));
  NOR2_X1   g521(.A1(new_n701), .A2(new_n633), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n356), .ZN(G18));
  NAND3_X1  g523(.A1(new_n432), .A2(new_n434), .A3(new_n643), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n699), .A2(new_n597), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n710), .A2(new_n552), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n354), .ZN(G21));
  INV_X1    g527(.A(new_n244), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n388), .B1(new_n411), .B2(new_n383), .ZN(new_n715));
  INV_X1    g529(.A(new_n421), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n427), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT111), .B(G472), .Z(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n714), .B(new_n717), .C1(new_n603), .C2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n698), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n658), .A2(new_n627), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT112), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n658), .A2(new_n724), .A3(new_n627), .A4(new_n721), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  INV_X1    g541(.A(new_n711), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n643), .B(new_n717), .C1(new_n603), .C2(new_n719), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT113), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n687), .A2(new_n689), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  AND3_X1   g546(.A1(new_n688), .A2(KEYINPUT109), .A3(new_n653), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT109), .B1(new_n688), .B2(new_n653), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n663), .A2(new_n554), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n346), .A2(new_n432), .A3(new_n434), .A4(new_n735), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n345), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n687), .A2(new_n689), .A3(new_n735), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n431), .A2(new_n714), .ZN(new_n741));
  OAI22_X1  g555(.A1(new_n737), .A2(KEYINPUT42), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  INV_X1    g557(.A(new_n736), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT114), .B1(new_n744), .B2(new_n655), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n736), .A2(new_n746), .A3(new_n654), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n523), .ZN(G36));
  NAND3_X1  g563(.A1(new_n510), .A2(new_n551), .A3(new_n684), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n604), .A3(new_n643), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n752), .A2(KEYINPUT44), .A3(new_n604), .A4(new_n643), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n735), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n335), .B1(new_n337), .B2(new_n327), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n335), .B(KEYINPUT45), .C1(new_n337), .C2(new_n327), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(G469), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(KEYINPUT46), .A3(new_n339), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n334), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n764), .A2(new_n339), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT46), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n765), .A2(KEYINPUT115), .A3(new_n334), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n768), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n773), .A2(new_n344), .A3(new_n678), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n755), .A2(KEYINPUT116), .A3(new_n735), .A4(new_n756), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n759), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G137), .ZN(G39));
  INV_X1    g591(.A(KEYINPUT47), .ZN(new_n778));
  INV_X1    g592(.A(new_n773), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n778), .B1(new_n779), .B2(new_n343), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n773), .A2(KEYINPUT47), .A3(new_n344), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n687), .A2(new_n689), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n783), .A2(new_n554), .A3(new_n663), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n782), .A2(new_n784), .A3(new_n648), .A4(new_n245), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  NAND2_X1  g600(.A1(new_n697), .A2(new_n334), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n787), .B(KEYINPUT117), .Z(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n343), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n780), .A2(new_n781), .A3(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n752), .A2(new_n543), .ZN(new_n791));
  INV_X1    g605(.A(new_n720), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n790), .A2(new_n791), .A3(new_n792), .A4(new_n735), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n699), .A2(new_n735), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n791), .A2(new_n730), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n675), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n795), .A2(new_n700), .A3(new_n543), .A4(new_n797), .ZN(new_n798));
  OR3_X1    g612(.A1(new_n798), .A2(new_n683), .A3(new_n684), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n793), .A2(new_n796), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n666), .A2(new_n553), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n791), .A2(new_n801), .A3(new_n721), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n800), .A2(KEYINPUT51), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n802), .B(KEYINPUT50), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n793), .A2(new_n796), .A3(new_n799), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n688), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n798), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n805), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT118), .B1(new_n683), .B2(new_n539), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n810), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n688), .A2(KEYINPUT118), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n622), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n599), .B1(new_n816), .B2(new_n607), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n712), .B1(new_n702), .B2(new_n704), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n708), .B1(new_n723), .B2(new_n725), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n817), .A2(new_n644), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n748), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n742), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n687), .A2(new_n689), .A3(new_n730), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n631), .A2(new_n504), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n489), .A2(new_n539), .A3(new_n643), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n648), .A2(new_n825), .A3(new_n652), .A4(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n638), .B(new_n735), .C1(new_n824), .C2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n829), .B1(new_n643), .B2(new_n652), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n661), .A2(KEYINPUT119), .A3(new_n653), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n638), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n797), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n659), .A2(new_n663), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n731), .A2(new_n690), .A3(new_n656), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n823), .A2(KEYINPUT53), .A3(new_n828), .A4(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n733), .A2(new_n734), .ZN(new_n840));
  INV_X1    g654(.A(new_n741), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n735), .A3(new_n841), .A4(new_n739), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n738), .B1(new_n783), .B2(new_n736), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n748), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n818), .A2(new_n644), .A3(new_n819), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n844), .A2(new_n845), .A3(new_n817), .A4(new_n828), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n835), .B(KEYINPUT52), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n839), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n838), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n838), .A2(new_n848), .A3(KEYINPUT54), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n812), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n791), .A2(new_n597), .A3(new_n721), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n741), .B1(new_n855), .B2(KEYINPUT48), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n791), .A2(new_n795), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n855), .A2(KEYINPUT48), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n857), .B(new_n858), .Z(new_n859));
  NAND4_X1  g673(.A1(new_n853), .A2(KEYINPUT120), .A3(new_n854), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(G953), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n853), .A2(new_n862), .A3(new_n854), .A4(new_n859), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n540), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n788), .B(KEYINPUT49), .Z(new_n865));
  NOR3_X1   g679(.A1(new_n865), .A2(new_n675), .A3(new_n750), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n666), .A2(new_n343), .A3(new_n554), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n714), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n861), .A2(new_n864), .A3(new_n868), .ZN(G75));
  OR2_X1    g683(.A1(new_n576), .A2(new_n578), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(new_n558), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT122), .Z(new_n872));
  AOI21_X1  g686(.A(new_n187), .B1(new_n838), .B2(new_n848), .ZN(new_n873));
  AOI211_X1 g687(.A(KEYINPUT55), .B(KEYINPUT56), .C1(new_n873), .C2(G210), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT55), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n849), .A2(G210), .A3(G902), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n872), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n216), .A2(G952), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(G210), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n882), .B(new_n187), .C1(new_n838), .C2(new_n848), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT55), .B1(new_n883), .B2(KEYINPUT56), .ZN(new_n884));
  INV_X1    g698(.A(new_n872), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n876), .A2(new_n875), .A3(new_n877), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n879), .A2(new_n881), .A3(new_n887), .ZN(G51));
  XOR2_X1   g702(.A(new_n339), .B(KEYINPUT57), .Z(new_n889));
  NAND3_X1  g703(.A1(new_n851), .A2(new_n852), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n695), .ZN(new_n891));
  INV_X1    g705(.A(new_n764), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n873), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n880), .B1(new_n891), .B2(new_n893), .ZN(G54));
  NAND2_X1  g708(.A1(KEYINPUT58), .A2(G475), .ZN(new_n895));
  AOI211_X1 g709(.A(new_n187), .B(new_n895), .C1(new_n838), .C2(new_n848), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n880), .B1(new_n896), .B2(new_n628), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n898));
  INV_X1    g712(.A(new_n895), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n898), .B(new_n628), .C1(new_n873), .C2(new_n899), .ZN(new_n900));
  AND4_X1   g714(.A1(new_n844), .A2(new_n845), .A3(new_n817), .A4(new_n828), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT53), .B1(new_n901), .B2(new_n837), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n846), .A2(new_n847), .A3(new_n839), .ZN(new_n903));
  OAI211_X1 g717(.A(G902), .B(new_n899), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT123), .B1(new_n904), .B2(new_n629), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n897), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g722(.A(KEYINPUT124), .B(new_n897), .C1(new_n900), .C2(new_n905), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(G60));
  NAND2_X1  g724(.A1(G478), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT59), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n851), .A2(new_n852), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n615), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(new_n880), .ZN(G63));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT60), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n838), .B2(new_n848), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n920), .A2(new_n240), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n641), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n881), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(G66));
  AOI21_X1  g739(.A(new_n216), .B1(new_n544), .B2(G224), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n820), .B2(new_n216), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT125), .Z(new_n928));
  INV_X1    g742(.A(G898), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n870), .B1(new_n929), .B2(G953), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n928), .B(new_n930), .ZN(G69));
  NAND2_X1  g745(.A1(G227), .A2(G900), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n216), .A2(G900), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n731), .A2(new_n656), .A3(new_n690), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n774), .A2(new_n841), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n659), .A2(new_n663), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n776), .A2(new_n937), .A3(new_n785), .A4(new_n844), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n933), .B1(new_n938), .B2(new_n216), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n399), .A2(new_n400), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n493), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  OAI211_X1 g758(.A(G953), .B(new_n932), .C1(new_n941), .C2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n939), .A2(new_n940), .ZN(new_n946));
  AOI211_X1 g760(.A(KEYINPUT126), .B(new_n933), .C1(new_n938), .C2(new_n216), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n932), .A2(G953), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n681), .A2(new_n934), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n814), .A2(new_n815), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n952), .A2(new_n678), .A3(new_n744), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n951), .A2(new_n776), .A3(new_n785), .A4(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n944), .B1(new_n955), .B2(G953), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n948), .A2(new_n949), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n945), .A2(new_n957), .ZN(G72));
  NAND2_X1  g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT63), .Z(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n954), .B2(new_n820), .ZN(new_n961));
  INV_X1    g775(.A(new_n402), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n403), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n880), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n960), .B1(new_n938), .B2(new_n820), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n965), .A2(new_n403), .A3(new_n962), .ZN(new_n966));
  INV_X1    g780(.A(new_n404), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n960), .B1(new_n967), .B2(new_n668), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n849), .A2(KEYINPUT127), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT127), .B1(new_n849), .B2(new_n969), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n964), .B(new_n966), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(G57));
endmodule


