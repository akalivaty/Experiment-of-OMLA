//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n627, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1237, new_n1238;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G221), .A4(G218), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT68), .Z(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n471), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n462), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n471), .A2(G136), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n484));
  INV_X1    g059(.A(new_n470), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  OAI211_X1 g061(.A(G126), .B(G2105), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n484), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n487), .A2(new_n489), .A3(new_n484), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n461), .C1(new_n485), .C2(new_n486), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n471), .A2(new_n495), .A3(G138), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n491), .A2(new_n492), .B1(new_n494), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n501), .A2(new_n503), .B1(new_n500), .B2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G62), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(KEYINPUT71), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n504), .A2(new_n507), .A3(G62), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n498), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n502), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n501), .A2(new_n503), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n500), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(new_n511), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n513), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n509), .A2(new_n519), .ZN(G166));
  XNOR2_X1  g095(.A(KEYINPUT72), .B(G89), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n504), .A2(new_n516), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  OAI211_X1 g104(.A(G51), .B(G543), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n514), .A2(G63), .A3(G651), .A4(new_n515), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n522), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n522), .A2(new_n531), .A3(KEYINPUT73), .A4(new_n532), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(G168));
  NAND2_X1  g112(.A1(new_n512), .A2(G52), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n504), .A2(G90), .A3(new_n516), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n538), .B(new_n539), .C1(new_n540), .C2(new_n498), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  NAND2_X1  g117(.A1(new_n504), .A2(G56), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n498), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT74), .B(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n512), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n517), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n552));
  XOR2_X1   g127(.A(new_n552), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(G78), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT77), .B1(new_n557), .B2(new_n502), .ZN(new_n558));
  OR3_X1    g133(.A1(new_n557), .A2(new_n502), .A3(KEYINPUT77), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n514), .A2(new_n515), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n558), .B(new_n559), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n516), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n512), .A2(new_n566), .A3(G53), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n562), .A2(G651), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n517), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n504), .A2(KEYINPUT76), .A3(new_n516), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n570), .A2(G91), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G168), .ZN(G286));
  INV_X1    g149(.A(G166), .ZN(G303));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  INV_X1    g151(.A(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n563), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n512), .A2(KEYINPUT78), .A3(G49), .ZN(new_n579));
  INV_X1    g154(.A(G74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n560), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n578), .A2(new_n579), .B1(new_n581), .B2(G651), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n570), .A2(G87), .A3(new_n571), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n560), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(G48), .B2(new_n512), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n570), .A2(new_n571), .ZN(new_n589));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n498), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n512), .A2(G47), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n517), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n570), .A2(G92), .A3(new_n571), .ZN(new_n600));
  XOR2_X1   g175(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n570), .A2(G92), .A3(new_n571), .A4(new_n601), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n512), .A2(G54), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n502), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT70), .B1(new_n502), .B2(KEYINPUT5), .ZN(new_n608));
  OAI211_X1 g183(.A(G66), .B(new_n515), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n609), .A2(KEYINPUT80), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G651), .ZN(new_n612));
  AOI21_X1  g187(.A(KEYINPUT80), .B1(new_n609), .B2(new_n610), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT81), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n609), .A2(new_n610), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n618), .A2(G651), .A3(new_n611), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT81), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n619), .A2(new_n620), .A3(new_n606), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n605), .B1(new_n615), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n599), .B1(new_n622), .B2(G868), .ZN(G284));
  XNOR2_X1  g198(.A(G284), .B(KEYINPUT82), .ZN(G321));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NOR2_X1   g200(.A1(G168), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g201(.A1(new_n626), .A2(KEYINPUT83), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n626), .A2(KEYINPUT83), .ZN(new_n628));
  NAND2_X1  g203(.A1(G299), .A2(new_n625), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(G297));
  AOI21_X1  g205(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n622), .B1(new_n632), .B2(G860), .ZN(G148));
  INV_X1    g208(.A(KEYINPUT84), .ZN(new_n634));
  INV_X1    g209(.A(new_n605), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n614), .A2(KEYINPUT81), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n620), .B1(new_n619), .B2(new_n606), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n634), .B1(new_n638), .B2(G559), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n622), .A2(KEYINPUT84), .A3(new_n632), .ZN(new_n640));
  AND3_X1   g215(.A1(new_n639), .A2(G868), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n625), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g218(.A1(new_n462), .A2(new_n472), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  INV_X1    g221(.A(G2100), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n471), .A2(G135), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n461), .A2(G111), .ZN(new_n651));
  OAI21_X1  g226(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n652));
  INV_X1    g227(.A(G123), .ZN(new_n653));
  OAI221_X1 g228(.A(new_n650), .B1(new_n651), .B2(new_n652), .C1(new_n653), .C2(new_n476), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  NAND3_X1  g230(.A1(new_n648), .A2(new_n649), .A3(new_n655), .ZN(G156));
  XNOR2_X1  g231(.A(KEYINPUT15), .B(G2435), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT87), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT86), .B(G2438), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2427), .B(G2430), .Z(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT85), .B(KEYINPUT14), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2451), .B(G2454), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1341), .B(G1348), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n665), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2443), .B(G2446), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  AND3_X1   g248(.A1(new_n672), .A2(G14), .A3(new_n673), .ZN(G401));
  NOR2_X1   g249(.A1(G2072), .A2(G2078), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n442), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT18), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n676), .B(KEYINPUT17), .ZN(new_n682));
  INV_X1    g257(.A(new_n678), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n683), .A2(new_n679), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n681), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n679), .B1(new_n677), .B2(KEYINPUT88), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(KEYINPUT88), .B2(new_n677), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n687), .A2(KEYINPUT89), .A3(new_n683), .ZN(new_n688));
  INV_X1    g263(.A(new_n679), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(new_n682), .ZN(new_n690));
  AOI21_X1  g265(.A(KEYINPUT89), .B1(new_n687), .B2(new_n683), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n685), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G2096), .B(G2100), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G227));
  XOR2_X1   g269(.A(G1971), .B(G1976), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT19), .ZN(new_n696));
  XOR2_X1   g271(.A(G1956), .B(G2474), .Z(new_n697));
  XOR2_X1   g272(.A(G1961), .B(G1966), .Z(new_n698));
  AND2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT20), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n697), .A2(new_n698), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n696), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n696), .B2(new_n702), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1991), .B(G1996), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1981), .B(G1986), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(G229));
  XNOR2_X1  g286(.A(KEYINPUT31), .B(G11), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT103), .B(G28), .Z(new_n713));
  AOI21_X1  g288(.A(G29), .B1(new_n713), .B2(KEYINPUT30), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(KEYINPUT30), .B2(new_n713), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n712), .B(new_n715), .C1(new_n654), .C2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT26), .Z(new_n719));
  INV_X1    g294(.A(G129), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n476), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n472), .A2(G105), .ZN(new_n722));
  INV_X1    g297(.A(new_n471), .ZN(new_n723));
  INV_X1    g298(.A(G141), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(new_n716), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n716), .B2(G32), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT27), .B(G1996), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n717), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G29), .A2(G33), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT100), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n462), .A2(G127), .ZN(new_n734));
  AND2_X1   g309(.A1(G115), .A2(G2104), .ZN(new_n735));
  OAI21_X1  g310(.A(G2105), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT25), .ZN(new_n737));
  NAND2_X1  g312(.A1(G103), .A2(G2104), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G2105), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n471), .A2(G139), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n733), .B1(new_n743), .B2(new_n716), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G2072), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n731), .B(new_n745), .C1(new_n729), .C2(new_n730), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n550), .A2(G16), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G16), .B2(G19), .ZN(new_n748));
  INV_X1    g323(.A(G1341), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n716), .A2(G35), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G162), .B2(new_n716), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT29), .Z(new_n753));
  INV_X1    g328(.A(G2090), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n746), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G34), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n757), .A2(KEYINPUT24), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(KEYINPUT24), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n716), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G160), .B2(new_n716), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT101), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2084), .ZN(new_n763));
  INV_X1    g338(.A(G16), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n764), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n756), .B(new_n763), .C1(G1966), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n716), .A2(G27), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G164), .B2(new_n716), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n753), .A2(new_n754), .B1(G2078), .B2(new_n769), .ZN(new_n770));
  OAI221_X1 g345(.A(new_n770), .B1(new_n749), .B2(new_n748), .C1(G2078), .C2(new_n769), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n766), .A2(G1966), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT102), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n471), .A2(G140), .ZN(new_n774));
  NOR2_X1   g349(.A1(G104), .A2(G2105), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT97), .ZN(new_n776));
  OAI21_X1  g351(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n777));
  AND3_X1   g352(.A1(new_n477), .A2(KEYINPUT96), .A3(G128), .ZN(new_n778));
  AOI21_X1  g353(.A(KEYINPUT96), .B1(new_n477), .B2(G128), .ZN(new_n779));
  OAI221_X1 g354(.A(new_n774), .B1(new_n776), .B2(new_n777), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G29), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT98), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n716), .A2(G26), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT99), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT28), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2067), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n767), .A2(new_n771), .A3(new_n773), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n764), .A2(G5), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G171), .B2(new_n764), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT104), .Z(new_n791));
  AND2_X1   g366(.A1(new_n791), .A2(G1961), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(G1961), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n764), .A2(G20), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT23), .Z(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G299), .B2(G16), .ZN(new_n796));
  INV_X1    g371(.A(G1956), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n792), .A2(new_n793), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n764), .A2(G4), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n622), .B2(new_n764), .ZN(new_n801));
  INV_X1    g376(.A(G1348), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n788), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n764), .A2(G24), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n597), .B2(new_n764), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(G1986), .Z(new_n807));
  INV_X1    g382(.A(G25), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n808), .A2(KEYINPUT90), .A3(G29), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT90), .B1(new_n808), .B2(G29), .ZN(new_n810));
  OR2_X1    g385(.A1(G95), .A2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n811), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT91), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n471), .A2(G131), .ZN(new_n814));
  INV_X1    g389(.A(G119), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(new_n476), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n809), .B(new_n810), .C1(new_n817), .C2(new_n716), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT35), .B(G1991), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n807), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT94), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT32), .B(G1981), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(G305), .A2(G16), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT92), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n764), .A2(G6), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n826), .B1(new_n825), .B2(new_n828), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n824), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n831), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n833), .A2(new_n829), .A3(new_n823), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n764), .A2(G22), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G166), .B2(new_n764), .ZN(new_n837));
  INV_X1    g412(.A(G1971), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(G16), .A2(G23), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT93), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n578), .A2(new_n579), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n581), .A2(G651), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n570), .A2(G87), .A3(new_n571), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n582), .A2(KEYINPUT93), .A3(new_n583), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n841), .B1(new_n849), .B2(new_n764), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT33), .B(G1976), .Z(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n852), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n839), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n822), .B1(new_n835), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n839), .A2(new_n854), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n832), .A2(new_n834), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n857), .A2(KEYINPUT94), .A3(new_n858), .A4(new_n853), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT34), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n821), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n856), .A2(new_n859), .A3(KEYINPUT34), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(KEYINPUT95), .A2(KEYINPUT36), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n862), .A2(new_n865), .A3(new_n863), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n804), .B1(new_n867), .B2(new_n868), .ZN(G311));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n868), .ZN(new_n870));
  INV_X1    g445(.A(new_n804), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(G150));
  NAND3_X1  g447(.A1(new_n504), .A2(G93), .A3(new_n516), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n512), .A2(G55), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n514), .A2(G67), .A3(new_n515), .ZN(new_n876));
  NAND2_X1  g451(.A1(G80), .A2(G543), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(G651), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n875), .A2(new_n879), .A3(KEYINPUT106), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n873), .A2(new_n874), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n498), .B1(new_n876), .B2(new_n877), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(G860), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT37), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n622), .A2(G559), .ZN(new_n888));
  XNOR2_X1  g463(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n550), .B1(new_n880), .B2(new_n884), .ZN(new_n891));
  NOR4_X1   g466(.A1(new_n545), .A2(new_n549), .A3(new_n882), .A4(new_n883), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n890), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT39), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT107), .ZN(new_n896));
  INV_X1    g471(.A(G860), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n894), .B2(KEYINPUT39), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n887), .B1(new_n896), .B2(new_n898), .ZN(G145));
  NAND2_X1  g474(.A1(new_n496), .A2(new_n494), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n487), .A2(new_n489), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n726), .B(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n780), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n742), .A2(KEYINPUT108), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n817), .B(new_n645), .ZN(new_n908));
  INV_X1    g483(.A(G130), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n461), .A2(G118), .ZN(new_n910));
  OAI21_X1  g485(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n911));
  OAI22_X1  g486(.A1(new_n476), .A2(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n912), .B1(G142), .B2(new_n471), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n908), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n742), .A2(KEYINPUT108), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n905), .A2(new_n906), .A3(new_n915), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n907), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT110), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n474), .B(new_n654), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(new_n482), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n907), .A2(new_n916), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n914), .A2(KEYINPUT110), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n914), .B1(new_n907), .B2(new_n916), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n920), .B1(new_n917), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(KEYINPUT109), .B(G37), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g504(.A(KEYINPUT111), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT42), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n930), .A2(KEYINPUT42), .ZN(new_n932));
  XNOR2_X1  g507(.A(G166), .B(new_n597), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n849), .B(new_n588), .C1(new_n590), .C2(new_n589), .ZN(new_n934));
  INV_X1    g509(.A(new_n848), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT93), .B1(new_n582), .B2(new_n583), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(G305), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n933), .A2(new_n934), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(G166), .A2(G290), .ZN(new_n940));
  NAND2_X1  g515(.A1(G303), .A2(new_n597), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n934), .A2(new_n938), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n931), .B(new_n932), .C1(new_n939), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n934), .A2(new_n938), .ZN(new_n944));
  INV_X1    g519(.A(new_n933), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n933), .A2(new_n934), .A3(new_n938), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n946), .A2(new_n930), .A3(new_n947), .A4(KEYINPUT42), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n893), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n639), .A2(new_n640), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n950), .B1(new_n639), .B2(new_n640), .ZN(new_n952));
  AOI211_X1 g527(.A(G299), .B(new_n605), .C1(new_n621), .C2(new_n615), .ZN(new_n953));
  INV_X1    g528(.A(G299), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n615), .A2(new_n621), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n955), .B2(new_n635), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  OR3_X1    g532(.A1(new_n951), .A2(new_n952), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n638), .A2(G299), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT41), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n622), .A2(new_n954), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT41), .B1(new_n953), .B2(new_n956), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n962), .B(new_n963), .C1(new_n951), .C2(new_n952), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n949), .A2(new_n958), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n949), .B1(new_n958), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g541(.A(G868), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n885), .A2(new_n625), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n968), .B1(new_n967), .B2(new_n969), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(G295));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n969), .ZN(G331));
  INV_X1    g548(.A(new_n550), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n885), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n550), .A2(new_n879), .A3(new_n875), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n535), .A2(G301), .A3(new_n536), .ZN(new_n977));
  NAND2_X1  g552(.A1(G168), .A2(G171), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n959), .A2(new_n961), .A3(new_n979), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n535), .A2(G301), .A3(new_n536), .ZN(new_n981));
  AOI21_X1  g556(.A(G301), .B1(new_n535), .B2(new_n536), .ZN(new_n982));
  OAI22_X1  g557(.A1(new_n891), .A2(new_n892), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n963), .A2(new_n985), .A3(new_n962), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  OAI221_X1 g563(.A(KEYINPUT113), .B1(new_n981), .B2(new_n982), .C1(new_n891), .C2(new_n892), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(new_n989), .A3(new_n979), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n962), .B2(new_n985), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n984), .B1(new_n986), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n939), .A2(new_n942), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n927), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n979), .A2(new_n983), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n963), .B2(new_n962), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n988), .A2(new_n989), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n959), .A2(new_n961), .A3(new_n979), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n946), .A2(new_n947), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n995), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n994), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1005));
  INV_X1    g580(.A(new_n996), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n953), .A2(new_n956), .A3(KEYINPUT41), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n960), .B1(new_n959), .B2(new_n961), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n980), .A2(new_n988), .A3(new_n989), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(new_n1002), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n993), .B1(new_n997), .B2(new_n1000), .ZN(new_n1012));
  INV_X1    g587(.A(G37), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1005), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT43), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n994), .A2(new_n1003), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1014), .A2(KEYINPUT43), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1016), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI211_X1 g597(.A(KEYINPUT115), .B(KEYINPUT44), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1015), .B1(new_n1022), .B2(new_n1023), .ZN(G397));
  INV_X1    g599(.A(G1384), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n903), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n472), .A2(G101), .ZN(new_n1028));
  INV_X1    g603(.A(G137), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1028), .B1(new_n723), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G40), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1030), .A2(new_n465), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1026), .A2(new_n1027), .A3(new_n1032), .ZN(new_n1033));
  XOR2_X1   g608(.A(new_n780), .B(G2067), .Z(new_n1034));
  NAND2_X1  g609(.A1(new_n726), .A2(G1996), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1033), .A2(G1996), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1036), .B1(new_n1039), .B2(new_n727), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1033), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n817), .A2(new_n819), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n819), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G290), .A2(G1986), .ZN(new_n1046));
  XOR2_X1   g621(.A(new_n1046), .B(KEYINPUT116), .Z(new_n1047));
  NAND2_X1  g622(.A1(G290), .A2(G1986), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1033), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n568), .B2(new_n572), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1055));
  INV_X1    g630(.A(new_n492), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n900), .B1(new_n1056), .B2(new_n490), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n1025), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1055), .A2(new_n1032), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n797), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1027), .B1(G164), .B2(G1384), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n466), .A2(G40), .A3(new_n473), .ZN(new_n1063));
  AOI21_X1  g638(.A(G1384), .B1(new_n900), .B2(new_n902), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1063), .B1(new_n1064), .B2(KEYINPUT45), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT56), .B(G2072), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1054), .A2(new_n1061), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1032), .A2(new_n1064), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(G2067), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1063), .B1(new_n1064), .B2(new_n1058), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1070), .B1(new_n1073), .B2(new_n802), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(new_n638), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1054), .B1(new_n1061), .B2(new_n1067), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1068), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(KEYINPUT124), .B(new_n1068), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT61), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1068), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(new_n1076), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n638), .B1(new_n1074), .B2(KEYINPUT60), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(KEYINPUT60), .B2(new_n1074), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1061), .A2(new_n1067), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1054), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(KEYINPUT61), .A3(new_n1068), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1083), .A2(new_n1085), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1069), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT58), .B(G1341), .ZN(new_n1093));
  OAI22_X1  g668(.A1(new_n1091), .A2(G1996), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n550), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(KEYINPUT59), .A3(new_n550), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1074), .A2(KEYINPUT60), .A3(new_n638), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1079), .B(new_n1080), .C1(new_n1090), .C2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n903), .A2(new_n1058), .A3(new_n1025), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n1032), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1058), .B1(new_n1057), .B2(new_n1025), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1106), .A2(G1961), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1091), .B2(G2078), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1064), .A2(KEYINPUT45), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n901), .B1(new_n494), .B2(new_n496), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1027), .B1(new_n1111), .B2(G1384), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1108), .A2(G2078), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1110), .A2(new_n1112), .A3(new_n1032), .A4(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1107), .A2(G301), .A3(new_n1109), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT126), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1057), .A2(KEYINPUT45), .A3(new_n1025), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1117), .A2(new_n1032), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1107), .A2(new_n1109), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G171), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1116), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1115), .A2(KEYINPUT126), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1102), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1069), .A2(G8), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT119), .B1(new_n1069), .B2(G8), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n847), .A2(G1976), .A3(new_n848), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n1126), .A2(new_n1127), .B1(new_n1128), .B2(KEYINPUT120), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(KEYINPUT120), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT52), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1124), .B(new_n1125), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n937), .A2(new_n1134), .A3(G1976), .ZN(new_n1135));
  INV_X1    g710(.A(G1976), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT52), .B1(G288), .B2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1133), .A2(new_n1135), .A3(new_n1130), .A4(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n588), .B1(new_n590), .B2(new_n517), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(G1981), .ZN(new_n1140));
  INV_X1    g715(.A(G1981), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n588), .B(new_n1141), .C1(new_n590), .C2(new_n589), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT49), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1140), .A2(KEYINPUT49), .A3(new_n1142), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1133), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1132), .A2(new_n1138), .A3(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT55), .ZN(new_n1150));
  INV_X1    g725(.A(G8), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(G166), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1110), .A2(new_n1032), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT45), .B1(new_n1057), .B2(new_n1025), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n838), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1055), .A2(new_n1059), .A3(new_n754), .A4(new_n1032), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1151), .B1(new_n1158), .B2(KEYINPUT122), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1156), .A2(new_n1160), .A3(new_n1157), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1153), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1071), .A2(new_n1072), .A3(new_n754), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT118), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1071), .A2(new_n1072), .A3(KEYINPUT118), .A4(new_n754), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1165), .A2(new_n1156), .A3(new_n1166), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1167), .A2(new_n1153), .A3(G8), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n1148), .A2(new_n1162), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT51), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n535), .A2(G8), .A3(new_n536), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1171), .B(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(G2084), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1117), .A2(new_n1032), .A3(new_n1112), .ZN(new_n1175));
  INV_X1    g750(.A(G1966), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1106), .A2(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1170), .B(new_n1173), .C1(new_n1177), .C2(new_n1151), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT51), .B1(new_n1177), .B2(new_n1173), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1171), .B(KEYINPUT125), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1071), .A2(new_n1072), .A3(new_n1174), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1180), .B1(new_n1183), .B2(G8), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1178), .B1(new_n1179), .B2(new_n1184), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1119), .A2(G171), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1107), .A2(new_n1109), .A3(new_n1114), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1102), .B1(new_n1187), .B2(G171), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1185), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1101), .A2(new_n1123), .A3(new_n1169), .A4(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1120), .B1(new_n1185), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1169), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n1185), .A2(new_n1191), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1193), .B1(new_n1169), .B2(new_n1192), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1190), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AND3_X1   g773(.A1(new_n1132), .A2(new_n1138), .A3(new_n1147), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT63), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1183), .A2(new_n1200), .A3(G8), .A4(G168), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1158), .A2(KEYINPUT122), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1202), .A2(G8), .A3(new_n1161), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1153), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1201), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1199), .B1(new_n1205), .B2(new_n1168), .ZN(new_n1206));
  NOR3_X1   g781(.A1(new_n1177), .A2(new_n1151), .A3(G286), .ZN(new_n1207));
  AOI22_X1  g782(.A1(new_n1163), .A2(new_n1164), .B1(new_n1091), .B2(new_n838), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1151), .B1(new_n1208), .B2(new_n1166), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1207), .B1(new_n1209), .B2(new_n1153), .ZN(new_n1210));
  OAI21_X1  g785(.A(KEYINPUT63), .B1(new_n1210), .B2(new_n1148), .ZN(new_n1211));
  NOR2_X1   g786(.A1(G288), .A2(G1976), .ZN(new_n1212));
  XOR2_X1   g787(.A(new_n1212), .B(KEYINPUT121), .Z(new_n1213));
  AOI21_X1  g788(.A(new_n1213), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1142), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1133), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1206), .A2(new_n1211), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT123), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND4_X1  g794(.A1(new_n1206), .A2(new_n1211), .A3(KEYINPUT123), .A4(new_n1216), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1050), .B1(new_n1198), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT46), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n1039), .B(new_n1223), .ZN(new_n1224));
  AND2_X1   g799(.A1(new_n1034), .A2(new_n727), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n1224), .B1(new_n1033), .B2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g801(.A(new_n1226), .B(KEYINPUT47), .ZN(new_n1227));
  AND2_X1   g802(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1228));
  NOR2_X1   g803(.A1(new_n780), .A2(G2067), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1041), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1047), .A2(new_n1033), .ZN(new_n1231));
  XNOR2_X1  g806(.A(new_n1231), .B(KEYINPUT48), .ZN(new_n1232));
  OAI211_X1 g807(.A(new_n1227), .B(new_n1230), .C1(new_n1045), .C2(new_n1232), .ZN(new_n1233));
  INV_X1    g808(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1222), .A2(new_n1234), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g810(.A(G319), .ZN(new_n1237));
  NOR4_X1   g811(.A1(G229), .A2(new_n1237), .A3(G401), .A4(G227), .ZN(new_n1238));
  NAND3_X1  g812(.A1(new_n1238), .A2(new_n928), .A3(new_n1020), .ZN(G225));
  INV_X1    g813(.A(G225), .ZN(G308));
endmodule


