

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778;

  XNOR2_X1 U369 ( .A(n597), .B(KEYINPUT42), .ZN(n775) );
  XNOR2_X1 U370 ( .A(G119), .B(G128), .ZN(n560) );
  INV_X2 U371 ( .A(n747), .ZN(n656) );
  INV_X2 U372 ( .A(KEYINPUT76), .ZN(n459) );
  XNOR2_X1 U373 ( .A(n443), .B(n460), .ZN(n645) );
  XNOR2_X2 U374 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X2 U375 ( .A(n660), .B(n659), .ZN(n661) );
  XOR2_X2 U376 ( .A(n654), .B(n653), .Z(n500) );
  NAND2_X1 U377 ( .A1(n349), .A2(n447), .ZN(n478) );
  INV_X1 U378 ( .A(n645), .ZN(n349) );
  XNOR2_X1 U379 ( .A(n481), .B(n523), .ZN(n563) );
  NOR2_X1 U380 ( .A1(n725), .A2(n605), .ZN(n597) );
  XNOR2_X1 U381 ( .A(n475), .B(n474), .ZN(n778) );
  XNOR2_X2 U382 ( .A(n472), .B(n469), .ZN(n408) );
  AND2_X2 U383 ( .A1(n456), .A2(n457), .ZN(n455) );
  XNOR2_X2 U384 ( .A(KEYINPUT38), .B(n585), .ZN(n709) );
  AND2_X2 U385 ( .A1(n399), .A2(n398), .ZN(n397) );
  AND2_X2 U386 ( .A1(n646), .A2(n494), .ZN(n479) );
  NAND2_X2 U387 ( .A1(n634), .A2(KEYINPUT44), .ZN(n646) );
  XNOR2_X2 U388 ( .A(n551), .B(n552), .ZN(n737) );
  INV_X1 U389 ( .A(n778), .ZN(n352) );
  XNOR2_X2 U390 ( .A(n578), .B(n752), .ZN(n472) );
  INV_X1 U391 ( .A(G146), .ZN(n361) );
  INV_X1 U392 ( .A(G125), .ZN(n362) );
  AND2_X1 U393 ( .A1(n422), .A2(n421), .ZN(n420) );
  XNOR2_X1 U394 ( .A(n351), .B(KEYINPUT103), .ZN(n496) );
  NAND2_X1 U395 ( .A1(n426), .A2(n425), .ZN(n424) );
  NAND2_X1 U396 ( .A1(n353), .A2(n352), .ZN(n351) );
  AND2_X1 U397 ( .A1(n429), .A2(n428), .ZN(n427) );
  AND2_X1 U398 ( .A1(n388), .A2(n386), .ZN(n385) );
  OR2_X1 U399 ( .A1(n674), .A2(n690), .ZN(n643) );
  XNOR2_X1 U400 ( .A(n394), .B(n393), .ZN(n725) );
  NOR2_X1 U401 ( .A1(n671), .A2(n430), .ZN(n425) );
  NAND2_X1 U402 ( .A1(n604), .A2(n708), .ZN(n497) );
  BUF_X1 U403 ( .A(n698), .Z(n444) );
  XNOR2_X1 U404 ( .A(n470), .B(n579), .ZN(n469) );
  XNOR2_X1 U405 ( .A(n440), .B(n574), .ZN(n470) );
  XNOR2_X1 U406 ( .A(n575), .B(n471), .ZN(n440) );
  XNOR2_X1 U407 ( .A(n452), .B(n450), .ZN(n753) );
  NAND2_X1 U408 ( .A1(n363), .A2(n364), .ZN(n573) );
  XNOR2_X1 U409 ( .A(n414), .B(KEYINPUT75), .ZN(n452) );
  INV_X1 U410 ( .A(KEYINPUT64), .ZN(n480) );
  NAND2_X1 U411 ( .A1(n643), .A2(n637), .ZN(n353) );
  NAND2_X1 U412 ( .A1(n427), .A2(n424), .ZN(n354) );
  NAND2_X1 U413 ( .A1(n427), .A2(n424), .ZN(n777) );
  OR2_X2 U414 ( .A1(n644), .A2(n366), .ZN(n634) );
  XNOR2_X1 U415 ( .A(KEYINPUT30), .B(n356), .ZN(n355) );
  NOR2_X1 U416 ( .A1(n539), .A2(n416), .ZN(n356) );
  AND2_X2 U417 ( .A1(n492), .A2(n491), .ZN(n357) );
  BUF_X1 U418 ( .A(n737), .Z(n358) );
  XNOR2_X1 U419 ( .A(n554), .B(n369), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n554), .B(n369), .ZN(n488) );
  BUF_X1 U421 ( .A(n729), .Z(n360) );
  NAND2_X1 U422 ( .A1(G146), .A2(n362), .ZN(n363) );
  NAND2_X1 U423 ( .A1(n361), .A2(G125), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n558), .B(n559), .ZN(n365) );
  XOR2_X2 U425 ( .A(G137), .B(G140), .Z(n559) );
  BUF_X1 U426 ( .A(n772), .Z(n366) );
  XNOR2_X1 U427 ( .A(n449), .B(n448), .ZN(n367) );
  BUF_X1 U428 ( .A(n726), .Z(n368) );
  XNOR2_X1 U429 ( .A(n628), .B(KEYINPUT35), .ZN(n772) );
  NAND2_X2 U430 ( .A1(n730), .A2(n652), .ZN(n449) );
  NAND2_X1 U431 ( .A1(n419), .A2(n418), .ZN(n417) );
  AND2_X1 U432 ( .A1(n423), .A2(KEYINPUT46), .ZN(n418) );
  NAND2_X1 U433 ( .A1(n775), .A2(n431), .ZN(n421) );
  INV_X1 U434 ( .A(KEYINPUT74), .ZN(n460) );
  NAND2_X1 U435 ( .A1(n420), .A2(n417), .ZN(n485) );
  XOR2_X1 U436 ( .A(KEYINPUT7), .B(KEYINPUT95), .Z(n519) );
  AND2_X1 U437 ( .A1(n631), .A2(n390), .ZN(n389) );
  INV_X1 U438 ( .A(KEYINPUT1), .ZN(n415) );
  INV_X1 U439 ( .A(KEYINPUT66), .ZN(n448) );
  INV_X1 U440 ( .A(KEYINPUT41), .ZN(n393) );
  NOR2_X1 U441 ( .A1(n712), .A2(n416), .ZN(n395) );
  INV_X1 U442 ( .A(n389), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n632), .B(KEYINPUT79), .ZN(n490) );
  XNOR2_X1 U444 ( .A(n411), .B(KEYINPUT77), .ZN(n586) );
  XNOR2_X1 U445 ( .A(n468), .B(n467), .ZN(n466) );
  XNOR2_X1 U446 ( .A(KEYINPUT107), .B(KEYINPUT28), .ZN(n467) );
  INV_X1 U447 ( .A(n445), .ZN(n636) );
  BUF_X1 U448 ( .A(n763), .Z(n412) );
  XNOR2_X1 U449 ( .A(n521), .B(n442), .ZN(n525) );
  XNOR2_X1 U450 ( .A(n522), .B(n373), .ZN(n442) );
  XOR2_X1 U451 ( .A(KEYINPUT5), .B(G137), .Z(n532) );
  NOR2_X1 U452 ( .A1(G953), .A2(G237), .ZN(n530) );
  NAND2_X1 U453 ( .A1(G234), .A2(G237), .ZN(n540) );
  XNOR2_X1 U454 ( .A(G902), .B(KEYINPUT15), .ZN(n649) );
  OR2_X1 U455 ( .A1(G237), .A2(G902), .ZN(n580) );
  XNOR2_X1 U456 ( .A(G131), .B(G134), .ZN(n529) );
  XNOR2_X1 U457 ( .A(n534), .B(n533), .ZN(n576) );
  XNOR2_X1 U458 ( .A(KEYINPUT3), .B(G119), .ZN(n533) );
  XOR2_X1 U459 ( .A(G113), .B(G116), .Z(n534) );
  NAND2_X1 U460 ( .A1(n495), .A2(n647), .ZN(n491) );
  XOR2_X1 U461 ( .A(G140), .B(KEYINPUT94), .Z(n502) );
  XNOR2_X1 U462 ( .A(G113), .B(G143), .ZN(n507) );
  XOR2_X1 U463 ( .A(G122), .B(G104), .Z(n508) );
  XNOR2_X1 U464 ( .A(G131), .B(KEYINPUT93), .ZN(n503) );
  XOR2_X1 U465 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n504) );
  INV_X1 U466 ( .A(KEYINPUT17), .ZN(n471) );
  NOR2_X1 U467 ( .A1(n770), .A2(n464), .ZN(n463) );
  INV_X1 U468 ( .A(n771), .ZN(n464) );
  XNOR2_X1 U469 ( .A(n576), .B(n441), .ZN(n752) );
  XNOR2_X1 U470 ( .A(KEYINPUT16), .B(G122), .ZN(n441) );
  XNOR2_X1 U471 ( .A(n451), .B(G110), .ZN(n450) );
  INV_X1 U472 ( .A(G104), .ZN(n451) );
  XNOR2_X1 U473 ( .A(KEYINPUT8), .B(KEYINPUT71), .ZN(n523) );
  XNOR2_X1 U474 ( .A(G116), .B(G134), .ZN(n516) );
  XNOR2_X1 U475 ( .A(G122), .B(KEYINPUT97), .ZN(n518) );
  INV_X1 U476 ( .A(KEYINPUT40), .ZN(n430) );
  NAND2_X1 U477 ( .A1(n671), .A2(n430), .ZN(n428) );
  AND2_X1 U478 ( .A1(n404), .A2(n402), .ZN(n401) );
  XOR2_X1 U479 ( .A(n527), .B(n526), .Z(n593) );
  XNOR2_X1 U480 ( .A(n486), .B(KEYINPUT91), .ZN(n638) );
  NAND2_X1 U481 ( .A1(n590), .A2(n593), .ZN(n671) );
  NAND2_X1 U482 ( .A1(n385), .A2(n382), .ZN(n774) );
  NAND2_X1 U483 ( .A1(n384), .A2(n376), .ZN(n382) );
  NAND2_X1 U484 ( .A1(n387), .A2(n490), .ZN(n386) );
  NOR2_X1 U485 ( .A1(n370), .A2(n605), .ZN(n606) );
  NAND2_X1 U486 ( .A1(n384), .A2(n391), .ZN(n679) );
  NOR2_X1 U487 ( .A1(n596), .A2(n444), .ZN(n392) );
  BUF_X1 U488 ( .A(G107), .Z(n446) );
  INV_X1 U489 ( .A(KEYINPUT102), .ZN(n474) );
  XNOR2_X1 U490 ( .A(n743), .B(n744), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n741), .B(n742), .ZN(n432) );
  INV_X1 U492 ( .A(KEYINPUT56), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n736), .B(n433), .ZN(G75) );
  XNOR2_X1 U494 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n433) );
  XOR2_X1 U495 ( .A(KEYINPUT73), .B(n553), .Z(n369) );
  XOR2_X1 U496 ( .A(n407), .B(KEYINPUT19), .Z(n370) );
  AND2_X1 U497 ( .A1(n697), .A2(n629), .ZN(n371) );
  AND2_X1 U498 ( .A1(G210), .A2(n580), .ZN(n372) );
  XNOR2_X1 U499 ( .A(KEYINPUT96), .B(KEYINPUT9), .ZN(n373) );
  AND2_X1 U500 ( .A1(n396), .A2(n627), .ZN(n374) );
  AND2_X1 U501 ( .A1(n638), .A2(n594), .ZN(n375) );
  NAND2_X1 U502 ( .A1(n492), .A2(n491), .ZN(n410) );
  AND2_X1 U503 ( .A1(n389), .A2(n383), .ZN(n376) );
  AND2_X1 U504 ( .A1(n357), .A2(n735), .ZN(n377) );
  INV_X1 U505 ( .A(n708), .ZN(n416) );
  INV_X1 U506 ( .A(KEYINPUT34), .ZN(n402) );
  XOR2_X1 U507 ( .A(n624), .B(KEYINPUT0), .Z(n378) );
  XOR2_X1 U508 ( .A(KEYINPUT6), .B(KEYINPUT101), .Z(n379) );
  XNOR2_X1 U509 ( .A(n611), .B(KEYINPUT48), .ZN(n380) );
  XOR2_X1 U510 ( .A(n664), .B(KEYINPUT86), .Z(n381) );
  INV_X1 U511 ( .A(n490), .ZN(n383) );
  INV_X1 U512 ( .A(n633), .ZN(n384) );
  NAND2_X1 U513 ( .A1(n633), .A2(n490), .ZN(n388) );
  NOR2_X1 U514 ( .A1(n633), .A2(n630), .ZN(n635) );
  INV_X1 U515 ( .A(n630), .ZN(n390) );
  NAND2_X1 U516 ( .A1(n774), .A2(n679), .ZN(n644) );
  AND2_X1 U517 ( .A1(n445), .A2(n392), .ZN(n391) );
  NAND2_X1 U518 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U519 ( .A1(n709), .A2(n395), .ZN(n394) );
  NAND2_X1 U520 ( .A1(n397), .A2(n374), .ZN(n628) );
  NAND2_X1 U521 ( .A1(n473), .A2(KEYINPUT34), .ZN(n396) );
  NAND2_X1 U522 ( .A1(n726), .A2(KEYINPUT34), .ZN(n398) );
  NAND2_X1 U523 ( .A1(n400), .A2(n401), .ZN(n399) );
  INV_X1 U524 ( .A(n726), .ZN(n400) );
  INV_X1 U525 ( .A(n404), .ZN(n473) );
  XNOR2_X2 U526 ( .A(n625), .B(n626), .ZN(n726) );
  NAND2_X1 U527 ( .A1(n404), .A2(n371), .ZN(n498) );
  XNOR2_X2 U528 ( .A(n623), .B(n378), .ZN(n404) );
  OR2_X1 U529 ( .A1(n473), .A2(n403), .ZN(n639) );
  INV_X1 U530 ( .A(n638), .ZN(n403) );
  NAND2_X1 U531 ( .A1(n704), .A2(n404), .ZN(n642) );
  AND2_X2 U532 ( .A1(n729), .A2(n650), .ZN(n652) );
  XNOR2_X1 U533 ( .A(n558), .B(n559), .ZN(n759) );
  BUF_X1 U534 ( .A(n695), .Z(n445) );
  XNOR2_X1 U535 ( .A(n745), .B(n746), .ZN(n413) );
  NAND2_X1 U536 ( .A1(n465), .A2(n463), .ZN(n762) );
  INV_X1 U537 ( .A(n354), .ZN(n419) );
  NOR2_X2 U538 ( .A1(n746), .A2(G902), .ZN(n571) );
  XNOR2_X1 U539 ( .A(n488), .B(n415), .ZN(n695) );
  NOR2_X2 U540 ( .A1(n737), .A2(G902), .ZN(n554) );
  XNOR2_X2 U541 ( .A(n405), .B(G472), .ZN(n539) );
  NOR2_X1 U542 ( .A1(n658), .A2(G902), .ZN(n405) );
  BUF_X1 U543 ( .A(n753), .Z(n406) );
  BUF_X1 U544 ( .A(n604), .Z(n615) );
  NOR2_X1 U545 ( .A1(n762), .A2(n459), .ZN(n454) );
  NOR2_X1 U546 ( .A1(n762), .A2(n459), .ZN(n458) );
  BUF_X1 U547 ( .A(n497), .Z(n407) );
  INV_X1 U548 ( .A(n539), .ZN(n596) );
  NAND2_X1 U549 ( .A1(n596), .A2(n598), .ZN(n468) );
  XNOR2_X1 U550 ( .A(n497), .B(KEYINPUT19), .ZN(n622) );
  BUF_X1 U551 ( .A(n730), .Z(n409) );
  NAND2_X1 U552 ( .A1(n410), .A2(n459), .ZN(n456) );
  NAND2_X1 U553 ( .A1(n439), .A2(n648), .ZN(n729) );
  NAND2_X1 U554 ( .A1(n408), .A2(n649), .ZN(n581) );
  NAND2_X1 U555 ( .A1(n375), .A2(n355), .ZN(n411) );
  NOR2_X1 U556 ( .A1(n413), .A2(n747), .ZN(G66) );
  XNOR2_X2 U557 ( .A(G107), .B(KEYINPUT87), .ZN(n414) );
  XNOR2_X2 U558 ( .A(n539), .B(n379), .ZN(n630) );
  INV_X1 U559 ( .A(n775), .ZN(n423) );
  NAND2_X1 U560 ( .A1(n777), .A2(n431), .ZN(n422) );
  INV_X1 U561 ( .A(n591), .ZN(n426) );
  NAND2_X1 U562 ( .A1(n591), .A2(n430), .ZN(n429) );
  INV_X1 U563 ( .A(KEYINPUT46), .ZN(n431) );
  NAND2_X1 U564 ( .A1(n740), .A2(G475), .ZN(n668) );
  XNOR2_X2 U565 ( .A(n449), .B(n448), .ZN(n740) );
  NOR2_X1 U566 ( .A1(n432), .A2(n747), .ZN(G54) );
  NOR2_X1 U567 ( .A1(n434), .A2(n747), .ZN(G63) );
  XNOR2_X1 U568 ( .A(n435), .B(n670), .ZN(G60) );
  NAND2_X1 U569 ( .A1(n669), .A2(n656), .ZN(n435) );
  XNOR2_X1 U570 ( .A(n437), .B(n436), .ZN(G51) );
  NAND2_X1 U571 ( .A1(n657), .A2(n656), .ZN(n437) );
  XNOR2_X1 U572 ( .A(n438), .B(n381), .ZN(G57) );
  NAND2_X1 U573 ( .A1(n663), .A2(n656), .ZN(n438) );
  XNOR2_X2 U574 ( .A(n753), .B(n547), .ZN(n578) );
  XNOR2_X1 U575 ( .A(n482), .B(n380), .ZN(n465) );
  NAND2_X1 U576 ( .A1(n357), .A2(n458), .ZN(n439) );
  NAND2_X1 U577 ( .A1(n762), .A2(n459), .ZN(n457) );
  NAND2_X1 U578 ( .A1(n461), .A2(n489), .ZN(n443) );
  XNOR2_X1 U579 ( .A(n551), .B(n538), .ZN(n658) );
  XNOR2_X2 U580 ( .A(n573), .B(KEYINPUT10), .ZN(n558) );
  XNOR2_X2 U581 ( .A(n583), .B(n582), .ZN(n591) );
  NAND2_X1 U582 ( .A1(n740), .A2(G210), .ZN(n655) );
  NAND2_X1 U583 ( .A1(n479), .A2(n496), .ZN(n447) );
  XNOR2_X2 U584 ( .A(n761), .B(G146), .ZN(n551) );
  NAND2_X1 U585 ( .A1(n455), .A2(n453), .ZN(n651) );
  NAND2_X1 U586 ( .A1(n357), .A2(n454), .ZN(n453) );
  XNOR2_X1 U587 ( .A(n462), .B(KEYINPUT70), .ZN(n461) );
  NOR2_X2 U588 ( .A1(n772), .A2(KEYINPUT44), .ZN(n462) );
  NAND2_X1 U589 ( .A1(n466), .A2(n359), .ZN(n605) );
  NAND2_X1 U590 ( .A1(n635), .A2(n476), .ZN(n475) );
  NOR2_X1 U591 ( .A1(n636), .A2(n477), .ZN(n476) );
  INV_X1 U592 ( .A(n444), .ZN(n477) );
  NAND2_X1 U593 ( .A1(n478), .A2(n493), .ZN(n492) );
  NAND2_X1 U594 ( .A1(n359), .A2(n487), .ZN(n486) );
  NOR2_X2 U595 ( .A1(n695), .A2(n694), .ZN(n640) );
  AND2_X1 U596 ( .A1(n610), .A2(n484), .ZN(n483) );
  XNOR2_X2 U597 ( .A(n480), .B(G953), .ZN(n763) );
  NAND2_X1 U598 ( .A1(n563), .A2(G221), .ZN(n564) );
  NAND2_X1 U599 ( .A1(n763), .A2(G234), .ZN(n481) );
  NAND2_X1 U600 ( .A1(n485), .A2(n483), .ZN(n482) );
  INV_X1 U601 ( .A(n683), .ZN(n484) );
  INV_X1 U602 ( .A(n694), .ZN(n487) );
  NAND2_X2 U603 ( .A1(n698), .A2(n697), .ZN(n694) );
  XNOR2_X2 U604 ( .A(n571), .B(n570), .ZN(n698) );
  INV_X1 U605 ( .A(n644), .ZN(n489) );
  NAND2_X1 U606 ( .A1(n645), .A2(n494), .ZN(n493) );
  INV_X1 U607 ( .A(n647), .ZN(n494) );
  NAND2_X1 U608 ( .A1(n646), .A2(n496), .ZN(n495) );
  INV_X1 U609 ( .A(n615), .ZN(n585) );
  XNOR2_X2 U610 ( .A(n581), .B(n372), .ZN(n604) );
  XNOR2_X2 U611 ( .A(n498), .B(KEYINPUT22), .ZN(n633) );
  XNOR2_X1 U612 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U613 ( .A(n550), .B(n578), .ZN(n552) );
  XNOR2_X1 U614 ( .A(n562), .B(KEYINPUT83), .ZN(n499) );
  INV_X1 U615 ( .A(KEYINPUT18), .ZN(n572) );
  XNOR2_X1 U616 ( .A(n573), .B(n572), .ZN(n574) );
  BUF_X1 U617 ( .A(n577), .Z(n579) );
  XNOR2_X1 U618 ( .A(n576), .B(n535), .ZN(n537) );
  XNOR2_X1 U619 ( .A(n537), .B(n547), .ZN(n538) );
  INV_X1 U620 ( .A(KEYINPUT67), .ZN(n624) );
  INV_X1 U621 ( .A(KEYINPUT39), .ZN(n582) );
  INV_X1 U622 ( .A(KEYINPUT63), .ZN(n664) );
  XNOR2_X1 U623 ( .A(n565), .B(n566), .ZN(n746) );
  NOR2_X1 U624 ( .A1(G952), .A2(n412), .ZN(n747) );
  XNOR2_X1 U625 ( .A(KEYINPUT13), .B(G475), .ZN(n514) );
  NAND2_X1 U626 ( .A1(G214), .A2(n530), .ZN(n501) );
  XNOR2_X1 U627 ( .A(n502), .B(n501), .ZN(n506) );
  XNOR2_X1 U628 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U629 ( .A(n506), .B(n505), .Z(n512) );
  INV_X1 U630 ( .A(n558), .ZN(n510) );
  XNOR2_X1 U631 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U632 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U633 ( .A(n512), .B(n511), .ZN(n666) );
  NOR2_X1 U634 ( .A1(G902), .A2(n666), .ZN(n513) );
  XNOR2_X1 U635 ( .A(n514), .B(n513), .ZN(n590) );
  XNOR2_X1 U636 ( .A(G478), .B(KEYINPUT99), .ZN(n515) );
  XNOR2_X1 U637 ( .A(n515), .B(KEYINPUT98), .ZN(n527) );
  XNOR2_X1 U638 ( .A(n516), .B(n446), .ZN(n522) );
  XNOR2_X2 U639 ( .A(G128), .B(KEYINPUT81), .ZN(n517) );
  XNOR2_X2 U640 ( .A(n517), .B(G143), .ZN(n528) );
  XNOR2_X1 U641 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U642 ( .A(n528), .B(n520), .ZN(n521) );
  NAND2_X1 U643 ( .A1(G217), .A2(n563), .ZN(n524) );
  XNOR2_X1 U644 ( .A(n525), .B(n524), .ZN(n744) );
  NOR2_X1 U645 ( .A1(G902), .A2(n744), .ZN(n526) );
  NOR2_X1 U646 ( .A1(n590), .A2(n593), .ZN(n689) );
  XOR2_X1 U647 ( .A(KEYINPUT100), .B(n689), .Z(n607) );
  XNOR2_X2 U648 ( .A(n528), .B(KEYINPUT4), .ZN(n577) );
  XNOR2_X2 U649 ( .A(n577), .B(n529), .ZN(n761) );
  NAND2_X1 U650 ( .A1(n530), .A2(G210), .ZN(n531) );
  XNOR2_X1 U651 ( .A(n532), .B(n531), .ZN(n535) );
  XNOR2_X1 U652 ( .A(G101), .B(KEYINPUT69), .ZN(n536) );
  XNOR2_X1 U653 ( .A(n536), .B(KEYINPUT68), .ZN(n547) );
  NAND2_X1 U654 ( .A1(G214), .A2(n580), .ZN(n708) );
  INV_X1 U655 ( .A(n412), .ZN(n542) );
  XNOR2_X1 U656 ( .A(n540), .B(KEYINPUT14), .ZN(n543) );
  NAND2_X1 U657 ( .A1(G902), .A2(n543), .ZN(n617) );
  NOR2_X1 U658 ( .A1(G900), .A2(n617), .ZN(n541) );
  NAND2_X1 U659 ( .A1(n542), .A2(n541), .ZN(n545) );
  NAND2_X1 U660 ( .A1(G952), .A2(n543), .ZN(n724) );
  NOR2_X1 U661 ( .A1(G953), .A2(n724), .ZN(n544) );
  XOR2_X1 U662 ( .A(KEYINPUT88), .B(n544), .Z(n619) );
  NAND2_X1 U663 ( .A1(n545), .A2(n619), .ZN(n546) );
  XNOR2_X1 U664 ( .A(n546), .B(KEYINPUT82), .ZN(n594) );
  XOR2_X1 U665 ( .A(n559), .B(KEYINPUT78), .Z(n549) );
  NAND2_X1 U666 ( .A1(G227), .A2(n763), .ZN(n548) );
  XNOR2_X1 U667 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U668 ( .A(G469), .B(KEYINPUT72), .Z(n553) );
  XOR2_X1 U669 ( .A(KEYINPUT90), .B(KEYINPUT21), .Z(n557) );
  NAND2_X1 U670 ( .A1(G234), .A2(n649), .ZN(n555) );
  XNOR2_X1 U671 ( .A(KEYINPUT20), .B(n555), .ZN(n567) );
  NAND2_X1 U672 ( .A1(G221), .A2(n567), .ZN(n556) );
  XNOR2_X1 U673 ( .A(n557), .B(n556), .ZN(n697) );
  XNOR2_X1 U674 ( .A(n759), .B(KEYINPUT23), .ZN(n566) );
  XOR2_X1 U675 ( .A(KEYINPUT24), .B(G110), .Z(n561) );
  XNOR2_X1 U676 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U677 ( .A(n499), .B(n564), .ZN(n565) );
  XOR2_X1 U678 ( .A(KEYINPUT89), .B(KEYINPUT25), .Z(n569) );
  NAND2_X1 U679 ( .A1(n567), .A2(G217), .ZN(n568) );
  XNOR2_X1 U680 ( .A(n569), .B(n568), .ZN(n570) );
  NAND2_X1 U681 ( .A1(G224), .A2(n763), .ZN(n575) );
  NAND2_X1 U682 ( .A1(n586), .A2(n709), .ZN(n583) );
  OR2_X1 U683 ( .A1(n607), .A2(n591), .ZN(n584) );
  XNOR2_X1 U684 ( .A(n584), .B(KEYINPUT109), .ZN(n770) );
  INV_X1 U685 ( .A(n590), .ZN(n592) );
  NOR2_X1 U686 ( .A1(n592), .A2(n593), .ZN(n627) );
  INV_X1 U687 ( .A(n627), .ZN(n589) );
  AND2_X1 U688 ( .A1(n586), .A2(n615), .ZN(n587) );
  XOR2_X1 U689 ( .A(KEYINPUT106), .B(n587), .Z(n588) );
  NOR2_X1 U690 ( .A1(n589), .A2(n588), .ZN(n683) );
  NAND2_X1 U691 ( .A1(n593), .A2(n592), .ZN(n712) );
  NAND2_X1 U692 ( .A1(n697), .A2(n594), .ZN(n595) );
  NOR2_X1 U693 ( .A1(n444), .A2(n595), .ZN(n598) );
  XOR2_X1 U694 ( .A(KEYINPUT36), .B(KEYINPUT108), .Z(n602) );
  NAND2_X1 U695 ( .A1(n630), .A2(n598), .ZN(n599) );
  NOR2_X1 U696 ( .A1(n671), .A2(n599), .ZN(n600) );
  NAND2_X1 U697 ( .A1(n600), .A2(n708), .ZN(n612) );
  NOR2_X1 U698 ( .A1(n612), .A2(n585), .ZN(n601) );
  XNOR2_X1 U699 ( .A(n602), .B(n601), .ZN(n603) );
  NOR2_X1 U700 ( .A1(n445), .A2(n603), .ZN(n692) );
  XNOR2_X1 U701 ( .A(n606), .B(KEYINPUT80), .ZN(n685) );
  NAND2_X1 U702 ( .A1(n607), .A2(n671), .ZN(n637) );
  NAND2_X1 U703 ( .A1(n685), .A2(n637), .ZN(n608) );
  XNOR2_X1 U704 ( .A(KEYINPUT47), .B(n608), .ZN(n609) );
  NOR2_X1 U705 ( .A1(n692), .A2(n609), .ZN(n610) );
  INV_X1 U706 ( .A(KEYINPUT84), .ZN(n611) );
  NOR2_X1 U707 ( .A1(n636), .A2(n612), .ZN(n613) );
  XNOR2_X1 U708 ( .A(n613), .B(KEYINPUT43), .ZN(n614) );
  NOR2_X1 U709 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U710 ( .A(KEYINPUT105), .B(n616), .ZN(n771) );
  INV_X1 U711 ( .A(n617), .ZN(n618) );
  INV_X1 U712 ( .A(G953), .ZN(n735) );
  NOR2_X1 U713 ( .A1(G898), .A2(n735), .ZN(n756) );
  NAND2_X1 U714 ( .A1(n618), .A2(n756), .ZN(n620) );
  NAND2_X1 U715 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U716 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U717 ( .A(KEYINPUT104), .B(KEYINPUT33), .Z(n626) );
  NAND2_X1 U718 ( .A1(n640), .A2(n630), .ZN(n625) );
  INV_X1 U719 ( .A(n712), .ZN(n629) );
  NOR2_X1 U720 ( .A1(n445), .A2(n444), .ZN(n631) );
  INV_X1 U721 ( .A(KEYINPUT32), .ZN(n632) );
  INV_X1 U722 ( .A(n637), .ZN(n714) );
  NOR2_X1 U723 ( .A1(n596), .A2(n639), .ZN(n674) );
  NAND2_X1 U724 ( .A1(n640), .A2(n596), .ZN(n641) );
  XOR2_X1 U725 ( .A(KEYINPUT92), .B(n641), .Z(n704) );
  XNOR2_X1 U726 ( .A(KEYINPUT31), .B(n642), .ZN(n690) );
  XNOR2_X1 U727 ( .A(KEYINPUT45), .B(KEYINPUT65), .ZN(n647) );
  INV_X1 U728 ( .A(KEYINPUT2), .ZN(n648) );
  INV_X1 U729 ( .A(n649), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(KEYINPUT2), .ZN(n730) );
  XOR2_X1 U731 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n654) );
  XNOR2_X1 U732 ( .A(n408), .B(KEYINPUT85), .ZN(n653) );
  XNOR2_X1 U733 ( .A(n655), .B(n500), .ZN(n657) );
  NAND2_X1 U734 ( .A1(n740), .A2(G472), .ZN(n662) );
  XOR2_X1 U735 ( .A(KEYINPUT111), .B(KEYINPUT62), .Z(n660) );
  XOR2_X1 U736 ( .A(n658), .B(KEYINPUT110), .Z(n659) );
  XNOR2_X1 U737 ( .A(n662), .B(n661), .ZN(n663) );
  INV_X1 U738 ( .A(KEYINPUT60), .ZN(n670) );
  XOR2_X1 U739 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n665) );
  INV_X1 U740 ( .A(n671), .ZN(n687) );
  NAND2_X1 U741 ( .A1(n674), .A2(n687), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n672), .B(KEYINPUT112), .ZN(n673) );
  XNOR2_X1 U743 ( .A(G104), .B(n673), .ZN(G6) );
  XOR2_X1 U744 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n676) );
  NAND2_X1 U745 ( .A1(n674), .A2(n689), .ZN(n675) );
  XNOR2_X1 U746 ( .A(n676), .B(n675), .ZN(n678) );
  XOR2_X1 U747 ( .A(n446), .B(KEYINPUT113), .Z(n677) );
  XNOR2_X1 U748 ( .A(n678), .B(n677), .ZN(G9) );
  XNOR2_X1 U749 ( .A(G110), .B(KEYINPUT114), .ZN(n680) );
  XNOR2_X1 U750 ( .A(n680), .B(n679), .ZN(G12) );
  XOR2_X1 U751 ( .A(G128), .B(KEYINPUT29), .Z(n682) );
  NAND2_X1 U752 ( .A1(n689), .A2(n685), .ZN(n681) );
  XNOR2_X1 U753 ( .A(n682), .B(n681), .ZN(G30) );
  XNOR2_X1 U754 ( .A(G143), .B(n683), .ZN(n684) );
  XNOR2_X1 U755 ( .A(n684), .B(KEYINPUT115), .ZN(G45) );
  NAND2_X1 U756 ( .A1(n685), .A2(n687), .ZN(n686) );
  XNOR2_X1 U757 ( .A(n686), .B(G146), .ZN(G48) );
  NAND2_X1 U758 ( .A1(n687), .A2(n690), .ZN(n688) );
  XNOR2_X1 U759 ( .A(G113), .B(n688), .ZN(G15) );
  NAND2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U761 ( .A(n691), .B(G116), .ZN(G18) );
  XNOR2_X1 U762 ( .A(G125), .B(n692), .ZN(n693) );
  XNOR2_X1 U763 ( .A(n693), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U764 ( .A1(n445), .A2(n694), .ZN(n696) );
  XNOR2_X1 U765 ( .A(n696), .B(KEYINPUT50), .ZN(n701) );
  NOR2_X1 U766 ( .A1(n444), .A2(n697), .ZN(n699) );
  XNOR2_X1 U767 ( .A(n699), .B(KEYINPUT49), .ZN(n700) );
  NAND2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U769 ( .A1(n596), .A2(n702), .ZN(n703) );
  NOR2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U771 ( .A(n705), .B(KEYINPUT51), .Z(n706) );
  XNOR2_X1 U772 ( .A(KEYINPUT116), .B(n706), .ZN(n707) );
  NOR2_X1 U773 ( .A1(n725), .A2(n707), .ZN(n720) );
  NOR2_X1 U774 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U775 ( .A(KEYINPUT117), .B(n710), .Z(n711) );
  NOR2_X1 U776 ( .A1(n712), .A2(n711), .ZN(n717) );
  NOR2_X1 U777 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U778 ( .A(n715), .B(KEYINPUT118), .ZN(n716) );
  NOR2_X1 U779 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U780 ( .A1(n368), .A2(n718), .ZN(n719) );
  NOR2_X1 U781 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U782 ( .A(n721), .B(KEYINPUT119), .Z(n722) );
  XNOR2_X1 U783 ( .A(KEYINPUT52), .B(n722), .ZN(n723) );
  NOR2_X1 U784 ( .A1(n724), .A2(n723), .ZN(n728) );
  NOR2_X1 U785 ( .A1(n368), .A2(n725), .ZN(n727) );
  NOR2_X1 U786 ( .A1(n728), .A2(n727), .ZN(n732) );
  NAND2_X1 U787 ( .A1(n409), .A2(n360), .ZN(n731) );
  NAND2_X1 U788 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U789 ( .A(KEYINPUT120), .B(n733), .Z(n734) );
  NAND2_X1 U790 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U791 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n739) );
  XNOR2_X1 U792 ( .A(n358), .B(KEYINPUT122), .ZN(n738) );
  XNOR2_X1 U793 ( .A(n739), .B(n738), .ZN(n742) );
  NAND2_X1 U794 ( .A1(G469), .A2(n367), .ZN(n741) );
  NAND2_X1 U795 ( .A1(G478), .A2(n367), .ZN(n743) );
  NAND2_X1 U796 ( .A1(G217), .A2(n367), .ZN(n745) );
  NAND2_X1 U797 ( .A1(G953), .A2(G224), .ZN(n748) );
  XNOR2_X1 U798 ( .A(KEYINPUT61), .B(n748), .ZN(n749) );
  NAND2_X1 U799 ( .A1(n749), .A2(G898), .ZN(n750) );
  XOR2_X1 U800 ( .A(KEYINPUT124), .B(n750), .Z(n751) );
  NOR2_X1 U801 ( .A1(n751), .A2(n377), .ZN(n758) );
  XNOR2_X1 U802 ( .A(n752), .B(G101), .ZN(n754) );
  XNOR2_X1 U803 ( .A(n406), .B(n754), .ZN(n755) );
  NOR2_X1 U804 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U805 ( .A(n758), .B(n757), .Z(G69) );
  XOR2_X1 U806 ( .A(n365), .B(KEYINPUT125), .Z(n760) );
  XNOR2_X1 U807 ( .A(n761), .B(n760), .ZN(n765) );
  XNOR2_X1 U808 ( .A(n762), .B(n765), .ZN(n764) );
  NAND2_X1 U809 ( .A1(n764), .A2(n412), .ZN(n769) );
  XNOR2_X1 U810 ( .A(G227), .B(n765), .ZN(n766) );
  NAND2_X1 U811 ( .A1(n766), .A2(G900), .ZN(n767) );
  NAND2_X1 U812 ( .A1(n767), .A2(G953), .ZN(n768) );
  NAND2_X1 U813 ( .A1(n769), .A2(n768), .ZN(G72) );
  XOR2_X1 U814 ( .A(G134), .B(n770), .Z(G36) );
  XNOR2_X1 U815 ( .A(G140), .B(n771), .ZN(G42) );
  XNOR2_X1 U816 ( .A(G122), .B(KEYINPUT126), .ZN(n773) );
  XOR2_X1 U817 ( .A(n773), .B(n366), .Z(G24) );
  XNOR2_X1 U818 ( .A(n774), .B(G119), .ZN(G21) );
  XNOR2_X1 U819 ( .A(G137), .B(KEYINPUT127), .ZN(n776) );
  XNOR2_X1 U820 ( .A(n776), .B(n775), .ZN(G39) );
  XOR2_X1 U821 ( .A(n354), .B(G131), .Z(G33) );
  XOR2_X1 U822 ( .A(G101), .B(n778), .Z(G3) );
endmodule

