//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986;
  AOI21_X1  g000(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT74), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(KEYINPUT74), .ZN(new_n204));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n203), .A2(new_n207), .A3(new_n204), .A4(new_n205), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT26), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT67), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n216), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(new_n213), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n214), .A2(new_n215), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT27), .B(G183gat), .ZN(new_n220));
  INV_X1    g019(.A(G190gat), .ZN(new_n221));
  OR2_X1    g020(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n222));
  NAND2_X1  g021(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT27), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT27), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G183gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n228), .A3(new_n221), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n222), .A2(new_n223), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n219), .A2(new_n224), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G226gat), .ZN(new_n234));
  INV_X1    g033(.A(G233gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n232), .A2(KEYINPUT24), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT24), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(G183gat), .A3(G190gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n221), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT23), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n245), .A2(G169gat), .A3(G176gat), .ZN(new_n246));
  INV_X1    g045(.A(new_n215), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n244), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n245), .B1(G169gat), .B2(G176gat), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n249), .A2(KEYINPUT25), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n212), .A2(KEYINPUT23), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT65), .A3(new_n215), .ZN(new_n252));
  AND4_X1   g051(.A1(new_n243), .A2(new_n248), .A3(new_n250), .A4(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(new_n225), .A3(new_n221), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n251), .A2(new_n249), .A3(new_n215), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT25), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n233), .B(new_n237), .C1(new_n253), .C2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n236), .A2(KEYINPUT29), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n243), .A2(new_n248), .A3(new_n250), .A4(new_n252), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n251), .A2(new_n249), .A3(new_n215), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n256), .A2(new_n254), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n264), .B1(new_n266), .B2(new_n241), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n263), .B1(new_n267), .B2(KEYINPUT25), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n262), .B1(new_n268), .B2(new_n233), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n211), .B1(new_n261), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n209), .A2(new_n210), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT25), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n225), .A2(KEYINPUT24), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n273), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n232), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(new_n265), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n272), .B1(new_n275), .B2(new_n264), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n232), .B1(new_n229), .B2(new_n230), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n220), .A2(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n276), .A2(new_n263), .B1(new_n279), .B2(new_n219), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n271), .B(new_n260), .C1(new_n280), .C2(new_n262), .ZN(new_n281));
  XNOR2_X1  g080(.A(G8gat), .B(G36gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT75), .ZN(new_n283));
  XNOR2_X1  g082(.A(G64gat), .B(G92gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT30), .ZN(new_n288));
  INV_X1    g087(.A(new_n281), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n233), .B1(new_n253), .B2(new_n259), .ZN(new_n290));
  INV_X1    g089(.A(new_n262), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n271), .B1(new_n292), .B2(new_n260), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n285), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(KEYINPUT76), .B(new_n285), .C1(new_n289), .C2(new_n293), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n288), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n300));
  INV_X1    g099(.A(G120gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G113gat), .ZN(new_n302));
  INV_X1    g101(.A(G113gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G120gat), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT1), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  OR2_X1    g104(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n306));
  AND2_X1   g105(.A1(G127gat), .A2(G134gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(G127gat), .A2(G134gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n305), .A2(new_n309), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n300), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G141gat), .B(G148gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n317), .B1(G155gat), .B2(G162gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n315), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G141gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G148gat), .ZN(new_n321));
  INV_X1    g120(.A(G148gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G141gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G155gat), .B(G162gat), .ZN(new_n325));
  INV_X1    g124(.A(G155gat), .ZN(new_n326));
  INV_X1    g125(.A(G162gat), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT2), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n324), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n319), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G127gat), .B(G134gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n306), .B(new_n332), .C1(new_n333), .C2(KEYINPUT1), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n305), .A2(new_n309), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT69), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n312), .A2(KEYINPUT4), .A3(new_n331), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n335), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(new_n319), .A3(new_n329), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n342));
  INV_X1    g141(.A(new_n338), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n319), .A2(new_n329), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n337), .A2(new_n341), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT5), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n330), .A2(new_n335), .A3(new_n334), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n339), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n347), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n312), .A2(new_n331), .A3(new_n336), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n340), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n344), .B1(new_n319), .B2(new_n329), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(new_n338), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n352), .B1(new_n358), .B2(new_n345), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n331), .A2(KEYINPUT4), .A3(new_n338), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n356), .A2(new_n359), .A3(new_n349), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(G1gat), .B(G29gat), .Z(new_n363));
  XNOR2_X1  g162(.A(G57gat), .B(G85gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n362), .A2(KEYINPUT6), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n367), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n361), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT6), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n360), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n373), .B1(new_n340), .B2(new_n355), .ZN(new_n374));
  AOI211_X1 g173(.A(KEYINPUT5), .B(new_n352), .C1(new_n358), .C2(new_n345), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n374), .A2(new_n375), .B1(new_n348), .B2(new_n353), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT78), .B1(new_n376), .B2(new_n369), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n378), .A3(new_n367), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n372), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n368), .B1(new_n380), .B2(KEYINPUT79), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT6), .B1(new_n376), .B2(new_n369), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n378), .B1(new_n362), .B2(new_n367), .ZN(new_n383));
  AOI211_X1 g182(.A(KEYINPUT78), .B(new_n369), .C1(new_n354), .C2(new_n361), .ZN(new_n384));
  OAI211_X1 g183(.A(KEYINPUT79), .B(new_n382), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n299), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT29), .B1(new_n209), .B2(new_n210), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n330), .B1(new_n388), .B2(KEYINPUT3), .ZN(new_n389));
  INV_X1    g188(.A(new_n345), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n211), .B1(KEYINPUT29), .B2(new_n390), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n389), .A2(new_n391), .A3(G22gat), .ZN(new_n392));
  AOI21_X1  g191(.A(G22gat), .B1(new_n389), .B2(new_n391), .ZN(new_n393));
  OAI211_X1 g192(.A(G228gat), .B(G233gat), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n389), .A2(new_n391), .ZN(new_n395));
  INV_X1    g194(.A(G22gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G228gat), .A2(G233gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n389), .A2(new_n391), .A3(G22gat), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G78gat), .B(G106gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT31), .B(G50gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT80), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n404), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(KEYINPUT80), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n394), .A2(new_n408), .A3(new_n400), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT81), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT81), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n406), .A2(new_n412), .A3(new_n409), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n387), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT37), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT84), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n271), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n417), .B1(new_n293), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n270), .A2(new_n418), .A3(new_n281), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n270), .A2(new_n417), .A3(new_n281), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT38), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n424), .A3(new_n285), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n416), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n423), .A2(new_n285), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n421), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n427), .A2(KEYINPUT85), .A3(new_n428), .A4(new_n424), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT83), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(new_n376), .B2(new_n369), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n362), .A2(KEYINPUT83), .A3(new_n367), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n382), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n287), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT37), .B1(new_n289), .B2(new_n293), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(new_n285), .A3(new_n423), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n435), .B1(new_n437), .B2(KEYINPUT38), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n430), .A2(new_n368), .A3(new_n434), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n432), .A2(new_n433), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(new_n298), .B2(new_n288), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT39), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n356), .A2(new_n346), .A3(new_n360), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT82), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n443), .A2(new_n444), .A3(new_n352), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n443), .B2(new_n352), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n352), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT82), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n443), .A2(new_n444), .A3(new_n352), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n351), .A2(new_n352), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(new_n442), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n447), .A2(new_n453), .A3(new_n369), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT40), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n447), .A2(new_n453), .A3(KEYINPUT40), .A4(new_n369), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n406), .A2(new_n409), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n439), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  XOR2_X1   g259(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n461));
  NAND2_X1  g260(.A1(G227gat), .A2(G233gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n312), .A2(new_n336), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n290), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n268), .A2(new_n233), .B1(new_n312), .B2(new_n336), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT32), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT33), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(G71gat), .B(G99gat), .Z(new_n471));
  XNOR2_X1  g270(.A(G15gat), .B(G43gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n468), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT32), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n290), .A2(new_n464), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n268), .A2(new_n336), .A3(new_n312), .A4(new_n233), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n475), .B1(new_n478), .B2(new_n463), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n473), .A2(KEYINPUT33), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT70), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n462), .B1(new_n476), .B2(new_n477), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT70), .ZN(new_n483));
  INV_X1    g282(.A(new_n480), .ZN(new_n484));
  NOR4_X1   g283(.A1(new_n482), .A2(new_n483), .A3(new_n475), .A4(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n474), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT34), .B1(new_n478), .B2(new_n463), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT34), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n476), .A2(new_n477), .A3(new_n488), .A4(new_n462), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT71), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n489), .A2(KEYINPUT71), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n486), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n491), .A2(new_n492), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n467), .A2(KEYINPUT32), .A3(new_n480), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n483), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n479), .A2(KEYINPUT70), .A3(new_n480), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n495), .B1(new_n499), .B2(new_n474), .ZN(new_n500));
  OAI211_X1 g299(.A(KEYINPUT73), .B(new_n461), .C1(new_n494), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n493), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n499), .A2(new_n495), .A3(new_n474), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(KEYINPUT36), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n502), .A2(new_n503), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT73), .B1(new_n506), .B2(new_n461), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n415), .B(new_n460), .C1(new_n505), .C2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n459), .A2(new_n503), .A3(new_n502), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT35), .B1(new_n387), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n506), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT35), .B1(new_n434), .B2(new_n368), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n511), .A2(new_n299), .A3(new_n459), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT86), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT86), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n508), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519));
  OR2_X1    g318(.A1(G43gat), .A2(G50gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(G43gat), .A2(G50gat), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT87), .B(G50gat), .Z(new_n523));
  OAI211_X1 g322(.A(new_n519), .B(new_n521), .C1(new_n523), .C2(G43gat), .ZN(new_n524));
  INV_X1    g323(.A(G29gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n526));
  XOR2_X1   g325(.A(KEYINPUT14), .B(G29gat), .Z(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(G36gat), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n522), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n528), .A2(new_n522), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(G1gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT16), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(G1gat), .B2(new_n532), .ZN(new_n536));
  INV_X1    g335(.A(G8gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n529), .A2(new_n530), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT17), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n539), .B1(new_n541), .B2(new_n538), .ZN(new_n542));
  NAND2_X1  g341(.A1(G229gat), .A2(G233gat), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n544), .A2(KEYINPUT18), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n542), .A2(KEYINPUT18), .A3(new_n543), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n531), .B(new_n538), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n543), .B(KEYINPUT13), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n545), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G197gat), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT11), .B(G169gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT12), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n555), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n545), .A2(new_n557), .A3(new_n546), .A4(new_n549), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n516), .A2(new_n518), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(G57gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(G64gat), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n562), .A2(KEYINPUT88), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(KEYINPUT88), .ZN(new_n564));
  INV_X1    g363(.A(G64gat), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n563), .B(new_n564), .C1(G57gat), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G71gat), .A2(G78gat), .ZN(new_n567));
  OR2_X1    g366(.A1(G71gat), .A2(G78gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT9), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n565), .A2(G57gat), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT9), .B1(new_n562), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(new_n567), .A3(new_n568), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT21), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G127gat), .B(G155gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT20), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n579), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G183gat), .B(G211gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n538), .B1(new_n575), .B2(new_n576), .ZN(new_n585));
  XOR2_X1   g384(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n584), .A2(new_n587), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT90), .B(KEYINPUT7), .ZN(new_n592));
  INV_X1    g391(.A(G85gat), .ZN(new_n593));
  INV_X1    g392(.A(G92gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n595), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n598), .B1(new_n593), .B2(new_n594), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G99gat), .B(G106gat), .Z(new_n601));
  OR2_X1    g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT41), .ZN(new_n605));
  NAND2_X1  g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606));
  OAI22_X1  g405(.A1(new_n604), .A2(new_n531), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(new_n541), .B2(new_n604), .ZN(new_n608));
  XNOR2_X1  g407(.A(G190gat), .B(G218gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n605), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT91), .Z(new_n614));
  OR2_X1    g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(KEYINPUT91), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n575), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n602), .A2(new_n571), .A3(new_n574), .A4(new_n603), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n624), .A2(new_n623), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n621), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n620), .B1(new_n622), .B2(new_n624), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G120gat), .B(G148gat), .Z(new_n630));
  XNOR2_X1  g429(.A(G176gat), .B(G204gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT92), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n629), .A2(new_n632), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n591), .A2(new_n619), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n560), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n381), .A2(new_n386), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n533), .ZN(G1324gat));
  NOR2_X1   g443(.A1(new_n640), .A2(new_n299), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT16), .B(G8gat), .Z(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(new_n537), .B2(new_n645), .ZN(new_n648));
  MUX2_X1   g447(.A(new_n647), .B(new_n648), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g448(.A(KEYINPUT93), .B1(new_n505), .B2(new_n507), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n461), .B1(new_n494), .B2(new_n500), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT73), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT93), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n654), .A2(new_n655), .A3(new_n504), .A4(new_n501), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(G15gat), .B1(new_n640), .B2(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n506), .A2(G15gat), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n640), .B2(new_n660), .ZN(G1326gat));
  INV_X1    g460(.A(new_n414), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n640), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT94), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT43), .B(G22gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  NAND3_X1  g465(.A1(new_n516), .A2(new_n518), .A3(new_n618), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT44), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n438), .A2(new_n368), .A3(new_n434), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n410), .B1(new_n669), .B2(new_n430), .ZN(new_n670));
  AOI22_X1  g469(.A1(new_n670), .A2(new_n458), .B1(new_n387), .B2(new_n414), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n650), .A2(new_n671), .A3(new_n656), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n514), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674));
  AND4_X1   g473(.A1(KEYINPUT96), .A2(new_n673), .A3(new_n674), .A4(new_n618), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n619), .B1(new_n672), .B2(new_n514), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT96), .B1(new_n676), .B2(new_n674), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n668), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n559), .B(KEYINPUT95), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n637), .A2(new_n590), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n525), .B1(new_n682), .B2(new_n641), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n680), .A2(new_n619), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n560), .A2(new_n525), .A3(new_n641), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT45), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT97), .ZN(G1328gat));
  NAND2_X1  g488(.A1(new_n678), .A2(new_n681), .ZN(new_n690));
  OAI21_X1  g489(.A(G36gat), .B1(new_n690), .B2(new_n299), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n560), .A2(new_n684), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(G36gat), .A3(new_n299), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(KEYINPUT98), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT98), .B(KEYINPUT46), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n691), .B(new_n695), .C1(new_n693), .C2(new_n696), .ZN(G1329gat));
  NOR2_X1   g496(.A1(new_n506), .A2(G43gat), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n560), .A2(new_n684), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT99), .ZN(new_n700));
  INV_X1    g499(.A(new_n658), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n682), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G43gat), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n702), .A2(new_n703), .ZN(new_n706));
  OAI211_X1 g505(.A(KEYINPUT47), .B(new_n700), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT100), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n702), .A2(G43gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n700), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AOI211_X1 g511(.A(KEYINPUT100), .B(KEYINPUT47), .C1(new_n709), .C2(new_n700), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n707), .B1(new_n712), .B2(new_n713), .ZN(G1330gat));
  OAI21_X1  g513(.A(new_n523), .B1(new_n690), .B2(new_n459), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n692), .A2(new_n662), .A3(new_n523), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT48), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n523), .B1(new_n690), .B2(new_n662), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n722), .A2(new_n723), .A3(new_n716), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n719), .B1(new_n724), .B2(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g524(.A1(new_n556), .A2(new_n558), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT95), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT95), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n559), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NOR4_X1   g529(.A1(new_n730), .A2(new_n590), .A3(new_n618), .A4(new_n637), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n673), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n642), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(new_n561), .ZN(G1332gat));
  INV_X1    g533(.A(new_n732), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n299), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT103), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1333gat));
  NOR3_X1   g539(.A1(new_n732), .A2(G71gat), .A3(new_n506), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n735), .A2(new_n701), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(G71gat), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g543(.A1(new_n735), .A2(new_n414), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g545(.A1(new_n730), .A2(new_n591), .A3(new_n637), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n678), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(G85gat), .B1(new_n748), .B2(new_n642), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n730), .A2(new_n591), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n676), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n751), .A2(new_n752), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n636), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n641), .A2(new_n593), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n749), .B1(new_n756), .B2(new_n757), .ZN(G1336gat));
  NOR3_X1   g557(.A1(new_n756), .A2(G92gat), .A3(new_n299), .ZN(new_n759));
  INV_X1    g558(.A(new_n748), .ZN(new_n760));
  INV_X1    g559(.A(new_n299), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n759), .B1(G92gat), .B2(new_n762), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT52), .Z(G1337gat));
  OR3_X1    g563(.A1(new_n756), .A2(G99gat), .A3(new_n506), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n760), .A2(new_n701), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT104), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G99gat), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n766), .A2(KEYINPUT104), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n765), .B1(new_n768), .B2(new_n769), .ZN(G1338gat));
  NOR2_X1   g569(.A1(new_n459), .A2(G106gat), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n755), .ZN(new_n773));
  AOI211_X1 g572(.A(new_n637), .B(new_n772), .C1(new_n773), .C2(new_n753), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776));
  OAI21_X1  g575(.A(G106gat), .B1(new_n748), .B2(new_n459), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT106), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n678), .A2(new_n414), .A3(new_n747), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G106gat), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n774), .B1(new_n781), .B2(KEYINPUT105), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT105), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n780), .A2(new_n783), .A3(G106gat), .ZN(new_n784));
  AOI211_X1 g583(.A(new_n779), .B(new_n776), .C1(new_n782), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n781), .A2(KEYINPUT105), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(new_n784), .A3(new_n775), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT106), .B1(new_n787), .B2(KEYINPUT53), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n778), .B1(new_n785), .B2(new_n788), .ZN(G1339gat));
  NOR2_X1   g588(.A1(new_n730), .A2(new_n638), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n625), .A2(new_n626), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n620), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n625), .A2(new_n626), .A3(new_n621), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(KEYINPUT54), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n632), .B1(new_n627), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n794), .A2(KEYINPUT55), .A3(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n634), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n794), .A2(new_n796), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n802), .B1(new_n727), .B2(new_n729), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n547), .A2(new_n548), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT107), .Z(new_n805));
  NOR2_X1   g604(.A1(new_n542), .A2(new_n543), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n554), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n558), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n636), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT109), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n809), .A2(KEYINPUT109), .A3(new_n636), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n619), .B1(new_n803), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n808), .B(KEYINPUT108), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n798), .A2(new_n801), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n816), .A2(new_n817), .A3(new_n618), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n790), .B1(new_n820), .B2(new_n590), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n414), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n511), .A2(new_n299), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n642), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n825), .A2(new_n303), .A3(new_n726), .ZN(new_n826));
  INV_X1    g625(.A(new_n790), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n812), .B(new_n813), .C1(new_n679), .C2(new_n802), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n818), .B1(new_n828), .B2(new_n619), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n829), .B2(new_n591), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n823), .A2(new_n410), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n641), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(G113gat), .B1(new_n833), .B2(new_n730), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n826), .A2(new_n834), .ZN(G1340gat));
  NOR3_X1   g634(.A1(new_n825), .A2(new_n301), .A3(new_n637), .ZN(new_n836));
  AOI21_X1  g635(.A(G120gat), .B1(new_n833), .B2(new_n636), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(G1341gat));
  OAI21_X1  g637(.A(G127gat), .B1(new_n825), .B2(new_n590), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n590), .A2(G127gat), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n832), .B2(new_n840), .ZN(G1342gat));
  NOR3_X1   g640(.A1(new_n832), .A2(G134gat), .A3(new_n619), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT110), .ZN(new_n846));
  INV_X1    g645(.A(new_n825), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n618), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n848), .B2(G134gat), .ZN(new_n849));
  INV_X1    g648(.A(G134gat), .ZN(new_n850));
  AOI211_X1 g649(.A(KEYINPUT110), .B(new_n850), .C1(new_n847), .C2(new_n618), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n844), .B(new_n845), .C1(new_n849), .C2(new_n851), .ZN(G1343gat));
  NOR2_X1   g651(.A1(new_n642), .A2(new_n761), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n701), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT111), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT55), .B1(new_n799), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n794), .A2(KEYINPUT111), .A3(new_n796), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(KEYINPUT112), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT112), .B1(new_n857), .B2(new_n858), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n798), .B(KEYINPUT113), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n559), .ZN(new_n863));
  INV_X1    g662(.A(new_n861), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n859), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT113), .B1(new_n865), .B2(new_n798), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n810), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n818), .B1(new_n867), .B2(new_n619), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n827), .B1(new_n868), .B2(new_n591), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n662), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(KEYINPUT114), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n821), .B2(new_n459), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT114), .B1(new_n869), .B2(new_n871), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n559), .B(new_n855), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G141gat), .ZN(new_n877));
  XOR2_X1   g676(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n878));
  OAI21_X1  g677(.A(KEYINPUT115), .B1(new_n821), .B2(new_n642), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n830), .A2(new_n880), .A3(new_n641), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n658), .A2(new_n410), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(new_n761), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n879), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n726), .A2(G141gat), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n878), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n877), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n730), .B(new_n855), .C1(new_n874), .C2(new_n875), .ZN(new_n888));
  AOI22_X1  g687(.A1(new_n888), .A2(G141gat), .B1(new_n884), .B2(new_n885), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(G1344gat));
  NAND3_X1  g690(.A1(new_n884), .A2(new_n322), .A3(new_n636), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(G148gat), .ZN(new_n894));
  INV_X1    g693(.A(new_n855), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n872), .A2(new_n873), .ZN(new_n896));
  INV_X1    g695(.A(new_n875), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n894), .B1(new_n898), .B2(new_n636), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n867), .A2(new_n619), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n798), .A2(new_n618), .A3(new_n801), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n901), .A2(KEYINPUT118), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(KEYINPUT118), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n816), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n591), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n638), .A2(new_n559), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n870), .B(new_n414), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT57), .B1(new_n821), .B2(new_n459), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n636), .B1(new_n855), .B2(KEYINPUT117), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(KEYINPUT117), .B2(new_n855), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n893), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n892), .B1(new_n899), .B2(new_n913), .ZN(G1345gat));
  NAND2_X1  g713(.A1(new_n591), .A2(G155gat), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT119), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n855), .B(new_n916), .C1(new_n874), .C2(new_n875), .ZN(new_n917));
  AND4_X1   g716(.A1(new_n591), .A2(new_n879), .A3(new_n881), .A4(new_n883), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(G155gat), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n917), .B(KEYINPUT120), .C1(new_n918), .C2(G155gat), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1346gat));
  AOI21_X1  g722(.A(G162gat), .B1(new_n884), .B2(new_n618), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n619), .A2(new_n327), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n898), .B2(new_n925), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n641), .A2(new_n299), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n511), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT121), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n822), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(G169gat), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n930), .A2(new_n931), .A3(new_n726), .ZN(new_n932));
  NOR4_X1   g731(.A1(new_n821), .A2(new_n641), .A3(new_n299), .A4(new_n509), .ZN(new_n933));
  AOI21_X1  g732(.A(G169gat), .B1(new_n933), .B2(new_n730), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n932), .A2(new_n934), .ZN(G1348gat));
  OAI21_X1  g734(.A(G176gat), .B1(new_n930), .B2(new_n637), .ZN(new_n936));
  INV_X1    g735(.A(G176gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n933), .A2(new_n937), .A3(new_n636), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1349gat));
  AND2_X1   g738(.A1(new_n591), .A2(new_n220), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n933), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n830), .A2(new_n662), .A3(new_n591), .A4(new_n929), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(G183gat), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n944), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n946));
  AOI22_X1  g745(.A1(new_n933), .A2(new_n940), .B1(new_n942), .B2(G183gat), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT60), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n950), .B1(new_n944), .B2(KEYINPUT60), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n947), .A2(KEYINPUT122), .A3(new_n948), .ZN(new_n952));
  OAI22_X1  g751(.A1(new_n945), .A2(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n933), .A2(new_n221), .A3(new_n618), .ZN(new_n954));
  OAI21_X1  g753(.A(G190gat), .B1(new_n930), .B2(new_n619), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n955), .A2(KEYINPUT61), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(KEYINPUT61), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(G1351gat));
  NAND2_X1  g757(.A1(new_n658), .A2(new_n927), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT124), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n909), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(G197gat), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n961), .A2(new_n962), .A3(new_n726), .ZN(new_n963));
  NOR4_X1   g762(.A1(new_n821), .A2(new_n641), .A3(new_n299), .A4(new_n882), .ZN(new_n964));
  AOI21_X1  g763(.A(G197gat), .B1(new_n964), .B2(new_n730), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n963), .A2(new_n965), .ZN(G1352gat));
  OAI21_X1  g765(.A(G204gat), .B1(new_n961), .B2(new_n637), .ZN(new_n967));
  INV_X1    g766(.A(G204gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n964), .A2(new_n968), .A3(new_n636), .ZN(new_n969));
  AND2_X1   g768(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n970));
  NOR2_X1   g769(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n967), .B(new_n972), .C1(new_n970), .C2(new_n969), .ZN(G1353gat));
  INV_X1    g772(.A(G211gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n964), .A2(new_n974), .A3(new_n591), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n909), .A2(new_n591), .A3(new_n960), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n976), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT63), .B1(new_n976), .B2(G211gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(G1354gat));
  AOI21_X1  g778(.A(G218gat), .B1(new_n964), .B2(new_n618), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n909), .A2(KEYINPUT126), .A3(new_n960), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n618), .A2(G218gat), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT127), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n961), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n980), .B1(new_n984), .B2(new_n986), .ZN(G1355gat));
endmodule


