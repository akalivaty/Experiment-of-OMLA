

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761;

  OR2_X1 U371 ( .A1(n637), .A2(G902), .ZN(n503) );
  XNOR2_X1 U372 ( .A(n429), .B(G107), .ZN(n484) );
  INV_X1 U373 ( .A(G104), .ZN(n428) );
  AND2_X1 U374 ( .A1(n553), .A2(n422), .ZN(n374) );
  NOR2_X1 U375 ( .A1(n659), .A2(n577), .ZN(n564) );
  BUF_X1 U376 ( .A(n649), .Z(n727) );
  XNOR2_X1 U377 ( .A(n406), .B(n405), .ZN(n607) );
  AND2_X1 U378 ( .A1(n545), .A2(n375), .ZN(n349) );
  OR2_X2 U379 ( .A1(n692), .A2(n533), .ZN(n358) );
  XNOR2_X2 U380 ( .A(n732), .B(n470), .ZN(n644) );
  XNOR2_X2 U381 ( .A(n462), .B(n461), .ZN(n732) );
  XNOR2_X2 U382 ( .A(n349), .B(KEYINPUT32), .ZN(n757) );
  NOR2_X1 U383 ( .A1(n533), .A2(n508), .ZN(n377) );
  XNOR2_X1 U384 ( .A(n377), .B(n376), .ZN(n541) );
  INV_X1 U385 ( .A(n669), .ZN(n574) );
  XNOR2_X1 U386 ( .A(n518), .B(n517), .ZN(n528) );
  INV_X1 U387 ( .A(n460), .ZN(n461) );
  XNOR2_X1 U388 ( .A(n402), .B(n401), .ZN(n460) );
  INV_X1 U389 ( .A(KEYINPUT35), .ZN(n354) );
  INV_X2 U390 ( .A(G953), .ZN(n746) );
  INV_X1 U391 ( .A(KEYINPUT22), .ZN(n376) );
  INV_X1 U392 ( .A(KEYINPUT4), .ZN(n352) );
  INV_X2 U393 ( .A(G131), .ZN(n373) );
  AND2_X1 U394 ( .A1(n655), .A2(n620), .ZN(n625) );
  XNOR2_X1 U395 ( .A(n420), .B(n419), .ZN(n418) );
  XNOR2_X1 U396 ( .A(n358), .B(n534), .ZN(n357) );
  NOR2_X1 U397 ( .A1(n595), .A2(n594), .ZN(n608) );
  NOR2_X1 U398 ( .A1(n541), .A2(n542), .ZN(n545) );
  AND2_X1 U399 ( .A1(n564), .A2(n563), .ZN(n565) );
  AND2_X1 U400 ( .A1(n544), .A2(n416), .ZN(n375) );
  INV_X1 U401 ( .A(n605), .ZN(n356) );
  XNOR2_X1 U402 ( .A(n417), .B(n524), .ZN(n596) );
  NAND2_X1 U403 ( .A1(n381), .A2(n380), .ZN(n659) );
  NAND2_X1 U404 ( .A1(n676), .A2(n380), .ZN(n508) );
  NOR2_X1 U405 ( .A1(n574), .A2(n597), .ZN(n576) );
  INV_X1 U406 ( .A(n662), .ZN(n381) );
  NAND2_X2 U407 ( .A1(n555), .A2(n679), .ZN(n600) );
  XNOR2_X1 U408 ( .A(n458), .B(n457), .ZN(n662) );
  XNOR2_X1 U409 ( .A(n528), .B(n519), .ZN(n540) );
  NOR2_X1 U410 ( .A1(G902), .A2(n728), .ZN(n458) );
  XNOR2_X1 U411 ( .A(n450), .B(n449), .ZN(n728) );
  XNOR2_X1 U412 ( .A(n516), .B(n515), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n427), .B(n424), .ZN(n462) );
  XNOR2_X1 U414 ( .A(n484), .B(n489), .ZN(n427) );
  XNOR2_X1 U415 ( .A(n459), .B(n425), .ZN(n424) );
  XNOR2_X1 U416 ( .A(n352), .B(KEYINPUT65), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n426), .B(G110), .ZN(n459) );
  INV_X1 U418 ( .A(KEYINPUT45), .ZN(n384) );
  INV_X2 U419 ( .A(G128), .ZN(n353) );
  OR2_X2 U420 ( .A1(n350), .A2(G902), .ZN(n518) );
  XNOR2_X1 U421 ( .A(n350), .B(n650), .ZN(n651) );
  XNOR2_X2 U422 ( .A(n480), .B(n351), .ZN(n469) );
  XNOR2_X2 U423 ( .A(n353), .B(G143), .ZN(n480) );
  XNOR2_X2 U424 ( .A(n355), .B(n354), .ZN(n755) );
  NAND2_X1 U425 ( .A1(n357), .A2(n356), .ZN(n355) );
  XNOR2_X2 U426 ( .A(n744), .B(G146), .ZN(n516) );
  NOR2_X1 U427 ( .A1(n597), .A2(n596), .ZN(n599) );
  XNOR2_X1 U428 ( .A(n532), .B(KEYINPUT33), .ZN(n692) );
  NOR2_X1 U429 ( .A1(n531), .A2(n530), .ZN(n532) );
  OR2_X1 U430 ( .A1(G237), .A2(G902), .ZN(n473) );
  INV_X1 U431 ( .A(G116), .ZN(n429) );
  AND2_X1 U432 ( .A1(n635), .A2(n713), .ZN(n363) );
  INV_X1 U433 ( .A(KEYINPUT79), .ZN(n453) );
  INV_X1 U434 ( .A(n591), .ZN(n388) );
  INV_X1 U435 ( .A(G119), .ZN(n426) );
  XNOR2_X1 U436 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n440) );
  XNOR2_X1 U437 ( .A(G113), .B(KEYINPUT95), .ZN(n497) );
  XNOR2_X1 U438 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n498) );
  INV_X1 U439 ( .A(G140), .ZN(n492) );
  XNOR2_X1 U440 ( .A(n439), .B(n464), .ZN(n490) );
  XNOR2_X1 U441 ( .A(KEYINPUT96), .B(G143), .ZN(n495) );
  INV_X1 U442 ( .A(G134), .ZN(n431) );
  INV_X1 U443 ( .A(KEYINPUT30), .ZN(n365) );
  INV_X1 U444 ( .A(n572), .ZN(n563) );
  XNOR2_X1 U445 ( .A(n488), .B(G478), .ZN(n583) );
  XNOR2_X1 U446 ( .A(n433), .B(n400), .ZN(n399) );
  XNOR2_X1 U447 ( .A(G137), .B(G119), .ZN(n433) );
  XNOR2_X1 U448 ( .A(G116), .B(KEYINPUT5), .ZN(n400) );
  NOR2_X2 U449 ( .A1(G953), .A2(G237), .ZN(n491) );
  XNOR2_X1 U450 ( .A(KEYINPUT73), .B(KEYINPUT3), .ZN(n401) );
  XNOR2_X1 U451 ( .A(n403), .B(G113), .ZN(n402) );
  INV_X1 U452 ( .A(G101), .ZN(n403) );
  XNOR2_X1 U453 ( .A(G134), .B(G122), .ZN(n485) );
  XNOR2_X1 U454 ( .A(G101), .B(G104), .ZN(n509) );
  XOR2_X1 U455 ( .A(G110), .B(G107), .Z(n510) );
  INV_X1 U456 ( .A(KEYINPUT105), .ZN(n369) );
  XNOR2_X1 U457 ( .A(n404), .B(KEYINPUT39), .ZN(n570) );
  NAND2_X1 U458 ( .A1(n416), .A2(n413), .ZN(n412) );
  NAND2_X1 U459 ( .A1(n600), .A2(n603), .ZN(n413) );
  OR2_X1 U460 ( .A1(n626), .A2(G902), .ZN(n437) );
  INV_X1 U461 ( .A(KEYINPUT0), .ZN(n430) );
  INV_X1 U462 ( .A(KEYINPUT72), .ZN(n397) );
  INV_X1 U463 ( .A(KEYINPUT48), .ZN(n393) );
  NAND2_X1 U464 ( .A1(n550), .A2(n549), .ZN(n422) );
  NAND2_X1 U465 ( .A1(G234), .A2(G237), .ZN(n474) );
  XNOR2_X1 U466 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U467 ( .A(n454), .B(n453), .ZN(n455) );
  AND2_X1 U468 ( .A1(n392), .A2(n385), .ZN(n420) );
  XNOR2_X1 U469 ( .A(n387), .B(n386), .ZN(n385) );
  INV_X1 U470 ( .A(KEYINPUT101), .ZN(n386) );
  INV_X1 U471 ( .A(KEYINPUT102), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n382), .B(KEYINPUT76), .ZN(n531) );
  XNOR2_X1 U473 ( .A(KEYINPUT15), .B(G902), .ZN(n619) );
  INV_X1 U474 ( .A(n583), .ZN(n523) );
  BUF_X1 U475 ( .A(n662), .Z(n372) );
  INV_X1 U476 ( .A(KEYINPUT16), .ZN(n425) );
  XNOR2_X1 U477 ( .A(G128), .B(KEYINPUT24), .ZN(n442) );
  XNOR2_X1 U478 ( .A(n490), .B(n512), .ZN(n743) );
  XNOR2_X1 U479 ( .A(n407), .B(n501), .ZN(n637) );
  XNOR2_X1 U480 ( .A(n371), .B(n370), .ZN(n657) );
  INV_X1 U481 ( .A(KEYINPUT84), .ZN(n370) );
  XNOR2_X1 U482 ( .A(n585), .B(KEYINPUT41), .ZN(n693) );
  INV_X1 U483 ( .A(KEYINPUT78), .ZN(n405) );
  XNOR2_X1 U484 ( .A(n557), .B(n365), .ZN(n364) );
  INV_X1 U485 ( .A(KEYINPUT19), .ZN(n367) );
  XNOR2_X1 U486 ( .A(n460), .B(n399), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n487), .B(n379), .ZN(n723) );
  XNOR2_X1 U488 ( .A(n486), .B(n359), .ZN(n379) );
  NOR2_X1 U489 ( .A1(n614), .A2(n555), .ZN(n722) );
  NAND2_X1 U490 ( .A1(n570), .A2(n714), .ZN(n571) );
  AND2_X1 U491 ( .A1(n601), .A2(n415), .ZN(n414) );
  INV_X1 U492 ( .A(KEYINPUT34), .ZN(n534) );
  INV_X1 U493 ( .A(n663), .ZN(n380) );
  XOR2_X1 U494 ( .A(KEYINPUT98), .B(KEYINPUT9), .Z(n359) );
  INV_X1 U495 ( .A(n660), .ZN(n416) );
  XOR2_X1 U496 ( .A(G137), .B(G140), .Z(n512) );
  AND2_X1 U497 ( .A1(n618), .A2(n621), .ZN(n360) );
  XOR2_X1 U498 ( .A(n626), .B(KEYINPUT62), .Z(n361) );
  XOR2_X1 U499 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n362) );
  NOR2_X1 U500 ( .A1(n700), .A2(G953), .ZN(n702) );
  XNOR2_X1 U501 ( .A(n446), .B(n743), .ZN(n450) );
  NAND2_X1 U502 ( .A1(n608), .A2(n363), .ZN(n398) );
  NAND2_X1 U503 ( .A1(n565), .A2(n364), .ZN(n406) );
  NOR2_X1 U504 ( .A1(n411), .A2(n412), .ZN(n410) );
  XNOR2_X1 U505 ( .A(n366), .B(n393), .ZN(n616) );
  NAND2_X1 U506 ( .A1(n394), .A2(n396), .ZN(n366) );
  NAND2_X1 U507 ( .A1(n383), .A2(n540), .ZN(n382) );
  NOR2_X1 U508 ( .A1(n755), .A2(n537), .ZN(n551) );
  XNOR2_X2 U509 ( .A(n600), .B(n367), .ZN(n588) );
  XNOR2_X1 U510 ( .A(n581), .B(KEYINPUT97), .ZN(n522) );
  NAND2_X1 U511 ( .A1(n368), .A2(n660), .ZN(n612) );
  XNOR2_X1 U512 ( .A(n611), .B(n369), .ZN(n368) );
  XNOR2_X1 U513 ( .A(n408), .B(n490), .ZN(n407) );
  NAND2_X1 U514 ( .A1(n745), .A2(n656), .ZN(n371) );
  XNOR2_X2 U515 ( .A(n373), .B(KEYINPUT71), .ZN(n496) );
  NAND2_X1 U516 ( .A1(n374), .A2(n423), .ZN(n421) );
  NOR2_X2 U517 ( .A1(n588), .A2(n478), .ZN(n479) );
  NOR2_X4 U518 ( .A1(n589), .A2(n588), .ZN(n715) );
  XNOR2_X2 U519 ( .A(n579), .B(n580), .ZN(n589) );
  XNOR2_X1 U520 ( .A(n398), .B(n397), .ZN(n396) );
  NOR2_X1 U521 ( .A1(n602), .A2(n415), .ZN(n411) );
  NAND2_X1 U522 ( .A1(n378), .A2(n656), .ZN(n624) );
  NAND2_X1 U523 ( .A1(n622), .A2(n623), .ZN(n378) );
  NAND2_X1 U524 ( .A1(n410), .A2(n409), .ZN(n635) );
  NAND2_X1 U525 ( .A1(n522), .A2(n583), .ZN(n417) );
  INV_X1 U526 ( .A(n659), .ZN(n383) );
  NAND2_X1 U527 ( .A1(n623), .A2(n360), .ZN(n655) );
  OR2_X1 U528 ( .A1(n623), .A2(KEYINPUT2), .ZN(n654) );
  AND2_X1 U529 ( .A1(n623), .A2(n746), .ZN(n739) );
  XNOR2_X2 U530 ( .A(n554), .B(n384), .ZN(n623) );
  NAND2_X1 U531 ( .A1(n389), .A2(n388), .ZN(n387) );
  NAND2_X1 U532 ( .A1(n391), .A2(n390), .ZN(n389) );
  INV_X1 U533 ( .A(n705), .ZN(n390) );
  INV_X1 U534 ( .A(n720), .ZN(n391) );
  INV_X1 U535 ( .A(n703), .ZN(n392) );
  XNOR2_X1 U536 ( .A(n395), .B(n362), .ZN(n394) );
  NAND2_X1 U537 ( .A1(n758), .A2(n760), .ZN(n395) );
  NAND2_X1 U538 ( .A1(n607), .A2(n680), .ZN(n404) );
  XNOR2_X2 U539 ( .A(n469), .B(n432), .ZN(n744) );
  AND2_X2 U540 ( .A1(n625), .A2(n624), .ZN(n649) );
  XNOR2_X1 U541 ( .A(n494), .B(n489), .ZN(n408) );
  NAND2_X1 U542 ( .A1(n602), .A2(n414), .ZN(n409) );
  INV_X1 U543 ( .A(n603), .ZN(n415) );
  NOR2_X2 U544 ( .A1(n421), .A2(n418), .ZN(n554) );
  NAND2_X1 U545 ( .A1(n546), .A2(n548), .ZN(n423) );
  XNOR2_X2 U546 ( .A(n428), .B(G122), .ZN(n489) );
  XNOR2_X2 U547 ( .A(n479), .B(n430), .ZN(n533) );
  NOR2_X1 U548 ( .A1(n658), .A2(n657), .ZN(n698) );
  INV_X1 U549 ( .A(n540), .ZN(n660) );
  BUF_X1 U550 ( .A(n528), .Z(n577) );
  XNOR2_X1 U551 ( .A(n445), .B(n444), .ZN(n446) );
  INV_X1 U552 ( .A(n731), .ZN(n629) );
  AND2_X1 U553 ( .A1(n628), .A2(G953), .ZN(n731) );
  XNOR2_X1 U554 ( .A(n496), .B(n431), .ZN(n432) );
  NAND2_X1 U555 ( .A1(n491), .A2(G210), .ZN(n434) );
  XNOR2_X1 U556 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U557 ( .A(n516), .B(n436), .ZN(n626) );
  XNOR2_X2 U558 ( .A(n437), .B(G472), .ZN(n669) );
  INV_X1 U559 ( .A(KEYINPUT6), .ZN(n438) );
  XNOR2_X1 U560 ( .A(n669), .B(n438), .ZN(n598) );
  XNOR2_X2 U561 ( .A(G146), .B(G125), .ZN(n464) );
  XNOR2_X1 U562 ( .A(KEYINPUT70), .B(KEYINPUT10), .ZN(n439) );
  NAND2_X1 U563 ( .A1(n746), .A2(G234), .ZN(n441) );
  XNOR2_X1 U564 ( .A(n441), .B(n440), .ZN(n481) );
  AND2_X1 U565 ( .A1(G221), .A2(n481), .ZN(n445) );
  XOR2_X1 U566 ( .A(KEYINPUT90), .B(KEYINPUT74), .Z(n443) );
  XNOR2_X1 U567 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U568 ( .A(KEYINPUT23), .B(KEYINPUT89), .ZN(n448) );
  INV_X1 U569 ( .A(n459), .ZN(n447) );
  XNOR2_X1 U570 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U571 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n452) );
  NAND2_X1 U572 ( .A1(G234), .A2(n619), .ZN(n451) );
  XNOR2_X1 U573 ( .A(n452), .B(n451), .ZN(n505) );
  NAND2_X1 U574 ( .A1(n505), .A2(G217), .ZN(n456) );
  XOR2_X1 U575 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n454) );
  INV_X1 U576 ( .A(n372), .ZN(n542) );
  XOR2_X1 U577 ( .A(KEYINPUT80), .B(KEYINPUT17), .Z(n463) );
  XNOR2_X1 U578 ( .A(n464), .B(n463), .ZN(n467) );
  NAND2_X1 U579 ( .A1(G224), .A2(n746), .ZN(n465) );
  XNOR2_X1 U580 ( .A(n465), .B(KEYINPUT18), .ZN(n466) );
  XNOR2_X1 U581 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U582 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U583 ( .A1(n644), .A2(n619), .ZN(n472) );
  AND2_X1 U584 ( .A1(G210), .A2(n473), .ZN(n471) );
  XNOR2_X2 U585 ( .A(n472), .B(n471), .ZN(n555) );
  NAND2_X1 U586 ( .A1(G214), .A2(n473), .ZN(n679) );
  XNOR2_X1 U587 ( .A(n474), .B(KEYINPUT14), .ZN(n475) );
  NAND2_X1 U588 ( .A1(n475), .A2(G952), .ZN(n690) );
  NOR2_X1 U589 ( .A1(G953), .A2(n690), .ZN(n562) );
  NAND2_X1 U590 ( .A1(n475), .A2(G902), .ZN(n476) );
  XNOR2_X1 U591 ( .A(n476), .B(KEYINPUT88), .ZN(n558) );
  XNOR2_X1 U592 ( .A(G898), .B(KEYINPUT87), .ZN(n737) );
  NAND2_X1 U593 ( .A1(G953), .A2(n737), .ZN(n734) );
  NOR2_X1 U594 ( .A1(n558), .A2(n734), .ZN(n477) );
  NOR2_X1 U595 ( .A1(n562), .A2(n477), .ZN(n478) );
  XOR2_X1 U596 ( .A(n480), .B(KEYINPUT7), .Z(n483) );
  NAND2_X1 U597 ( .A1(G217), .A2(n481), .ZN(n482) );
  XNOR2_X1 U598 ( .A(n483), .B(n482), .ZN(n487) );
  XNOR2_X1 U599 ( .A(n485), .B(n484), .ZN(n486) );
  NOR2_X1 U600 ( .A1(n723), .A2(G902), .ZN(n488) );
  NAND2_X1 U601 ( .A1(n491), .A2(G214), .ZN(n493) );
  XNOR2_X1 U602 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U603 ( .A(n496), .B(n495), .ZN(n500) );
  XNOR2_X1 U604 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U605 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U606 ( .A(KEYINPUT13), .B(G475), .ZN(n502) );
  XNOR2_X2 U607 ( .A(n503), .B(n502), .ZN(n581) );
  INV_X1 U608 ( .A(n581), .ZN(n504) );
  NOR2_X1 U609 ( .A1(n523), .A2(n504), .ZN(n676) );
  NAND2_X1 U610 ( .A1(G221), .A2(n505), .ZN(n506) );
  XNOR2_X1 U611 ( .A(n506), .B(KEYINPUT93), .ZN(n507) );
  XOR2_X1 U612 ( .A(KEYINPUT21), .B(n507), .Z(n663) );
  XNOR2_X1 U613 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U614 ( .A(n512), .B(n511), .Z(n514) );
  NAND2_X1 U615 ( .A1(G227), .A2(n746), .ZN(n513) );
  XNOR2_X1 U616 ( .A(n514), .B(n513), .ZN(n515) );
  INV_X1 U617 ( .A(G469), .ZN(n517) );
  INV_X1 U618 ( .A(KEYINPUT1), .ZN(n519) );
  NOR2_X1 U619 ( .A1(n541), .A2(n416), .ZN(n520) );
  NAND2_X1 U620 ( .A1(n542), .A2(n520), .ZN(n521) );
  NOR2_X1 U621 ( .A1(n598), .A2(n521), .ZN(n703) );
  OR2_X1 U622 ( .A1(n583), .A2(n522), .ZN(n704) );
  XNOR2_X1 U623 ( .A(n704), .B(KEYINPUT100), .ZN(n566) );
  INV_X1 U624 ( .A(KEYINPUT99), .ZN(n524) );
  NAND2_X1 U625 ( .A1(n566), .A2(n596), .ZN(n681) );
  XNOR2_X1 U626 ( .A(n681), .B(KEYINPUT83), .ZN(n591) );
  NOR2_X1 U627 ( .A1(n531), .A2(n574), .ZN(n525) );
  XNOR2_X1 U628 ( .A(n525), .B(KEYINPUT94), .ZN(n672) );
  INV_X1 U629 ( .A(n533), .ZN(n526) );
  NAND2_X1 U630 ( .A1(n672), .A2(n526), .ZN(n527) );
  XNOR2_X1 U631 ( .A(n527), .B(KEYINPUT31), .ZN(n720) );
  NAND2_X1 U632 ( .A1(n564), .A2(n574), .ZN(n529) );
  NOR2_X1 U633 ( .A1(n533), .A2(n529), .ZN(n705) );
  INV_X1 U634 ( .A(n598), .ZN(n530) );
  OR2_X1 U635 ( .A1(n583), .A2(n581), .ZN(n536) );
  INV_X1 U636 ( .A(KEYINPUT103), .ZN(n535) );
  XNOR2_X1 U637 ( .A(n536), .B(n535), .ZN(n605) );
  INV_X1 U638 ( .A(KEYINPUT67), .ZN(n547) );
  XNOR2_X1 U639 ( .A(n755), .B(n547), .ZN(n538) );
  INV_X1 U640 ( .A(KEYINPUT44), .ZN(n537) );
  NAND2_X1 U641 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U642 ( .A1(n539), .A2(KEYINPUT66), .ZN(n546) );
  NAND2_X1 U643 ( .A1(n660), .A2(n545), .ZN(n543) );
  NOR2_X1 U644 ( .A1(n669), .A2(n543), .ZN(n709) );
  XNOR2_X1 U645 ( .A(n598), .B(KEYINPUT81), .ZN(n544) );
  NOR2_X2 U646 ( .A1(n709), .A2(n757), .ZN(n548) );
  NAND2_X1 U647 ( .A1(n548), .A2(n547), .ZN(n550) );
  AND2_X1 U648 ( .A1(KEYINPUT44), .A2(KEYINPUT66), .ZN(n549) );
  NOR2_X1 U649 ( .A1(KEYINPUT44), .A2(KEYINPUT66), .ZN(n552) );
  NOR2_X1 U650 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U651 ( .A(n555), .B(KEYINPUT75), .ZN(n556) );
  XNOR2_X1 U652 ( .A(n556), .B(KEYINPUT38), .ZN(n680) );
  NAND2_X1 U653 ( .A1(n669), .A2(n679), .ZN(n557) );
  OR2_X1 U654 ( .A1(n746), .A2(n558), .ZN(n559) );
  NOR2_X1 U655 ( .A1(G900), .A2(n559), .ZN(n560) );
  XNOR2_X1 U656 ( .A(n560), .B(KEYINPUT104), .ZN(n561) );
  NOR2_X1 U657 ( .A1(n562), .A2(n561), .ZN(n572) );
  INV_X1 U658 ( .A(n566), .ZN(n567) );
  NAND2_X1 U659 ( .A1(n570), .A2(n567), .ZN(n568) );
  XNOR2_X1 U660 ( .A(n568), .B(KEYINPUT110), .ZN(n759) );
  NAND2_X1 U661 ( .A1(KEYINPUT2), .A2(n759), .ZN(n569) );
  XOR2_X1 U662 ( .A(KEYINPUT82), .B(n569), .Z(n618) );
  INV_X1 U663 ( .A(n596), .ZN(n714) );
  XNOR2_X2 U664 ( .A(n571), .B(KEYINPUT40), .ZN(n758) );
  INV_X1 U665 ( .A(KEYINPUT108), .ZN(n580) );
  NOR2_X1 U666 ( .A1(n572), .A2(n663), .ZN(n573) );
  NAND2_X1 U667 ( .A1(n662), .A2(n573), .ZN(n597) );
  XNOR2_X1 U668 ( .A(KEYINPUT107), .B(KEYINPUT28), .ZN(n575) );
  XNOR2_X1 U669 ( .A(n576), .B(n575), .ZN(n578) );
  NOR2_X1 U670 ( .A1(n578), .A2(n577), .ZN(n579) );
  INV_X1 U671 ( .A(n589), .ZN(n586) );
  AND2_X1 U672 ( .A1(n581), .A2(n679), .ZN(n582) );
  AND2_X1 U673 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U674 ( .A1(n680), .A2(n584), .ZN(n585) );
  NAND2_X1 U675 ( .A1(n586), .A2(n693), .ZN(n587) );
  XNOR2_X1 U676 ( .A(n587), .B(KEYINPUT42), .ZN(n760) );
  XOR2_X1 U677 ( .A(KEYINPUT68), .B(KEYINPUT47), .Z(n590) );
  NAND2_X1 U678 ( .A1(n715), .A2(n590), .ZN(n592) );
  NOR2_X1 U679 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U680 ( .A1(n715), .A2(n681), .ZN(n593) );
  AND2_X1 U681 ( .A1(n593), .A2(KEYINPUT47), .ZN(n594) );
  NAND2_X1 U682 ( .A1(n599), .A2(n598), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n610), .B(KEYINPUT109), .ZN(n602) );
  INV_X1 U684 ( .A(n600), .ZN(n601) );
  XNOR2_X1 U685 ( .A(KEYINPUT86), .B(KEYINPUT36), .ZN(n603) );
  INV_X1 U686 ( .A(n555), .ZN(n604) );
  NOR2_X1 U687 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U688 ( .A1(n607), .A2(n606), .ZN(n713) );
  INV_X1 U689 ( .A(n679), .ZN(n609) );
  NOR2_X1 U690 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U691 ( .A(n612), .B(KEYINPUT43), .Z(n613) );
  XNOR2_X1 U692 ( .A(n613), .B(KEYINPUT106), .ZN(n614) );
  INV_X1 U693 ( .A(n722), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X2 U695 ( .A(n617), .B(KEYINPUT85), .ZN(n621) );
  INV_X1 U696 ( .A(n619), .ZN(n620) );
  NAND2_X2 U697 ( .A1(n621), .A2(n759), .ZN(n745) );
  XNOR2_X1 U698 ( .A(n745), .B(KEYINPUT77), .ZN(n622) );
  INV_X1 U699 ( .A(KEYINPUT2), .ZN(n656) );
  NAND2_X1 U700 ( .A1(n649), .A2(G472), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(n361), .ZN(n630) );
  INV_X1 U702 ( .A(G952), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U704 ( .A(n631), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U705 ( .A1(n705), .A2(n714), .ZN(n632) );
  XNOR2_X1 U706 ( .A(n632), .B(G104), .ZN(G6) );
  NAND2_X1 U707 ( .A1(n720), .A2(n714), .ZN(n633) );
  XNOR2_X1 U708 ( .A(n633), .B(G113), .ZN(G15) );
  XOR2_X1 U709 ( .A(G125), .B(KEYINPUT37), .Z(n634) );
  XNOR2_X1 U710 ( .A(n635), .B(n634), .ZN(G27) );
  NAND2_X1 U711 ( .A1(n649), .A2(G475), .ZN(n639) );
  XNOR2_X1 U712 ( .A(KEYINPUT119), .B(KEYINPUT59), .ZN(n636) );
  XNOR2_X1 U713 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U714 ( .A(n639), .B(n638), .ZN(n640) );
  NOR2_X2 U715 ( .A1(n640), .A2(n731), .ZN(n642) );
  XNOR2_X1 U716 ( .A(KEYINPUT120), .B(KEYINPUT60), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n642), .B(n641), .ZN(G60) );
  NAND2_X1 U718 ( .A1(n649), .A2(G210), .ZN(n646) );
  XNOR2_X1 U719 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n643) );
  XNOR2_X1 U720 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n646), .B(n645), .ZN(n647) );
  NOR2_X2 U722 ( .A1(n647), .A2(n731), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n648), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U724 ( .A1(n727), .A2(G469), .ZN(n652) );
  XNOR2_X1 U725 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n650) );
  XNOR2_X1 U726 ( .A(n652), .B(n651), .ZN(n653) );
  AND2_X1 U727 ( .A1(n653), .A2(n629), .ZN(G54) );
  NAND2_X1 U728 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U730 ( .A(KEYINPUT50), .B(n661), .ZN(n667) );
  XOR2_X1 U731 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n665) );
  NAND2_X1 U732 ( .A1(n663), .A2(n372), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U736 ( .A(KEYINPUT115), .B(n670), .Z(n671) );
  NOR2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U738 ( .A(KEYINPUT51), .B(n673), .ZN(n674) );
  NAND2_X1 U739 ( .A1(n674), .A2(n693), .ZN(n675) );
  XOR2_X1 U740 ( .A(KEYINPUT116), .B(n675), .Z(n688) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n678) );
  INV_X1 U742 ( .A(n676), .ZN(n677) );
  NOR2_X1 U743 ( .A1(n678), .A2(n677), .ZN(n685) );
  NAND2_X1 U744 ( .A1(n680), .A2(n679), .ZN(n683) );
  INV_X1 U745 ( .A(n681), .ZN(n682) );
  NOR2_X1 U746 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U747 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U748 ( .A1(n686), .A2(n692), .ZN(n687) );
  NOR2_X1 U749 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U750 ( .A(n689), .B(KEYINPUT52), .ZN(n691) );
  OR2_X1 U751 ( .A1(n691), .A2(n690), .ZN(n696) );
  INV_X1 U752 ( .A(n692), .ZN(n694) );
  NAND2_X1 U753 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U754 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U755 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U756 ( .A(n699), .B(KEYINPUT117), .ZN(n700) );
  XNOR2_X1 U757 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n701) );
  XNOR2_X1 U758 ( .A(n702), .B(n701), .ZN(G75) );
  XOR2_X1 U759 ( .A(G101), .B(n703), .Z(G3) );
  XOR2_X1 U760 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n707) );
  INV_X1 U761 ( .A(n704), .ZN(n719) );
  NAND2_X1 U762 ( .A1(n705), .A2(n719), .ZN(n706) );
  XNOR2_X1 U763 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U764 ( .A(G107), .B(n708), .ZN(G9) );
  XNOR2_X1 U765 ( .A(G110), .B(n709), .ZN(n710) );
  XNOR2_X1 U766 ( .A(n710), .B(KEYINPUT111), .ZN(G12) );
  XOR2_X1 U767 ( .A(G128), .B(KEYINPUT29), .Z(n712) );
  NAND2_X1 U768 ( .A1(n715), .A2(n719), .ZN(n711) );
  XNOR2_X1 U769 ( .A(n712), .B(n711), .ZN(G30) );
  XNOR2_X1 U770 ( .A(G143), .B(n713), .ZN(G45) );
  NAND2_X1 U771 ( .A1(n715), .A2(n714), .ZN(n717) );
  XOR2_X1 U772 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n716) );
  XNOR2_X1 U773 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U774 ( .A(G146), .B(n718), .ZN(G48) );
  NAND2_X1 U775 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U776 ( .A(n721), .B(G116), .ZN(G18) );
  XOR2_X1 U777 ( .A(G140), .B(n722), .Z(G42) );
  NAND2_X1 U778 ( .A1(n727), .A2(G478), .ZN(n725) );
  XOR2_X1 U779 ( .A(n723), .B(KEYINPUT121), .Z(n724) );
  XNOR2_X1 U780 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U781 ( .A1(n731), .A2(n726), .ZN(G63) );
  NAND2_X1 U782 ( .A1(n727), .A2(G217), .ZN(n729) );
  XNOR2_X1 U783 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U784 ( .A1(n731), .A2(n730), .ZN(G66) );
  XOR2_X1 U785 ( .A(n732), .B(KEYINPUT123), .Z(n733) );
  NAND2_X1 U786 ( .A1(n734), .A2(n733), .ZN(n742) );
  XOR2_X1 U787 ( .A(KEYINPUT61), .B(KEYINPUT122), .Z(n736) );
  NAND2_X1 U788 ( .A1(G224), .A2(G953), .ZN(n735) );
  XNOR2_X1 U789 ( .A(n736), .B(n735), .ZN(n738) );
  NOR2_X1 U790 ( .A1(n738), .A2(n737), .ZN(n740) );
  NOR2_X1 U791 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U792 ( .A(n742), .B(n741), .ZN(G69) );
  XNOR2_X1 U793 ( .A(n744), .B(n743), .ZN(n748) );
  XNOR2_X1 U794 ( .A(n745), .B(n748), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n747), .A2(n746), .ZN(n753) );
  XNOR2_X1 U796 ( .A(n748), .B(G227), .ZN(n749) );
  XNOR2_X1 U797 ( .A(n749), .B(KEYINPUT124), .ZN(n750) );
  NAND2_X1 U798 ( .A1(n750), .A2(G900), .ZN(n751) );
  NAND2_X1 U799 ( .A1(G953), .A2(n751), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U801 ( .A(KEYINPUT125), .B(n754), .Z(G72) );
  XNOR2_X1 U802 ( .A(n755), .B(G122), .ZN(G24) );
  XOR2_X1 U803 ( .A(G119), .B(KEYINPUT126), .Z(n756) );
  XNOR2_X1 U804 ( .A(n757), .B(n756), .ZN(G21) );
  XNOR2_X1 U805 ( .A(n758), .B(G131), .ZN(G33) );
  XNOR2_X1 U806 ( .A(G134), .B(n759), .ZN(G36) );
  XOR2_X1 U807 ( .A(n760), .B(G137), .Z(n761) );
  XNOR2_X1 U808 ( .A(KEYINPUT127), .B(n761), .ZN(G39) );
endmodule

