

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591;

  XNOR2_X1 U325 ( .A(n388), .B(n387), .ZN(n573) );
  XNOR2_X1 U326 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n387) );
  XNOR2_X1 U327 ( .A(n334), .B(n306), .ZN(n307) );
  XNOR2_X1 U328 ( .A(n308), .B(n307), .ZN(n310) );
  XNOR2_X1 U329 ( .A(n364), .B(KEYINPUT41), .ZN(n551) );
  XNOR2_X1 U330 ( .A(n452), .B(G190GAT), .ZN(n453) );
  XNOR2_X1 U331 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XNOR2_X1 U332 ( .A(KEYINPUT32), .B(KEYINPUT69), .ZN(n294) );
  AND2_X1 U333 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U335 ( .A(n295), .B(KEYINPUT68), .ZN(n304) );
  INV_X1 U336 ( .A(G92GAT), .ZN(n296) );
  NAND2_X1 U337 ( .A1(n296), .A2(G64GAT), .ZN(n299) );
  INV_X1 U338 ( .A(G64GAT), .ZN(n297) );
  NAND2_X1 U339 ( .A1(n297), .A2(G92GAT), .ZN(n298) );
  NAND2_X1 U340 ( .A1(n299), .A2(n298), .ZN(n301) );
  XNOR2_X1 U341 ( .A(G176GAT), .B(G204GAT), .ZN(n300) );
  XNOR2_X1 U342 ( .A(n301), .B(n300), .ZN(n379) );
  XNOR2_X1 U343 ( .A(G106GAT), .B(G78GAT), .ZN(n302) );
  XNOR2_X1 U344 ( .A(n302), .B(G148GAT), .ZN(n402) );
  XNOR2_X1 U345 ( .A(n379), .B(n402), .ZN(n303) );
  XNOR2_X1 U346 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U347 ( .A(G120GAT), .B(G57GAT), .Z(n419) );
  XNOR2_X1 U348 ( .A(n305), .B(n419), .ZN(n308) );
  XOR2_X1 U349 ( .A(G99GAT), .B(G85GAT), .Z(n334) );
  XNOR2_X1 U350 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n306) );
  XOR2_X1 U351 ( .A(G71GAT), .B(KEYINPUT13), .Z(n352) );
  INV_X1 U352 ( .A(n352), .ZN(n309) );
  XOR2_X1 U353 ( .A(n310), .B(n309), .Z(n580) );
  INV_X1 U354 ( .A(n580), .ZN(n364) );
  XOR2_X1 U355 ( .A(G29GAT), .B(G43GAT), .Z(n312) );
  XNOR2_X1 U356 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n311) );
  XNOR2_X1 U357 ( .A(n312), .B(n311), .ZN(n329) );
  XOR2_X1 U358 ( .A(n329), .B(KEYINPUT29), .Z(n314) );
  NAND2_X1 U359 ( .A1(G229GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U360 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U361 ( .A(G169GAT), .B(G8GAT), .Z(n382) );
  XOR2_X1 U362 ( .A(n315), .B(n382), .Z(n317) );
  XNOR2_X1 U363 ( .A(G50GAT), .B(G36GAT), .ZN(n316) );
  XNOR2_X1 U364 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U365 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n319) );
  XNOR2_X1 U366 ( .A(G197GAT), .B(G15GAT), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U368 ( .A(n321), .B(n320), .Z(n323) );
  XOR2_X1 U369 ( .A(G141GAT), .B(G22GAT), .Z(n394) );
  XOR2_X1 U370 ( .A(G113GAT), .B(G1GAT), .Z(n420) );
  XNOR2_X1 U371 ( .A(n394), .B(n420), .ZN(n322) );
  XNOR2_X1 U372 ( .A(n323), .B(n322), .ZN(n576) );
  NAND2_X1 U373 ( .A1(n551), .A2(n576), .ZN(n325) );
  XOR2_X1 U374 ( .A(KEYINPUT46), .B(KEYINPUT107), .Z(n324) );
  XNOR2_X1 U375 ( .A(n325), .B(n324), .ZN(n361) );
  XOR2_X1 U376 ( .A(G134GAT), .B(KEYINPUT70), .Z(n414) );
  XOR2_X1 U377 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n327) );
  XNOR2_X1 U378 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U380 ( .A(n414), .B(n328), .Z(n331) );
  XOR2_X1 U381 ( .A(G50GAT), .B(G162GAT), .Z(n390) );
  XNOR2_X1 U382 ( .A(n329), .B(n390), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n339) );
  XOR2_X1 U384 ( .A(KEYINPUT66), .B(G92GAT), .Z(n333) );
  NAND2_X1 U385 ( .A1(G232GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U386 ( .A(n333), .B(n332), .ZN(n335) );
  XOR2_X1 U387 ( .A(n335), .B(n334), .Z(n337) );
  XOR2_X1 U388 ( .A(G36GAT), .B(G190GAT), .Z(n378) );
  XNOR2_X1 U389 ( .A(G106GAT), .B(n378), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U391 ( .A(n339), .B(n338), .Z(n557) );
  XOR2_X1 U392 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n341) );
  XNOR2_X1 U393 ( .A(KEYINPUT12), .B(KEYINPUT72), .ZN(n340) );
  XNOR2_X1 U394 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U395 ( .A(G57GAT), .B(G64GAT), .Z(n343) );
  XNOR2_X1 U396 ( .A(KEYINPUT73), .B(KEYINPUT71), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n359) );
  XOR2_X1 U399 ( .A(G155GAT), .B(G211GAT), .Z(n347) );
  XNOR2_X1 U400 ( .A(G22GAT), .B(G78GAT), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U402 ( .A(KEYINPUT15), .B(G183GAT), .Z(n349) );
  XNOR2_X1 U403 ( .A(G15GAT), .B(G127GAT), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U405 ( .A(n351), .B(n350), .Z(n357) );
  XOR2_X1 U406 ( .A(G8GAT), .B(n352), .Z(n354) );
  NAND2_X1 U407 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U409 ( .A(G1GAT), .B(n355), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n359), .B(n358), .ZN(n583) );
  NOR2_X1 U412 ( .A1(n557), .A2(n583), .ZN(n360) );
  NAND2_X1 U413 ( .A1(n361), .A2(n360), .ZN(n363) );
  XOR2_X1 U414 ( .A(KEYINPUT47), .B(KEYINPUT108), .Z(n362) );
  XNOR2_X1 U415 ( .A(n363), .B(n362), .ZN(n371) );
  XOR2_X1 U416 ( .A(KEYINPUT45), .B(KEYINPUT109), .Z(n367) );
  XNOR2_X1 U417 ( .A(n557), .B(KEYINPUT96), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n365), .B(KEYINPUT36), .ZN(n586) );
  NAND2_X1 U419 ( .A1(n583), .A2(n586), .ZN(n366) );
  XNOR2_X1 U420 ( .A(n367), .B(n366), .ZN(n368) );
  NOR2_X1 U421 ( .A1(n368), .A2(n576), .ZN(n369) );
  NAND2_X1 U422 ( .A1(n364), .A2(n369), .ZN(n370) );
  AND2_X1 U423 ( .A1(n371), .A2(n370), .ZN(n373) );
  XOR2_X1 U424 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n372) );
  XNOR2_X1 U425 ( .A(n373), .B(n372), .ZN(n545) );
  XOR2_X1 U426 ( .A(G211GAT), .B(KEYINPUT21), .Z(n375) );
  XNOR2_X1 U427 ( .A(G197GAT), .B(G218GAT), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n401) );
  XOR2_X1 U429 ( .A(KEYINPUT86), .B(n401), .Z(n377) );
  NAND2_X1 U430 ( .A1(G226GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U431 ( .A(n377), .B(n376), .ZN(n386) );
  XOR2_X1 U432 ( .A(n379), .B(n378), .Z(n384) );
  XOR2_X1 U433 ( .A(G183GAT), .B(KEYINPUT18), .Z(n381) );
  XNOR2_X1 U434 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n380) );
  XNOR2_X1 U435 ( .A(n381), .B(n380), .ZN(n446) );
  XNOR2_X1 U436 ( .A(n382), .B(n446), .ZN(n383) );
  XNOR2_X1 U437 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U438 ( .A(n386), .B(n385), .Z(n518) );
  NAND2_X1 U439 ( .A1(n545), .A2(n518), .ZN(n388) );
  XNOR2_X1 U440 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n389) );
  XNOR2_X1 U441 ( .A(n389), .B(KEYINPUT2), .ZN(n424) );
  XOR2_X1 U442 ( .A(n424), .B(n390), .Z(n392) );
  NAND2_X1 U443 ( .A1(G228GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U444 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U445 ( .A(n393), .B(KEYINPUT24), .Z(n396) );
  XNOR2_X1 U446 ( .A(n394), .B(KEYINPUT79), .ZN(n395) );
  XNOR2_X1 U447 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U448 ( .A(G204GAT), .B(KEYINPUT80), .Z(n398) );
  XNOR2_X1 U449 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U451 ( .A(n400), .B(n399), .Z(n404) );
  XNOR2_X1 U452 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U453 ( .A(n404), .B(n403), .ZN(n463) );
  XOR2_X1 U454 ( .A(KEYINPUT85), .B(KEYINPUT83), .Z(n406) );
  XNOR2_X1 U455 ( .A(KEYINPUT6), .B(KEYINPUT81), .ZN(n405) );
  XNOR2_X1 U456 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U457 ( .A(KEYINPUT82), .B(KEYINPUT4), .Z(n408) );
  XNOR2_X1 U458 ( .A(G141GAT), .B(KEYINPUT1), .ZN(n407) );
  XNOR2_X1 U459 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U460 ( .A(n410), .B(n409), .ZN(n428) );
  XOR2_X1 U461 ( .A(G85GAT), .B(G162GAT), .Z(n412) );
  XNOR2_X1 U462 ( .A(G29GAT), .B(G148GAT), .ZN(n411) );
  XNOR2_X1 U463 ( .A(n412), .B(n411), .ZN(n418) );
  XNOR2_X1 U464 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n413) );
  XNOR2_X1 U465 ( .A(n413), .B(KEYINPUT75), .ZN(n447) );
  XOR2_X1 U466 ( .A(n414), .B(n447), .Z(n416) );
  NAND2_X1 U467 ( .A1(G225GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U468 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U469 ( .A(n418), .B(n417), .Z(n422) );
  XNOR2_X1 U470 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U471 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U472 ( .A(n423), .B(KEYINPUT5), .Z(n426) );
  XNOR2_X1 U473 ( .A(n424), .B(KEYINPUT84), .ZN(n425) );
  XNOR2_X1 U474 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U475 ( .A(n428), .B(n427), .ZN(n572) );
  INV_X1 U476 ( .A(n572), .ZN(n516) );
  NOR2_X1 U477 ( .A1(n463), .A2(n516), .ZN(n429) );
  AND2_X1 U478 ( .A1(n573), .A2(n429), .ZN(n430) );
  XNOR2_X1 U479 ( .A(n430), .B(KEYINPUT55), .ZN(n450) );
  XOR2_X1 U480 ( .A(G99GAT), .B(G190GAT), .Z(n432) );
  XNOR2_X1 U481 ( .A(G43GAT), .B(G134GAT), .ZN(n431) );
  XNOR2_X1 U482 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U483 ( .A(KEYINPUT76), .B(KEYINPUT20), .Z(n434) );
  XNOR2_X1 U484 ( .A(G120GAT), .B(KEYINPUT65), .ZN(n433) );
  XNOR2_X1 U485 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U486 ( .A(n436), .B(n435), .Z(n441) );
  XOR2_X1 U487 ( .A(KEYINPUT78), .B(G71GAT), .Z(n438) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U490 ( .A(G113GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U491 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U492 ( .A(G176GAT), .B(KEYINPUT77), .Z(n443) );
  XNOR2_X1 U493 ( .A(G169GAT), .B(G15GAT), .ZN(n442) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U495 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U496 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U497 ( .A(n449), .B(n448), .ZN(n497) );
  NOR2_X1 U498 ( .A1(n450), .A2(n497), .ZN(n451) );
  XOR2_X1 U499 ( .A(KEYINPUT120), .B(n451), .Z(n568) );
  INV_X1 U500 ( .A(n557), .ZN(n539) );
  NOR2_X1 U501 ( .A1(n568), .A2(n539), .ZN(n454) );
  INV_X1 U502 ( .A(KEYINPUT58), .ZN(n452) );
  XOR2_X1 U503 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n456) );
  XNOR2_X1 U504 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n455) );
  XNOR2_X1 U505 ( .A(n456), .B(n455), .ZN(n472) );
  INV_X1 U506 ( .A(n576), .ZN(n560) );
  NOR2_X1 U507 ( .A1(n580), .A2(n560), .ZN(n487) );
  INV_X1 U508 ( .A(n497), .ZN(n526) );
  XOR2_X1 U509 ( .A(n463), .B(KEYINPUT28), .Z(n508) );
  XOR2_X1 U510 ( .A(n518), .B(KEYINPUT27), .Z(n461) );
  NOR2_X1 U511 ( .A1(n572), .A2(n461), .ZN(n457) );
  NAND2_X1 U512 ( .A1(n508), .A2(n457), .ZN(n528) );
  NOR2_X1 U513 ( .A1(n526), .A2(n528), .ZN(n468) );
  XOR2_X1 U514 ( .A(KEYINPUT88), .B(KEYINPUT26), .Z(n459) );
  NAND2_X1 U515 ( .A1(n463), .A2(n497), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U517 ( .A(KEYINPUT87), .B(n460), .ZN(n574) );
  NOR2_X1 U518 ( .A1(n461), .A2(n574), .ZN(n546) );
  INV_X1 U519 ( .A(n518), .ZN(n492) );
  NOR2_X1 U520 ( .A1(n497), .A2(n492), .ZN(n462) );
  NOR2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n464) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n464), .Z(n465) );
  NOR2_X1 U523 ( .A1(n546), .A2(n465), .ZN(n466) );
  NOR2_X1 U524 ( .A1(n466), .A2(n516), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n468), .A2(n467), .ZN(n483) );
  INV_X1 U526 ( .A(n583), .ZN(n567) );
  NOR2_X1 U527 ( .A1(n557), .A2(n567), .ZN(n469) );
  XOR2_X1 U528 ( .A(KEYINPUT16), .B(n469), .Z(n470) );
  NOR2_X1 U529 ( .A1(n483), .A2(n470), .ZN(n502) );
  NAND2_X1 U530 ( .A1(n487), .A2(n502), .ZN(n480) );
  NOR2_X1 U531 ( .A1(n572), .A2(n480), .ZN(n471) );
  XOR2_X1 U532 ( .A(n472), .B(n471), .Z(G1324GAT) );
  NOR2_X1 U533 ( .A1(n492), .A2(n480), .ZN(n474) );
  XNOR2_X1 U534 ( .A(G8GAT), .B(KEYINPUT91), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n474), .B(n473), .ZN(G1325GAT) );
  NOR2_X1 U536 ( .A1(n497), .A2(n480), .ZN(n479) );
  XOR2_X1 U537 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n476) );
  XNOR2_X1 U538 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n475) );
  XNOR2_X1 U539 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U540 ( .A(KEYINPUT92), .B(n477), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  NOR2_X1 U542 ( .A1(n508), .A2(n480), .ZN(n482) );
  XNOR2_X1 U543 ( .A(G22GAT), .B(KEYINPUT95), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n482), .B(n481), .ZN(G1327GAT) );
  XNOR2_X1 U545 ( .A(KEYINPUT98), .B(KEYINPUT39), .ZN(n490) );
  NOR2_X1 U546 ( .A1(n583), .A2(n483), .ZN(n484) );
  NAND2_X1 U547 ( .A1(n586), .A2(n484), .ZN(n485) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n485), .ZN(n486) );
  XOR2_X1 U549 ( .A(KEYINPUT97), .B(n486), .Z(n513) );
  NAND2_X1 U550 ( .A1(n487), .A2(n513), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n488), .B(KEYINPUT38), .ZN(n500) );
  NOR2_X1 U552 ( .A1(n572), .A2(n500), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(n491), .ZN(G1328GAT) );
  NOR2_X1 U555 ( .A1(n500), .A2(n492), .ZN(n494) );
  XNOR2_X1 U556 ( .A(G36GAT), .B(KEYINPUT99), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(G1329GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n496) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(n499) );
  NOR2_X1 U561 ( .A1(n497), .A2(n500), .ZN(n498) );
  XOR2_X1 U562 ( .A(n499), .B(n498), .Z(G1330GAT) );
  NOR2_X1 U563 ( .A1(n508), .A2(n500), .ZN(n501) );
  XOR2_X1 U564 ( .A(G50GAT), .B(n501), .Z(G1331GAT) );
  XOR2_X1 U565 ( .A(n551), .B(KEYINPUT102), .Z(n563) );
  NOR2_X1 U566 ( .A1(n576), .A2(n563), .ZN(n514) );
  NAND2_X1 U567 ( .A1(n514), .A2(n502), .ZN(n503) );
  XNOR2_X1 U568 ( .A(KEYINPUT103), .B(n503), .ZN(n509) );
  NAND2_X1 U569 ( .A1(n516), .A2(n509), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(KEYINPUT42), .ZN(n505) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U572 ( .A1(n509), .A2(n518), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n506), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n526), .A2(n509), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n511) );
  INV_X1 U577 ( .A(n508), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n509), .A2(n521), .ZN(n510) );
  XNOR2_X1 U579 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  NAND2_X1 U581 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(KEYINPUT105), .ZN(n522) );
  NAND2_X1 U583 ( .A1(n522), .A2(n516), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n522), .A2(n518), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n526), .A2(n522), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n520), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT106), .B(KEYINPUT44), .Z(n524) );
  NAND2_X1 U590 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U592 ( .A(G106GAT), .B(n525), .Z(G1339GAT) );
  NAND2_X1 U593 ( .A1(n526), .A2(n545), .ZN(n527) );
  NOR2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n534), .A2(n576), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n529), .B(KEYINPUT110), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  INV_X1 U598 ( .A(n534), .ZN(n540) );
  NOR2_X1 U599 ( .A1(n563), .A2(n540), .ZN(n532) );
  XNOR2_X1 U600 ( .A(KEYINPUT111), .B(KEYINPUT49), .ZN(n531) );
  XNOR2_X1 U601 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U602 ( .A(G120GAT), .B(n533), .Z(G1341GAT) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(KEYINPUT113), .ZN(n538) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT112), .Z(n536) );
  NAND2_X1 U605 ( .A1(n534), .A2(n583), .ZN(n535) );
  XNOR2_X1 U606 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U607 ( .A(n538), .B(n537), .ZN(G1342GAT) );
  NOR2_X1 U608 ( .A1(n540), .A2(n539), .ZN(n544) );
  XOR2_X1 U609 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n542) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT114), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  XOR2_X1 U613 ( .A(G141GAT), .B(KEYINPUT117), .Z(n550) );
  NAND2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U615 ( .A1(n547), .A2(n572), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(KEYINPUT116), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n576), .A2(n558), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(G1344GAT) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n555) );
  XOR2_X1 U620 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n553) );
  NAND2_X1 U621 ( .A1(n551), .A2(n558), .ZN(n552) );
  XNOR2_X1 U622 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n583), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U628 ( .A1(n568), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(G1348GAT) );
  XNOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n565) );
  NOR2_X1 U632 ( .A1(n568), .A2(n563), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n566), .B(G176GAT), .ZN(G1349GAT) );
  NOR2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U636 ( .A(G183GAT), .B(n569), .Z(G1350GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n571) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n571), .B(n570), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n575) );
  NOR2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n587) );
  NAND2_X1 U642 ( .A1(n587), .A2(n576), .ZN(n577) );
  XOR2_X1 U643 ( .A(n578), .B(n577), .Z(n579) );
  XNOR2_X1 U644 ( .A(KEYINPUT59), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  NAND2_X1 U646 ( .A1(n587), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n587), .A2(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(KEYINPUT124), .ZN(n585) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(n585), .ZN(G1354GAT) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n591) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n589) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(G1355GAT) );
endmodule

