//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n465), .C1(new_n459), .C2(new_n460), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n470), .B1(new_n468), .B2(new_n469), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n464), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  OR2_X1    g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n465), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n465), .B1(new_n475), .B2(new_n476), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n488), .B(new_n489), .C1(new_n460), .C2(new_n459), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT67), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(new_n465), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n481), .A2(G126), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n465), .A2(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n475), .B2(new_n476), .ZN(new_n499));
  AOI21_X1  g074(.A(KEYINPUT67), .B1(new_n499), .B2(new_n489), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n488), .B(KEYINPUT67), .C1(new_n460), .C2(new_n459), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n493), .B(new_n497), .C1(new_n500), .C2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n505), .A2(new_n509), .A3(G88), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI211_X1 g087(.A(G50), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT69), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n510), .A2(new_n516), .A3(new_n513), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n508), .B1(new_n515), .B2(new_n517), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT70), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT7), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n524), .A2(new_n525), .B1(new_n511), .B2(new_n512), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n509), .A2(G543), .ZN(new_n529));
  OAI221_X1 g104(.A(new_n523), .B1(new_n526), .B2(new_n527), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  OR3_X1    g105(.A1(new_n522), .A2(new_n530), .A3(KEYINPUT71), .ZN(new_n531));
  OAI21_X1  g106(.A(KEYINPUT71), .B1(new_n522), .B2(new_n530), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(G168));
  NAND2_X1  g108(.A1(new_n505), .A2(G64), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n507), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  INV_X1    g114(.A(new_n526), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n511), .A2(new_n512), .ZN(new_n541));
  INV_X1    g116(.A(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n540), .A2(G90), .B1(new_n543), .B2(G52), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n538), .A2(new_n539), .A3(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n525), .A2(new_n524), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G651), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI221_X1 g128(.A(new_n551), .B1(new_n552), .B2(new_n529), .C1(new_n553), .C2(new_n526), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT73), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n505), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n505), .A2(new_n563), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  XOR2_X1   g143(.A(new_n568), .B(KEYINPUT75), .Z(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(KEYINPUT74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n543), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n543), .A2(new_n576), .A3(new_n573), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n575), .A2(new_n577), .B1(G91), .B2(new_n540), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n571), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G168), .ZN(G286));
  INV_X1    g155(.A(new_n517), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n516), .B1(new_n510), .B2(new_n513), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n581), .A2(new_n582), .B1(new_n507), .B2(new_n506), .ZN(G303));
  NAND2_X1  g158(.A1(new_n540), .A2(G87), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n543), .A2(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  INV_X1    g162(.A(G48), .ZN(new_n588));
  INV_X1    g163(.A(G86), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n529), .A2(new_n588), .B1(new_n526), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n505), .A2(G61), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n507), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n507), .ZN(new_n597));
  INV_X1    g172(.A(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n529), .A2(new_n598), .B1(new_n526), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(new_n565), .B2(new_n566), .ZN(new_n605));
  AND2_X1   g180(.A1(G79), .A2(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(G651), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n526), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n540), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n529), .A2(KEYINPUT77), .ZN(new_n612));
  INV_X1    g187(.A(G54), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n529), .B2(KEYINPUT77), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n610), .A2(new_n611), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n603), .B1(new_n617), .B2(G868), .ZN(G284));
  XNOR2_X1  g193(.A(G284), .B(KEYINPUT78), .ZN(G321));
  NOR2_X1   g194(.A1(G299), .A2(G868), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g196(.A(new_n620), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(G148));
  NOR2_X1   g199(.A1(new_n554), .A2(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n617), .A2(new_n623), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT79), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n625), .B1(new_n627), .B2(G868), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g204(.A1(new_n461), .A2(new_n466), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT13), .B(G2100), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n481), .A2(G123), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n465), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(G135), .ZN(new_n637));
  OAI221_X1 g212(.A(new_n634), .B1(new_n635), .B2(new_n636), .C1(new_n637), .C2(new_n478), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(KEYINPUT80), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(KEYINPUT80), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  AND2_X1   g217(.A1(new_n642), .A2(G2096), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(G2096), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n633), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT81), .Z(G156));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT82), .ZN(new_n660));
  INV_X1    g235(.A(G14), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n657), .B2(new_n658), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT83), .Z(G401));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT17), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT85), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n665), .A3(new_n667), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT84), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT18), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n666), .A2(new_n667), .ZN(new_n676));
  INV_X1    g251(.A(new_n665), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n669), .B1(new_n677), .B2(new_n668), .ZN(new_n678));
  AOI211_X1 g253(.A(new_n672), .B(new_n675), .C1(new_n676), .C2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G227));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT86), .ZN(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  NAND3_X1  g266(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT20), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n693), .B(new_n696), .C1(new_n687), .C2(new_n695), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1991), .B(G1996), .Z(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n699), .A2(new_n701), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n685), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n704), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n706), .A2(new_n684), .A3(new_n702), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(G229));
  NOR2_X1   g284(.A1(G6), .A2(G16), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n594), .B2(G16), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT88), .Z(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT32), .B(G1981), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G1971), .ZN(new_n716));
  NAND2_X1  g291(.A1(G166), .A2(G16), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G16), .B2(G22), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n712), .A2(new_n714), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G23), .ZN(new_n721));
  AND3_X1   g296(.A1(new_n584), .A2(new_n586), .A3(new_n585), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n720), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT33), .B(G1976), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n718), .A2(new_n716), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n715), .A2(new_n719), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G25), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n479), .A2(G131), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n481), .A2(G119), .ZN(new_n733));
  OR2_X1    g308(.A1(G95), .A2(G2105), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n734), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n731), .B1(new_n737), .B2(new_n730), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT35), .B(G1991), .Z(new_n739));
  XOR2_X1   g314(.A(new_n738), .B(new_n739), .Z(new_n740));
  INV_X1    g315(.A(G24), .ZN(new_n741));
  OR3_X1    g316(.A1(new_n741), .A2(KEYINPUT87), .A3(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(KEYINPUT87), .B1(new_n741), .B2(G16), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n742), .B(new_n743), .C1(new_n601), .C2(new_n720), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1986), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n728), .A2(new_n729), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(KEYINPUT36), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n728), .A2(new_n749), .A3(new_n729), .A4(new_n746), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n720), .A2(G21), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G168), .B2(new_n720), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n753), .A2(G1966), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n720), .A2(G20), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT23), .Z(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G299), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1956), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n753), .A2(G1966), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n754), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n730), .A2(G26), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT28), .ZN(new_n763));
  OAI21_X1  g338(.A(KEYINPUT91), .B1(G104), .B2(G2105), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NOR3_X1   g340(.A1(KEYINPUT91), .A2(G104), .A3(G2105), .ZN(new_n766));
  OAI221_X1 g341(.A(G2104), .B1(G116), .B2(new_n465), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT92), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n479), .A2(G140), .B1(G128), .B2(new_n481), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n763), .B1(new_n771), .B2(new_n730), .ZN(new_n772));
  INV_X1    g347(.A(G2067), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G1961), .ZN(new_n775));
  NOR2_X1   g350(.A1(G171), .A2(new_n720), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G5), .B2(new_n720), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n774), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G16), .A2(G19), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n555), .B2(G16), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(G1341), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(G1341), .ZN(new_n782));
  INV_X1    g357(.A(G28), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(KEYINPUT30), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n730), .B1(new_n785), .B2(G28), .ZN(new_n786));
  NOR2_X1   g361(.A1(KEYINPUT31), .A2(G11), .ZN(new_n787));
  AND2_X1   g362(.A1(KEYINPUT31), .A2(G11), .ZN(new_n788));
  OAI221_X1 g363(.A(new_n782), .B1(new_n784), .B2(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n730), .A2(G35), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G162), .B2(new_n730), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT29), .B(G2090), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n641), .A2(new_n730), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n778), .A2(new_n781), .A3(new_n789), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G29), .A2(G33), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT93), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n479), .A2(G139), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT94), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(new_n465), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT25), .Z(new_n805));
  NAND3_X1  g380(.A1(new_n801), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n799), .B1(new_n806), .B2(new_n730), .ZN(new_n807));
  INV_X1    g382(.A(G2072), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n730), .A2(G32), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n479), .A2(G141), .B1(G105), .B2(new_n467), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n481), .A2(G129), .ZN(new_n812));
  NAND3_X1  g387(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT26), .Z(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n810), .B1(new_n816), .B2(new_n730), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT27), .B(G1996), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n795), .A2(new_n794), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n807), .A2(new_n808), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n809), .A2(new_n819), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n730), .A2(G27), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT97), .Z(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n503), .B2(G29), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT98), .B(G2078), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n777), .A2(new_n775), .ZN(new_n829));
  INV_X1    g404(.A(G2084), .ZN(new_n830));
  INV_X1    g405(.A(G34), .ZN(new_n831));
  AOI21_X1  g406(.A(G29), .B1(new_n831), .B2(KEYINPUT24), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(KEYINPUT24), .B2(new_n831), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n473), .B2(new_n730), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n829), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n830), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT96), .Z(new_n837));
  NOR2_X1   g412(.A1(G4), .A2(G16), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT89), .Z(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n616), .B2(new_n720), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT90), .B(G1348), .Z(new_n841));
  XOR2_X1   g416(.A(new_n840), .B(new_n841), .Z(new_n842));
  NOR3_X1   g417(.A1(new_n835), .A2(new_n837), .A3(new_n842), .ZN(new_n843));
  AND4_X1   g418(.A1(new_n761), .A2(new_n797), .A3(new_n828), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n751), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT99), .ZN(G311));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(G150));
  NOR2_X1   g423(.A1(new_n616), .A2(new_n623), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(new_n507), .ZN(new_n853));
  INV_X1    g428(.A(G55), .ZN(new_n854));
  INV_X1    g429(.A(G93), .ZN(new_n855));
  OAI22_X1  g430(.A1(new_n529), .A2(new_n854), .B1(new_n526), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n554), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n851), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n860));
  AOI21_X1  g435(.A(G860), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n860), .B2(new_n859), .ZN(new_n862));
  OAI21_X1  g437(.A(G860), .B1(new_n853), .B2(new_n856), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT37), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(G145));
  NOR2_X1   g440(.A1(new_n770), .A2(new_n503), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n770), .A2(new_n503), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n867), .A2(new_n806), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n806), .B1(new_n867), .B2(new_n868), .ZN(new_n870));
  OR3_X1    g445(.A1(new_n869), .A2(new_n870), .A3(new_n815), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n815), .B1(new_n869), .B2(new_n870), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n481), .A2(G130), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n465), .A2(G118), .ZN(new_n876));
  OAI21_X1  g451(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n877));
  INV_X1    g452(.A(G142), .ZN(new_n878));
  OAI221_X1 g453(.A(new_n875), .B1(new_n876), .B2(new_n877), .C1(new_n878), .C2(new_n478), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n631), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n736), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n880), .A2(new_n736), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n874), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(KEYINPUT102), .A3(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n873), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n887), .B1(new_n871), .B2(new_n872), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT103), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n871), .A2(new_n887), .A3(new_n872), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n485), .B(new_n473), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n641), .ZN(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n892), .A2(new_n897), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n871), .A2(new_n872), .A3(new_n885), .A4(new_n881), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(KEYINPUT104), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n898), .A2(new_n905), .A3(KEYINPUT40), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT40), .B1(new_n898), .B2(new_n905), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(G395));
  INV_X1    g483(.A(new_n858), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n627), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n627), .A2(new_n909), .ZN(new_n911));
  AND2_X1   g486(.A1(G299), .A2(new_n616), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n571), .A2(new_n607), .A3(new_n578), .A4(new_n615), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n910), .B(new_n911), .C1(new_n912), .C2(new_n914), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n910), .A2(new_n911), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT41), .B1(new_n912), .B2(new_n914), .ZN(new_n917));
  NAND2_X1  g492(.A1(G299), .A2(new_n616), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n913), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n915), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(G303), .B(KEYINPUT105), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(G305), .ZN(new_n926));
  XNOR2_X1  g501(.A(G166), .B(KEYINPUT105), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n594), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G290), .A2(G288), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n722), .A2(new_n601), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT106), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n931), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n932), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n928), .B2(new_n926), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n915), .B(KEYINPUT42), .C1(new_n916), .C2(new_n921), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n924), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n924), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g517(.A(G868), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n857), .A2(G868), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(G295));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n944), .ZN(G331));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n531), .A2(new_n532), .A3(G301), .ZN(new_n948));
  AOI21_X1  g523(.A(G301), .B1(new_n531), .B2(new_n532), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n909), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(G168), .A2(G171), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n531), .A2(new_n532), .A3(G301), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n858), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n912), .A2(new_n914), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n950), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n950), .A2(new_n953), .B1(new_n917), .B2(new_n920), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT107), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n939), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n950), .A2(new_n953), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n921), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n950), .A2(new_n953), .A3(new_n954), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n957), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n955), .A2(new_n956), .ZN(new_n965));
  AOI21_X1  g540(.A(G37), .B1(new_n965), .B2(new_n939), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n947), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT109), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n920), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n918), .A2(KEYINPUT109), .A3(new_n919), .A4(new_n913), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n917), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n959), .A3(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n972), .A2(new_n959), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n962), .A2(KEYINPUT110), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n958), .B(new_n974), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n966), .ZN(new_n978));
  OAI22_X1  g553(.A1(new_n967), .A2(new_n968), .B1(new_n978), .B2(KEYINPUT43), .ZN(new_n979));
  AOI211_X1 g554(.A(KEYINPUT108), .B(new_n947), .C1(new_n964), .C2(new_n966), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n979), .A2(KEYINPUT44), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n964), .A2(new_n966), .A3(new_n947), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n983), .A2(KEYINPUT111), .B1(new_n978), .B2(KEYINPUT43), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n983), .A2(KEYINPUT111), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n981), .A2(new_n986), .ZN(G397));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n503), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n464), .B(G40), .C1(new_n471), .C2(new_n472), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n770), .B(new_n773), .ZN(new_n994));
  INV_X1    g569(.A(G1996), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n815), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n737), .A2(new_n739), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n737), .A2(new_n739), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n994), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n601), .B(G1986), .Z(new_n1000));
  OAI21_X1  g575(.A(new_n993), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n992), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n991), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1966), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n503), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n494), .A2(new_n496), .ZN(new_n1009));
  OAI211_X1 g584(.A(G126), .B(G2105), .C1(new_n459), .C2(new_n460), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n500), .B2(new_n492), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n490), .A2(new_n491), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1013), .A2(KEYINPUT4), .A3(new_n501), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1384), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1002), .B(new_n1008), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  OAI22_X1  g592(.A1(new_n1006), .A2(KEYINPUT117), .B1(G2084), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT45), .B1(new_n503), .B2(new_n988), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(new_n992), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1966), .B1(new_n1020), .B2(new_n1003), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(G8), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G168), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT51), .B1(new_n1026), .B2(KEYINPUT125), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1024), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1016), .B1(new_n503), .B2(new_n988), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1007), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1031), .A2(new_n1033), .A3(new_n992), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1021), .A2(new_n1022), .B1(new_n830), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1006), .A2(KEYINPUT117), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(G8), .B(new_n1028), .C1(new_n1037), .C2(G286), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1026), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(KEYINPUT124), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT124), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n1037), .B2(new_n1026), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1030), .B(new_n1038), .C1(new_n1040), .C2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT62), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1039), .A2(KEYINPUT124), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1037), .A2(new_n1041), .A3(new_n1026), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT62), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(new_n1030), .A4(new_n1038), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n722), .A2(G1976), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1050), .B(G8), .C1(new_n989), .C2(new_n992), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT52), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT49), .ZN(new_n1053));
  OAI21_X1  g628(.A(G1981), .B1(new_n590), .B2(new_n593), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n590), .A2(new_n593), .A3(G1981), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1015), .A2(new_n1002), .ZN(new_n1058));
  INV_X1    g633(.A(G1981), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n594), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1060), .A2(KEYINPUT49), .A3(new_n1054), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1057), .A2(new_n1058), .A3(new_n1061), .A4(G8), .ZN(new_n1062));
  INV_X1    g637(.A(G1976), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT52), .B1(G288), .B2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1058), .A2(G8), .A3(new_n1050), .A4(new_n1064), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1052), .A2(new_n1062), .A3(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT112), .B(G1971), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n1020), .B2(new_n1003), .ZN(new_n1068));
  NOR4_X1   g643(.A1(new_n1031), .A2(new_n1033), .A3(G2090), .A4(new_n992), .ZN(new_n1069));
  OAI21_X1  g644(.A(G8), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AND2_X1   g645(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1071));
  NOR2_X1   g646(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1072));
  OAI22_X1  g647(.A1(G166), .A2(new_n1025), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1072), .ZN(new_n1074));
  NAND3_X1  g649(.A1(G303), .A2(G8), .A3(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1073), .A2(new_n1075), .A3(KEYINPUT114), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT114), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1066), .B1(new_n1070), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1067), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1004), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n992), .B1(new_n989), .B2(KEYINPUT50), .ZN(new_n1082));
  INV_X1    g657(.A(G2090), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT115), .B1(new_n503), .B2(new_n1007), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n503), .A2(KEYINPUT115), .A3(new_n1007), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1082), .B(new_n1083), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1081), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT116), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1081), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(G8), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1079), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1095), .A2(new_n1019), .A3(new_n992), .ZN(new_n1096));
  INV_X1    g671(.A(G2078), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT53), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(G2078), .ZN(new_n1100));
  AND4_X1   g675(.A1(new_n991), .A2(new_n1002), .A3(new_n1003), .A4(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(G1961), .B1(new_n1082), .B2(new_n1008), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT126), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1020), .A2(new_n1003), .A3(new_n1100), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1017), .A2(new_n775), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT126), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1098), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1108), .A2(G301), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1094), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1044), .A2(new_n1049), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n989), .A2(KEYINPUT50), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1112), .B(new_n1002), .C1(new_n1085), .C2(new_n1084), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n758), .A2(new_n1113), .B1(new_n1096), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n540), .A2(G91), .ZN(new_n1118));
  INV_X1    g693(.A(new_n577), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n576), .B1(new_n543), .B2(new_n573), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n566), .ZN(new_n1122));
  OAI21_X1  g697(.A(G65), .B1(new_n1122), .B2(new_n564), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n507), .B1(new_n1123), .B2(new_n569), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1117), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n571), .A2(new_n578), .A3(new_n1116), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT120), .B1(new_n1115), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT115), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1008), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n503), .A2(KEYINPUT115), .A3(new_n1007), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(G1956), .B1(new_n1133), .B2(new_n1082), .ZN(new_n1134));
  AND4_X1   g709(.A1(new_n991), .A2(new_n1002), .A3(new_n1003), .A4(new_n1114), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n1136));
  NOR4_X1   g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .A4(new_n1127), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1129), .A2(new_n1137), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n989), .A2(G2067), .A3(new_n992), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1034), .B2(G1348), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n617), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1127), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1138), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n616), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(G1348), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1139), .B1(new_n1017), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1148), .A2(new_n1149), .A3(KEYINPUT60), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1148), .B2(KEYINPUT60), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1146), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n991), .A2(new_n995), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1153));
  XOR2_X1   g728(.A(KEYINPUT58), .B(G1341), .Z(new_n1154));
  NAND2_X1  g729(.A1(new_n1058), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n554), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT59), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  OAI211_X1 g733(.A(KEYINPUT60), .B(new_n1140), .C1(new_n1034), .C2(G1348), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT123), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n617), .B1(new_n1148), .B2(KEYINPUT60), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1148), .A2(new_n1149), .A3(KEYINPUT60), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1113), .A2(new_n758), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1096), .A2(new_n1114), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1164), .A2(new_n1165), .A3(new_n1128), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1143), .A2(new_n1166), .A3(KEYINPUT61), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1152), .A2(new_n1158), .A3(new_n1163), .A4(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1143), .B1(new_n1129), .B2(new_n1137), .ZN(new_n1169));
  XOR2_X1   g744(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1168), .B1(new_n1171), .B2(KEYINPUT122), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1169), .A2(new_n1173), .A3(new_n1170), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1144), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1099), .B1(new_n1004), .B2(G2078), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1101), .A2(new_n1102), .A3(KEYINPUT126), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1106), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1178));
  OAI211_X1 g753(.A(G301), .B(new_n1176), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1176), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1180), .B1(new_n1181), .B2(G171), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1079), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1176), .A2(G301), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1187), .B1(new_n1108), .B2(G301), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1188), .A2(KEYINPUT127), .A3(new_n1180), .ZN(new_n1189));
  AOI21_X1  g764(.A(KEYINPUT127), .B1(new_n1188), .B2(new_n1180), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n1043), .B(new_n1186), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1111), .B1(new_n1175), .B2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g767(.A(G8), .B(G168), .C1(new_n1018), .C2(new_n1023), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1034), .A2(new_n1083), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1025), .B1(new_n1194), .B2(new_n1081), .ZN(new_n1195));
  OAI21_X1  g770(.A(KEYINPUT63), .B1(new_n1195), .B2(new_n1092), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1193), .A2(new_n1196), .A3(new_n1079), .ZN(new_n1197));
  AOI211_X1 g772(.A(new_n1025), .B(G286), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1184), .A2(new_n1185), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT63), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1197), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI211_X1 g776(.A(new_n1066), .B(new_n1195), .C1(new_n1077), .C2(new_n1076), .ZN(new_n1202));
  AND3_X1   g777(.A1(new_n1062), .A2(new_n1063), .A3(new_n722), .ZN(new_n1203));
  OAI211_X1 g778(.A(G8), .B(new_n1058), .C1(new_n1203), .C2(new_n1056), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(KEYINPUT118), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1205), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT118), .ZN(new_n1208));
  AOI21_X1  g783(.A(KEYINPUT63), .B1(new_n1094), .B2(new_n1198), .ZN(new_n1209));
  OAI211_X1 g784(.A(new_n1207), .B(new_n1208), .C1(new_n1209), .C2(new_n1197), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1206), .A2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1001), .B1(new_n1192), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n994), .A2(new_n996), .ZN(new_n1213));
  OAI22_X1  g788(.A1(new_n1213), .A2(new_n997), .B1(G2067), .B2(new_n770), .ZN(new_n1214));
  AND2_X1   g789(.A1(new_n1214), .A2(new_n993), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n993), .A2(new_n995), .ZN(new_n1216));
  XOR2_X1   g791(.A(new_n1216), .B(KEYINPUT46), .Z(new_n1217));
  INV_X1    g792(.A(new_n993), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1218), .B1(new_n994), .B2(new_n816), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n1220), .B(KEYINPUT47), .ZN(new_n1221));
  OR3_X1    g796(.A1(new_n1218), .A2(G1986), .A3(G290), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT48), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1225), .B1(new_n999), .B2(new_n993), .ZN(new_n1226));
  AOI211_X1 g801(.A(new_n1215), .B(new_n1221), .C1(new_n1224), .C2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1212), .A2(new_n1227), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g803(.A1(new_n682), .A2(G319), .ZN(new_n1230));
  AND3_X1   g804(.A1(new_n708), .A2(new_n663), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g805(.A(new_n893), .ZN(new_n1232));
  OAI21_X1  g806(.A(new_n894), .B1(new_n892), .B2(KEYINPUT103), .ZN(new_n1233));
  OAI21_X1  g807(.A(new_n897), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g808(.A(G37), .ZN(new_n1235));
  NAND2_X1  g809(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g810(.A(new_n897), .ZN(new_n1237));
  AND4_X1   g811(.A1(KEYINPUT104), .A2(new_n889), .A3(new_n900), .A4(new_n1237), .ZN(new_n1238));
  AOI21_X1  g812(.A(KEYINPUT104), .B1(new_n899), .B2(new_n900), .ZN(new_n1239));
  NOR2_X1   g813(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g814(.A(new_n1231), .B1(new_n1236), .B2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g815(.A1(new_n979), .A2(new_n980), .ZN(new_n1242));
  NOR2_X1   g816(.A1(new_n1241), .A2(new_n1242), .ZN(G308));
  OAI221_X1 g817(.A(new_n1231), .B1(new_n979), .B2(new_n980), .C1(new_n1240), .C2(new_n1236), .ZN(G225));
endmodule


