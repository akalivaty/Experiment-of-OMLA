//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n204));
  INV_X1    g0004(.A(G87), .ZN(new_n205));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G257), .ZN(new_n208));
  OAI221_X1 g0008(.A(new_n204), .B1(new_n205), .B2(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(KEYINPUT67), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n209), .A2(new_n210), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n203), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT68), .Z(new_n217));
  INV_X1    g0017(.A(KEYINPUT1), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT64), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n221), .B1(new_n203), .B2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G13), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n223), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT65), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(G50), .B1(G58), .B2(G68), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT66), .Z(new_n234));
  AOI21_X1  g0034(.A(new_n227), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  AND3_X1   g0035(.A1(new_n219), .A2(new_n220), .A3(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(KEYINPUT76), .ZN(new_n252));
  INV_X1    g0052(.A(G226), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G232), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G1698), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n255), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G97), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G41), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  AOI21_X1  g0066(.A(G1), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G1), .A3(G13), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(new_n269), .A3(G274), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(G238), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT13), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n264), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT73), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n269), .B1(new_n260), .B2(new_n261), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n270), .A2(new_n273), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT13), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n264), .A2(new_n274), .A3(KEYINPUT73), .A4(new_n275), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n278), .A2(G179), .A3(new_n281), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n276), .A2(new_n281), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT14), .B1(new_n284), .B2(G169), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT14), .ZN(new_n286));
  INV_X1    g0086(.A(G169), .ZN(new_n287));
  AOI211_X1 g0087(.A(new_n286), .B(new_n287), .C1(new_n276), .C2(new_n281), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n283), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n271), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT72), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n271), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT12), .B1(new_n294), .B2(G68), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n223), .A2(G1), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT12), .ZN(new_n297));
  INV_X1    g0097(.A(G68), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n296), .A2(new_n297), .A3(G20), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n228), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(new_n292), .B2(new_n293), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n271), .A2(G20), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(G68), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n229), .A2(G33), .A3(G77), .ZN(new_n306));
  NOR2_X1   g0106(.A1(G20), .A2(G33), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G50), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n306), .B1(new_n229), .B2(G68), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT11), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n310), .A2(new_n311), .A3(new_n302), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n310), .B2(new_n302), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n300), .B(new_n305), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n289), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n304), .ZN(new_n316));
  INV_X1    g0116(.A(G77), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n303), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(G77), .B2(new_n294), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G20), .A2(G77), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT8), .B(G58), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(new_n308), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT15), .B(G87), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n229), .A2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n302), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT71), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI221_X1 g0129(.A(new_n321), .B1(new_n322), .B2(new_n308), .C1(new_n325), .C2(new_n324), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n330), .A2(KEYINPUT71), .A3(new_n302), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n320), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n269), .A2(G244), .A3(new_n272), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n270), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n258), .A2(new_n259), .ZN(new_n336));
  INV_X1    g0136(.A(G107), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n269), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n256), .A2(new_n254), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(G238), .B2(new_n254), .ZN(new_n340));
  OR2_X1    g0140(.A1(KEYINPUT3), .A2(G33), .ZN(new_n341));
  NAND2_X1  g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n335), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G200), .ZN(new_n347));
  INV_X1    g0147(.A(G190), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n332), .B(new_n347), .C1(new_n348), .C2(new_n346), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n331), .A2(new_n329), .ZN(new_n350));
  INV_X1    g0150(.A(new_n320), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n346), .A2(new_n287), .ZN(new_n353));
  INV_X1    g0153(.A(G179), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n335), .A2(new_n345), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G200), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(new_n276), .B2(new_n281), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(new_n314), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n278), .A2(G190), .A3(new_n281), .A4(new_n282), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n315), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  XOR2_X1   g0163(.A(KEYINPUT8), .B(G58), .Z(new_n364));
  INV_X1    g0164(.A(KEYINPUT75), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(new_n304), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n290), .A2(new_n228), .A3(new_n301), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT75), .B1(new_n322), .B2(new_n316), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n290), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n322), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n343), .B2(G20), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n336), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n298), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G58), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(new_n298), .ZN(new_n381));
  NOR2_X1   g0181(.A1(G58), .A2(G68), .ZN(new_n382));
  OAI21_X1  g0182(.A(G20), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n307), .A2(G159), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n375), .B1(new_n379), .B2(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n301), .A2(new_n228), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT7), .B1(new_n336), .B2(new_n229), .ZN(new_n388));
  NOR4_X1   g0188(.A1(new_n258), .A2(new_n259), .A3(new_n376), .A4(G20), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n384), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n387), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n373), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(G223), .B(new_n254), .C1(new_n258), .C2(new_n259), .ZN(new_n395));
  OAI211_X1 g0195(.A(G226), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n396));
  INV_X1    g0196(.A(G33), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n395), .B(new_n396), .C1(new_n397), .C2(new_n205), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n263), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n269), .A2(new_n272), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n270), .B1(new_n256), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n348), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n401), .B1(new_n263), .B2(new_n398), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(G200), .B2(new_n404), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n394), .A2(KEYINPUT17), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT17), .B1(new_n394), .B2(new_n405), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n399), .A2(new_n354), .A3(new_n402), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(G169), .B2(new_n404), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n409), .B1(new_n394), .B2(new_n411), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n399), .A2(new_n354), .A3(new_n402), .ZN(new_n413));
  AOI21_X1  g0213(.A(G169), .B1(new_n399), .B2(new_n402), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n373), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n302), .B1(new_n379), .B2(new_n391), .ZN(new_n417));
  INV_X1    g0217(.A(new_n385), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n374), .B1(new_n390), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n416), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n415), .A2(new_n420), .A3(KEYINPUT18), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n412), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n408), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n363), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n270), .B1(new_n253), .B2(new_n400), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n336), .A2(G77), .ZN(new_n426));
  OAI211_X1 g0226(.A(G222), .B(new_n254), .C1(new_n258), .C2(new_n259), .ZN(new_n427));
  OAI211_X1 g0227(.A(G223), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n269), .B1(new_n429), .B2(KEYINPUT69), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT69), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n426), .A2(new_n431), .A3(new_n427), .A4(new_n428), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n425), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n433), .A2(new_n354), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n304), .A2(G50), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n367), .A2(new_n435), .B1(G50), .B2(new_n290), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT70), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n371), .A2(new_n309), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(KEYINPUT70), .C1(new_n367), .C2(new_n435), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G150), .ZN(new_n442));
  OAI22_X1  g0242(.A1(new_n322), .A2(new_n325), .B1(new_n442), .B2(new_n308), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n229), .B1(new_n382), .B2(new_n309), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n302), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n433), .B2(G169), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n434), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n429), .A2(KEYINPUT69), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(new_n432), .A3(new_n263), .ZN(new_n450));
  INV_X1    g0250(.A(new_n425), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n358), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n440), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n387), .A2(G50), .A3(new_n290), .A4(new_n304), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT70), .B1(new_n454), .B2(new_n439), .ZN(new_n455));
  OAI211_X1 g0255(.A(KEYINPUT9), .B(new_n445), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT9), .B1(new_n441), .B2(new_n445), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n452), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT10), .ZN(new_n460));
  AOI211_X1 g0260(.A(new_n348), .B(new_n425), .C1(new_n430), .C2(new_n432), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT9), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n446), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n465), .B(new_n456), .C1(new_n358), .C2(new_n433), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT10), .B1(new_n466), .B2(new_n461), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n448), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n252), .B1(new_n424), .B2(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n289), .A2(new_n314), .B1(new_n361), .B2(new_n360), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n470), .A2(new_n408), .A3(new_n422), .A4(new_n357), .ZN(new_n471));
  INV_X1    g0271(.A(new_n448), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n460), .B1(new_n459), .B2(new_n462), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n465), .A2(new_n456), .ZN(new_n474));
  NOR4_X1   g0274(.A1(new_n474), .A2(new_n461), .A3(KEYINPUT10), .A4(new_n452), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n472), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n471), .A2(new_n476), .A3(KEYINPUT76), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(G97), .A2(G107), .ZN(new_n479));
  NOR2_X1   g0279(.A1(G97), .A2(G107), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n479), .A2(new_n480), .B1(KEYINPUT77), .B2(KEYINPUT6), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(KEYINPUT6), .B2(new_n207), .ZN(new_n483));
  XNOR2_X1  g0283(.A(G97), .B(G107), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n481), .B(G20), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n307), .A2(G77), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n337), .B1(new_n377), .B2(new_n378), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n302), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n290), .A2(G97), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n397), .A2(G1), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n367), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n490), .B1(new_n492), .B2(G97), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G250), .A2(G1698), .ZN(new_n494));
  NAND2_X1  g0294(.A1(KEYINPUT4), .A2(G244), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(G1698), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n343), .A2(new_n496), .B1(G33), .B2(G283), .ZN(new_n497));
  OAI211_X1 g0297(.A(G244), .B(new_n254), .C1(new_n258), .C2(new_n259), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n269), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n271), .A2(G45), .ZN(new_n503));
  OR2_X1    g0303(.A1(KEYINPUT5), .A2(G41), .ZN(new_n504));
  NAND2_X1  g0304(.A1(KEYINPUT5), .A2(G41), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G274), .ZN(new_n507));
  INV_X1    g0307(.A(new_n228), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n268), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n266), .A2(G1), .ZN(new_n511));
  AND2_X1   g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  NOR2_X1   g0312(.A1(KEYINPUT5), .A2(G41), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n269), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n510), .B1(new_n515), .B2(new_n208), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(G200), .B1(new_n502), .B2(new_n517), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n501), .A2(new_n516), .A3(G190), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n489), .B(new_n493), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n489), .A2(new_n493), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n287), .B1(new_n501), .B2(new_n516), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n501), .A2(new_n516), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n354), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(G244), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n527));
  OAI211_X1 g0327(.A(G238), .B(new_n254), .C1(new_n258), .C2(new_n259), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G116), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n263), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n503), .A2(G250), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n269), .A2(new_n533), .B1(new_n509), .B2(new_n511), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G200), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT19), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n229), .B1(new_n261), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n480), .A2(new_n205), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n229), .B(G68), .C1(new_n258), .C2(new_n259), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n537), .B1(new_n325), .B2(new_n207), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n302), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n292), .A2(new_n324), .A3(new_n293), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n492), .A2(G87), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n531), .A2(G190), .A3(new_n534), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n536), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OR3_X1    g0349(.A1(new_n367), .A2(new_n324), .A3(new_n491), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n544), .A2(new_n550), .A3(new_n545), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n531), .A2(new_n354), .A3(new_n534), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n269), .A2(G274), .ZN(new_n553));
  OAI22_X1  g0353(.A1(new_n553), .A2(new_n503), .B1(new_n263), .B2(new_n532), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n263), .B2(new_n530), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n551), .B(new_n552), .C1(G169), .C2(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n206), .A2(new_n254), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n208), .A2(G1698), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n558), .B(new_n559), .C1(new_n258), .C2(new_n259), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G33), .A2(G294), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n269), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n514), .A2(G264), .A3(new_n269), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n564), .A3(new_n510), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(G190), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT80), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(KEYINPUT79), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT79), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n514), .A2(new_n569), .A3(G264), .A4(new_n269), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n567), .B1(new_n571), .B2(new_n563), .ZN(new_n572));
  AOI211_X1 g0372(.A(KEYINPUT80), .B(new_n562), .C1(new_n568), .C2(new_n570), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n510), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n566), .B1(new_n574), .B2(new_n358), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n229), .B(G87), .C1(new_n258), .C2(new_n259), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT22), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT22), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n343), .A2(new_n578), .A3(new_n229), .A4(G87), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT24), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n529), .A2(G20), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT23), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n229), .B2(G107), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n337), .A2(KEYINPUT23), .A3(G20), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n580), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n581), .B1(new_n580), .B2(new_n586), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n302), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n371), .A2(new_n337), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n590), .B(KEYINPUT25), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(G107), .B2(new_n492), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n526), .B(new_n557), .C1(new_n575), .C2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n354), .B1(new_n506), .B2(new_n509), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n572), .B2(new_n573), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n565), .A2(G169), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n596), .A2(new_n597), .B1(new_n589), .B2(new_n592), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT21), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n491), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n294), .A2(new_n387), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n292), .A2(new_n600), .A3(new_n293), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n600), .A2(G20), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n302), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(G20), .B1(G33), .B2(G283), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n397), .A2(G97), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT78), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT78), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n608), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n607), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT20), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n612), .B1(new_n608), .B2(new_n609), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n606), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(KEYINPUT20), .A3(new_n613), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n604), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(G303), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n341), .A2(new_n621), .A3(new_n342), .ZN(new_n622));
  MUX2_X1   g0422(.A(G257), .B(G264), .S(G1698), .Z(new_n623));
  OAI211_X1 g0423(.A(new_n263), .B(new_n622), .C1(new_n623), .C2(new_n336), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n514), .A2(G270), .A3(new_n269), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n510), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G169), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n599), .B1(new_n620), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n602), .A2(new_n603), .ZN(new_n629));
  AND4_X1   g0429(.A1(KEYINPUT20), .A2(new_n607), .A3(new_n613), .A4(new_n611), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT20), .B1(new_n618), .B2(new_n613), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n627), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n633), .A3(KEYINPUT21), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n626), .A2(new_n348), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n626), .A2(G200), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n620), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n595), .A2(new_n624), .A3(new_n625), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n628), .A2(new_n634), .A3(new_n637), .A4(new_n639), .ZN(new_n640));
  NOR4_X1   g0440(.A1(new_n478), .A2(new_n594), .A3(new_n598), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(KEYINPUT81), .ZN(G372));
  NAND2_X1  g0442(.A1(new_n463), .A2(new_n467), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n353), .A2(new_n355), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n332), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n362), .A2(new_n645), .ZN(new_n646));
  AOI211_X1 g0446(.A(new_n407), .B(new_n406), .C1(new_n315), .C2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT83), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n422), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n412), .A2(new_n421), .A3(KEYINPUT83), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n643), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n472), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT26), .B1(new_n557), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n549), .A2(new_n556), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n657), .A2(new_n525), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n556), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n628), .A2(new_n634), .A3(new_n639), .ZN(new_n661));
  AOI221_X4 g0461(.A(KEYINPUT82), .B1(new_n589), .B2(new_n592), .C1(new_n596), .C2(new_n597), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT82), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n596), .A2(new_n597), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(new_n593), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n661), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n575), .A2(new_n593), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n557), .A2(new_n520), .A3(new_n525), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n660), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n654), .B1(new_n478), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g0471(.A(new_n671), .B(KEYINPUT84), .Z(G369));
  NAND2_X1  g0472(.A1(new_n296), .A2(new_n229), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n620), .A2(new_n679), .ZN(new_n680));
  MUX2_X1   g0480(.A(new_n640), .B(new_n661), .S(new_n680), .Z(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT85), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  INV_X1    g0483(.A(new_n595), .ZN(new_n684));
  XNOR2_X1  g0484(.A(KEYINPUT5), .B(G41), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n685), .A2(new_n511), .B1(new_n508), .B2(new_n268), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n569), .B1(new_n686), .B2(G264), .ZN(new_n687));
  INV_X1    g0487(.A(new_n570), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n563), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT80), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n571), .A2(new_n567), .A3(new_n563), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n684), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n597), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n593), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n593), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(new_n679), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n667), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n598), .A2(new_n678), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n683), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n661), .A2(new_n678), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n697), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n694), .A2(KEYINPUT82), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n598), .A2(new_n663), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n704), .B1(new_n707), .B2(new_n678), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n702), .A2(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n225), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n710), .A2(KEYINPUT87), .A3(G41), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT87), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n225), .B2(new_n265), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n480), .A2(new_n205), .A3(new_n600), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT86), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(G1), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n233), .B2(new_n715), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n572), .A2(new_n573), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n523), .A2(new_n638), .A3(new_n555), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n690), .A2(new_n691), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n523), .A2(new_n638), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(KEYINPUT30), .A4(new_n555), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n626), .A2(new_n354), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n523), .A2(new_n729), .A3(new_n555), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n574), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n725), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n678), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n598), .A2(new_n640), .ZN(new_n736));
  AOI21_X1  g0536(.A(G200), .B1(new_n726), .B2(new_n510), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n695), .B1(new_n737), .B2(new_n566), .ZN(new_n738));
  AND4_X1   g0538(.A1(new_n520), .A2(new_n525), .A3(new_n556), .A4(new_n549), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n736), .A2(new_n738), .A3(new_n739), .A4(new_n679), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n735), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT29), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n670), .B2(new_n678), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n679), .A2(KEYINPUT29), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n694), .A2(new_n661), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(new_n738), .A3(new_n739), .ZN(new_n749));
  INV_X1    g0549(.A(new_n556), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n557), .A2(KEYINPUT26), .A3(new_n655), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n658), .B1(new_n657), .B2(new_n525), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n747), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n744), .B1(new_n746), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n721), .B1(new_n756), .B2(G1), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT88), .ZN(G364));
  INV_X1    g0558(.A(new_n683), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n223), .A2(G20), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n271), .B1(new_n760), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n714), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(G330), .B2(new_n682), .ZN(new_n765));
  INV_X1    g0565(.A(new_n763), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n228), .B1(G20), .B2(new_n287), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n348), .A2(new_n358), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n229), .A2(new_n354), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT90), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n348), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n229), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n777), .A2(G326), .B1(G294), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT92), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n358), .A2(G190), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n229), .A2(G179), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G283), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n336), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n770), .A2(G190), .A3(new_n358), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G190), .A2(G200), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n789), .A2(G322), .B1(new_n792), .B2(G329), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n769), .A2(new_n784), .ZN(new_n794));
  INV_X1    g0594(.A(G311), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n770), .A2(new_n790), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n793), .B1(new_n621), .B2(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n770), .A2(new_n783), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n798), .A2(KEYINPUT91), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(KEYINPUT91), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT33), .B(G317), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n787), .B(new_n797), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n782), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT32), .ZN(new_n806));
  INV_X1    g0606(.A(G159), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n791), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n792), .A2(KEYINPUT32), .A3(G159), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n777), .A2(G50), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n785), .A2(new_n337), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n794), .A2(new_n205), .ZN(new_n812));
  INV_X1    g0612(.A(new_n796), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n811), .B(new_n812), .C1(G77), .C2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n779), .A2(new_n207), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n336), .B(new_n815), .C1(G58), .C2(new_n789), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n802), .A2(G68), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n810), .A2(new_n814), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n768), .B1(new_n805), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G13), .A2(G33), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(G20), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n767), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n710), .A2(new_n343), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n266), .B2(new_n234), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n247), .A2(new_n266), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n225), .A2(G355), .A3(new_n343), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(G116), .B2(new_n225), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n826), .A2(new_n827), .B1(KEYINPUT89), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(KEYINPUT89), .B2(new_n829), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n766), .B(new_n819), .C1(new_n823), .C2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n822), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n682), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n765), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G396));
  NAND2_X1  g0636(.A1(new_n352), .A2(new_n678), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n357), .A2(KEYINPUT93), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n349), .A2(new_n356), .A3(new_n837), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT93), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n594), .B1(new_n707), .B2(new_n661), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n679), .B(new_n842), .C1(new_n843), .C2(new_n660), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n670), .A2(new_n678), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n838), .B(new_n841), .C1(new_n356), .C2(new_n679), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n763), .B1(new_n847), .B2(new_n743), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n743), .B2(new_n847), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n767), .A2(new_n820), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n763), .B1(G77), .B2(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n777), .A2(G303), .B1(new_n802), .B2(G283), .ZN(new_n853));
  INV_X1    g0653(.A(new_n794), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G116), .A2(new_n813), .B1(new_n854), .B2(G107), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n789), .A2(G294), .B1(new_n792), .B2(G311), .ZN(new_n856));
  INV_X1    g0656(.A(new_n785), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n343), .B(new_n815), .C1(G87), .C2(new_n857), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n853), .A2(new_n855), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n789), .A2(G143), .B1(new_n813), .B2(G159), .ZN(new_n860));
  INV_X1    g0660(.A(G137), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n860), .B1(new_n801), .B2(new_n442), .C1(new_n776), .C2(new_n861), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT34), .Z(new_n863));
  AOI22_X1  g0663(.A1(new_n857), .A2(G68), .B1(new_n792), .B2(G132), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n336), .B1(new_n854), .B2(G50), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n864), .B(new_n865), .C1(new_n380), .C2(new_n779), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n859), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n852), .B1(new_n867), .B2(new_n767), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n846), .B2(new_n821), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n849), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT94), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n849), .A2(KEYINPUT94), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(G384));
  INV_X1    g0674(.A(KEYINPUT35), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n232), .B(G116), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n875), .B2(new_n876), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT36), .Z(new_n879));
  OAI21_X1  g0679(.A(G77), .B1(new_n380), .B2(new_n298), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n880), .A2(new_n233), .B1(G50), .B2(new_n298), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(G1), .A3(new_n223), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT95), .Z(new_n884));
  INV_X1    g0684(.A(KEYINPUT98), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n314), .A2(new_n678), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n360), .A2(new_n361), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n887), .B1(new_n888), .B2(new_n289), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT97), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n470), .A2(new_n886), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT97), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n892), .B(new_n887), .C1(new_n888), .C2(new_n289), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n676), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n420), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n423), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n415), .A2(new_n420), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n394), .A2(new_n405), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT37), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n899), .A2(new_n896), .A3(new_n900), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  INV_X1    g0707(.A(new_n905), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n896), .B1(new_n408), .B2(new_n422), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n645), .A2(new_n679), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT96), .Z(new_n912));
  AOI221_X4 g0712(.A(new_n894), .B1(new_n906), .B2(new_n910), .C1(new_n844), .C2(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n412), .A2(new_n421), .A3(KEYINPUT83), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT83), .B1(new_n412), .B2(new_n421), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n916), .A2(new_n895), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n885), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n908), .A2(new_n907), .A3(new_n909), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT38), .B1(new_n898), .B2(new_n905), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n648), .B1(new_n394), .B2(new_n411), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n415), .A2(new_n420), .A3(KEYINPUT83), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n923), .A2(new_n924), .A3(new_n900), .A4(new_n896), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT37), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(KEYINPUT99), .A3(new_n904), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT99), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n925), .A2(new_n928), .A3(KEYINPUT37), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n896), .B1(new_n916), .B2(new_n408), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n907), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n906), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n922), .B1(new_n933), .B2(new_n921), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n315), .A2(new_n678), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n917), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n844), .A2(new_n912), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n919), .A2(new_n920), .ZN(new_n941));
  OAI211_X1 g0741(.A(KEYINPUT98), .B(new_n937), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n918), .A2(new_n936), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT76), .B1(new_n471), .B2(new_n476), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n315), .A2(new_n357), .A3(new_n362), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n408), .A2(new_n422), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n945), .A2(new_n468), .A3(new_n946), .A4(new_n252), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n754), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n653), .B1(new_n948), .B2(new_n746), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n943), .B(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT40), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n932), .B2(new_n906), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n741), .A2(KEYINPUT100), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT100), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n732), .A2(new_n954), .A3(KEYINPUT31), .A4(new_n678), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n953), .A2(new_n735), .A3(new_n740), .A4(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(new_n846), .A3(new_n939), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT101), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT101), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n956), .A2(new_n959), .A3(new_n846), .A4(new_n939), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n952), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n951), .B1(new_n957), .B2(new_n941), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n956), .B1(new_n469), .B2(new_n477), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(G330), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n950), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n271), .B2(new_n760), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n950), .A2(new_n967), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n884), .B1(new_n969), .B2(new_n970), .ZN(G367));
  INV_X1    g0771(.A(new_n702), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n521), .A2(new_n678), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n526), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n655), .A2(new_n678), .ZN(new_n975));
  AND3_X1   g0775(.A1(new_n974), .A2(KEYINPUT105), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT105), .B1(new_n974), .B2(new_n975), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n972), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(KEYINPUT42), .B1(new_n978), .B2(new_n704), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n978), .A2(KEYINPUT42), .A3(new_n704), .ZN(new_n981));
  INV_X1    g0781(.A(new_n978), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n655), .B1(new_n982), .B2(new_n598), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n980), .B(new_n981), .C1(new_n983), .C2(new_n678), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(KEYINPUT106), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(KEYINPUT106), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n679), .A2(new_n547), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n557), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n990), .A2(KEYINPUT102), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(KEYINPUT102), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n991), .B(new_n992), .C1(new_n556), .C2(new_n989), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT103), .Z(new_n994));
  MUX2_X1   g0794(.A(new_n988), .B(KEYINPUT43), .S(new_n994), .Z(new_n995));
  NAND2_X1  g0795(.A1(new_n987), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n994), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n998), .A2(new_n988), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n987), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n979), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n996), .B1(new_n972), .B2(new_n978), .C1(new_n999), .C2(new_n987), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n714), .B(KEYINPUT41), .Z(new_n1003));
  NAND2_X1  g0803(.A1(new_n708), .A2(new_n978), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT44), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT45), .ZN(new_n1007));
  OR3_X1    g0807(.A1(new_n708), .A2(new_n1007), .A3(new_n978), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1007), .B1(new_n708), .B2(new_n978), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT107), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n972), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n704), .B1(new_n700), .B2(new_n703), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n683), .B(new_n1014), .Z(new_n1015));
  NAND2_X1  g0815(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1016), .A2(KEYINPUT107), .A3(new_n702), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1013), .A2(new_n756), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1003), .B1(new_n1018), .B2(new_n756), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1001), .B(new_n1002), .C1(new_n1019), .C2(new_n762), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n823), .B1(new_n225), .B2(new_n324), .C1(new_n825), .C2(new_n243), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1021), .A2(new_n763), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n789), .A2(G150), .B1(new_n854), .B2(G58), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n861), .B2(new_n791), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n779), .A2(new_n298), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n343), .B1(new_n785), .B2(new_n317), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n801), .A2(new_n807), .B1(new_n309), .B2(new_n796), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(KEYINPUT109), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n777), .A2(G143), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1028), .A2(KEYINPUT109), .ZN(new_n1032));
  INV_X1    g0832(.A(G294), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n776), .A2(new_n795), .B1(new_n801), .B2(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n857), .A2(G97), .B1(new_n792), .B2(G317), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n336), .C1(new_n621), .C2(new_n788), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n794), .A2(new_n600), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT46), .ZN(new_n1038));
  OR3_X1    g0838(.A1(new_n1034), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n779), .A2(new_n337), .B1(new_n796), .B2(new_n786), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT108), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n1031), .A2(new_n1032), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1022), .B1(new_n768), .B2(new_n1044), .C1(new_n994), .C2(new_n833), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1020), .A2(new_n1045), .ZN(G387));
  NAND3_X1  g0846(.A1(new_n717), .A2(new_n225), .A3(new_n343), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(G107), .B2(new_n225), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT111), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n322), .A2(G50), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1050), .B(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n718), .A3(new_n1053), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1054), .B(new_n824), .C1(new_n240), .C2(new_n266), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1049), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n766), .B1(new_n1056), .B2(new_n823), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT113), .Z(new_n1058));
  AOI22_X1  g0858(.A1(new_n789), .A2(G317), .B1(new_n813), .B2(G303), .ZN(new_n1059));
  INV_X1    g0859(.A(G322), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1059), .B1(new_n776), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G311), .B2(new_n802), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1062), .A2(KEYINPUT48), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1062), .A2(KEYINPUT48), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n779), .A2(new_n786), .B1(new_n794), .B2(new_n1033), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT49), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(KEYINPUT49), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n336), .B1(new_n785), .B2(new_n600), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G326), .B2(new_n792), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n777), .A2(G159), .B1(new_n802), .B2(new_n364), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n794), .A2(new_n317), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n796), .A2(new_n298), .B1(new_n791), .B2(new_n442), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(G50), .C2(new_n789), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n779), .A2(new_n324), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n336), .B(new_n1076), .C1(G97), .C2(new_n857), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1072), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n768), .B1(new_n1071), .B2(new_n1078), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1058), .B(new_n1079), .C1(new_n701), .C2(new_n822), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n1015), .B2(new_n762), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1015), .A2(new_n756), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n714), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1015), .A2(new_n756), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(G393));
  NOR2_X1   g0885(.A1(new_n1011), .A2(new_n972), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT114), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1016), .A2(new_n702), .ZN(new_n1088));
  OR3_X1    g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1087), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n762), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n823), .B1(new_n207), .B2(new_n225), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n250), .B2(new_n824), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n801), .A2(new_n309), .B1(new_n322), .B2(new_n796), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT116), .Z(new_n1095));
  AOI22_X1  g0895(.A1(G68), .A2(new_n854), .B1(new_n792), .B2(G143), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1096), .B(new_n343), .C1(new_n205), .C2(new_n785), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT115), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n779), .A2(new_n317), .ZN(new_n1099));
  OR3_X1    g0899(.A1(new_n1095), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n776), .A2(new_n442), .B1(new_n807), .B2(new_n788), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT51), .Z(new_n1102));
  AOI22_X1  g0902(.A1(new_n777), .A2(G317), .B1(G311), .B2(new_n789), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT52), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n336), .B1(new_n785), .B2(new_n337), .C1(new_n779), .C2(new_n600), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n794), .A2(new_n786), .B1(new_n791), .B2(new_n1060), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(G294), .C2(new_n813), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n621), .B2(new_n801), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n1100), .A2(new_n1102), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n766), .B(new_n1093), .C1(new_n1109), .C2(new_n767), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n982), .B2(new_n833), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1082), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1018), .A2(new_n1112), .A3(new_n714), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1091), .A2(new_n1111), .A3(new_n1113), .ZN(G390));
  NAND2_X1  g0914(.A1(new_n749), .A2(new_n753), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n678), .B1(new_n838), .B2(new_n841), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n912), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n939), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n935), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n933), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n742), .A2(G330), .A3(new_n846), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1122), .A2(new_n894), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n956), .A2(G330), .A3(new_n846), .A4(new_n939), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1123), .B1(KEYINPUT117), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1121), .B(new_n1125), .C1(new_n934), .C2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n649), .A2(new_n408), .A3(new_n650), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n897), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1129), .A2(new_n929), .A3(new_n927), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n919), .B1(new_n1130), .B2(new_n907), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n894), .B1(new_n1117), .B2(new_n912), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1131), .A2(new_n1132), .A3(new_n935), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n912), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n845), .B2(new_n842), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1120), .B1(new_n1135), .B2(new_n894), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n941), .A2(KEYINPUT39), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n1131), .B2(KEYINPUT39), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1133), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT117), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1124), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1127), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n948), .A2(new_n746), .ZN(new_n1144));
  OAI211_X1 g0944(.A(G330), .B(new_n956), .C1(new_n469), .C2(new_n477), .ZN(new_n1145));
  AND4_X1   g0945(.A1(KEYINPUT118), .A2(new_n1144), .A3(new_n654), .A4(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT118), .B1(new_n949), .B2(new_n1145), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1123), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n956), .A2(G330), .A3(new_n846), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1118), .B1(new_n1151), .B2(new_n894), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1122), .A2(new_n894), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1124), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1150), .A2(new_n1152), .B1(new_n1154), .B2(new_n938), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1143), .B1(new_n1149), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1121), .B1(new_n934), .B2(new_n1126), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n1141), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1154), .A2(new_n938), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1127), .A3(new_n1148), .A4(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1156), .A2(new_n1162), .A3(new_n714), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT119), .B1(new_n1143), .B2(new_n761), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT119), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1158), .A2(new_n1165), .A3(new_n762), .A4(new_n1127), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G97), .A2(new_n813), .B1(new_n792), .B2(G294), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n298), .B2(new_n785), .C1(new_n600), .C2(new_n788), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n1169), .A2(new_n343), .A3(new_n812), .A4(new_n1099), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n337), .B2(new_n801), .C1(new_n786), .C2(new_n776), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT54), .B(G143), .ZN(new_n1172));
  INV_X1    g0972(.A(G125), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n796), .A2(new_n1172), .B1(new_n791), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(G132), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n343), .B1(new_n788), .B2(new_n1175), .C1(new_n807), .C2(new_n779), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1174), .B(new_n1176), .C1(G50), .C2(new_n857), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n777), .A2(G128), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n854), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT53), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n794), .B2(new_n442), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n802), .A2(G137), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1177), .A2(new_n1178), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n768), .B1(new_n1171), .B2(new_n1183), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n766), .B(new_n1184), .C1(new_n322), .C2(new_n850), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT120), .Z(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n934), .B2(new_n821), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1163), .A2(new_n1167), .A3(new_n1187), .ZN(G378));
  NAND3_X1  g0988(.A1(new_n918), .A2(new_n936), .A3(new_n942), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n961), .A2(G330), .A3(new_n962), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n476), .A2(new_n446), .A3(new_n895), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n446), .A2(new_n895), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n468), .A2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1194), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1190), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT121), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1197), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1202), .A2(KEYINPUT121), .A3(new_n1195), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n961), .A2(new_n1204), .A3(G330), .A4(new_n962), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1189), .A2(new_n1199), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1189), .B1(new_n1205), .B2(new_n1199), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1148), .B1(new_n1143), .B2(new_n1155), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT57), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1199), .A2(new_n1205), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n943), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1210), .A2(new_n1213), .A3(KEYINPUT57), .A4(new_n1206), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n714), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1211), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1213), .A2(new_n762), .A3(new_n1206), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n763), .B1(G50), .B2(new_n851), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(G33), .A2(G41), .ZN(new_n1219));
  AOI211_X1 g1019(.A(G50), .B(new_n1219), .C1(new_n336), .C2(new_n265), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n777), .A2(G116), .B1(new_n802), .B2(G97), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n785), .A2(new_n380), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n788), .A2(new_n337), .B1(new_n796), .B2(new_n324), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(G283), .C2(new_n792), .ZN(new_n1224));
  NOR4_X1   g1024(.A1(new_n1025), .A2(new_n1073), .A3(G41), .A4(new_n343), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1221), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT58), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1220), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n789), .A2(G128), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n794), .B2(new_n1172), .C1(new_n861), .C2(new_n796), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n776), .A2(new_n1173), .B1(new_n801), .B2(new_n1175), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(G150), .C2(new_n780), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1233), .A2(KEYINPUT59), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1219), .B1(new_n785), .B2(new_n807), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G124), .B2(new_n792), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT59), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1236), .B1(new_n1232), .B2(new_n1237), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1228), .B1(new_n1227), .B2(new_n1226), .C1(new_n1234), .C2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1218), .B1(new_n1239), .B2(new_n767), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1204), .B2(new_n821), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1217), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1216), .A2(new_n1242), .ZN(G375));
  AOI21_X1  g1043(.A(new_n1003), .B1(new_n1148), .B2(new_n1161), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1148), .B2(new_n1161), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n761), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n894), .A2(new_n820), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n763), .B1(G68), .B2(new_n851), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n343), .B(new_n1076), .C1(G77), .C2(new_n857), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G107), .A2(new_n813), .B1(new_n854), .B2(G97), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n789), .A2(G283), .B1(new_n792), .B2(G303), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n776), .A2(new_n1033), .B1(new_n801), .B2(new_n600), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n336), .B(new_n1222), .C1(G50), .C2(new_n780), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G150), .A2(new_n813), .B1(new_n854), .B2(G159), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n789), .A2(G137), .B1(new_n792), .B2(G128), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n776), .A2(new_n1175), .B1(new_n801), .B2(new_n1172), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n1252), .A2(new_n1253), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1248), .B1(new_n1259), .B2(new_n767), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1247), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT122), .B1(new_n1246), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT122), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1264), .B(new_n1261), .C1(new_n1155), .C2(new_n761), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1245), .A2(new_n1266), .ZN(G381));
  AND2_X1   g1067(.A1(new_n1020), .A2(new_n1045), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1091), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1269));
  INV_X1    g1069(.A(G378), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n835), .B(new_n1081), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT123), .ZN(new_n1272));
  OR3_X1    g1072(.A1(new_n1271), .A2(G384), .A3(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1272), .B1(new_n1271), .B2(G384), .ZN(new_n1274));
  AOI21_X1  g1074(.A(G381), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .A4(new_n1275), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1276), .A2(G375), .ZN(G407));
  OAI21_X1  g1077(.A(G213), .B1(new_n1276), .B2(G375), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n677), .A2(G213), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(G375), .A2(G378), .A3(new_n1279), .ZN(new_n1280));
  OR3_X1    g1080(.A1(new_n1278), .A2(KEYINPUT124), .A3(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(KEYINPUT124), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(G409));
  INV_X1    g1083(.A(G2897), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1279), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT60), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n1148), .B2(new_n1161), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n715), .B1(new_n1148), .B2(new_n1161), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1155), .B(KEYINPUT60), .C1(new_n1147), .C2(new_n1146), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1288), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1291), .A2(G384), .A3(new_n1266), .ZN(new_n1292));
  AOI21_X1  g1092(.A(G384), .B1(new_n1291), .B2(new_n1266), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT125), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1292), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1291), .A2(new_n1266), .ZN(new_n1296));
  INV_X1    g1096(.A(G384), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1291), .A2(G384), .A3(new_n1266), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT125), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1286), .B1(new_n1295), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1286), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(KEYINPUT126), .A3(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT126), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1294), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1298), .A2(KEYINPUT125), .A3(new_n1299), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1285), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1305), .B1(new_n1308), .B2(new_n1302), .ZN(new_n1309));
  OAI211_X1 g1109(.A(G378), .B(new_n1242), .C1(new_n1211), .C2(new_n1215), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1210), .A2(new_n1213), .A3(new_n1206), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1217), .B(new_n1241), .C1(new_n1311), .C2(new_n1003), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1270), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1310), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1279), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1304), .A2(new_n1309), .A3(new_n1315), .ZN(new_n1316));
  XOR2_X1   g1116(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1317));
  NAND2_X1  g1117(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1314), .A2(new_n1279), .A3(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(KEYINPUT62), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1314), .A2(new_n1321), .A3(new_n1279), .A4(new_n1318), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1316), .A2(new_n1317), .A3(new_n1320), .A4(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(G393), .A2(G396), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1271), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1269), .A2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(G390), .A2(new_n1271), .A3(new_n1324), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(G387), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1268), .A2(new_n1327), .A3(new_n1326), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1323), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT61), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1329), .A2(new_n1330), .A3(new_n1333), .ZN(new_n1334));
  AND2_X1   g1134(.A1(new_n1319), .A2(KEYINPUT63), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1319), .A2(KEYINPUT63), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1334), .B(new_n1316), .C1(new_n1335), .C2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1332), .A2(new_n1337), .ZN(G405));
  NAND2_X1  g1138(.A1(G375), .A2(new_n1270), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1339), .B(new_n1310), .C1(new_n1293), .C2(new_n1292), .ZN(new_n1340));
  AOI21_X1  g1140(.A(G378), .B1(new_n1216), .B2(new_n1242), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1310), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1318), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1340), .A2(new_n1331), .A3(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1331), .B1(new_n1340), .B2(new_n1343), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1344), .A2(new_n1345), .ZN(G402));
endmodule


