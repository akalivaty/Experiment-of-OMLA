//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n546, new_n548, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G137), .ZN(new_n465));
  NAND2_X1  g040(.A1(G101), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n464), .A2(new_n467), .ZN(G160));
  NAND2_X1  g043(.A1(new_n461), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G124), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n473), .A2(new_n475), .A3(new_n460), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n471), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  NOR2_X1   g056(.A1(new_n472), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G102), .ZN(new_n483));
  NAND2_X1  g058(.A1(G114), .A2(G2104), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(new_n461), .B2(G126), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n483), .B1(new_n486), .B2(new_n460), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT67), .B(KEYINPUT4), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n476), .A2(KEYINPUT68), .A3(G138), .A4(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n473), .A2(new_n475), .A3(G138), .A4(new_n460), .ZN(new_n491));
  AND2_X1   g066(.A1(KEYINPUT67), .A2(KEYINPUT4), .ZN(new_n492));
  NOR2_X1   g067(.A1(KEYINPUT67), .A2(KEYINPUT4), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n490), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n491), .A2(KEYINPUT66), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n461), .A2(new_n498), .A3(G138), .A4(new_n460), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT4), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n487), .B1(new_n496), .B2(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(KEYINPUT69), .A2(G651), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n502), .B(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(G62), .A3(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n504), .A2(new_n512), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n507), .A2(new_n516), .ZN(G166));
  NOR2_X1   g092(.A1(new_n502), .A2(new_n503), .ZN(new_n518));
  AOI21_X1  g093(.A(KEYINPUT6), .B1(KEYINPUT69), .B2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n520), .A2(new_n506), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n520), .A2(new_n511), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n522), .A2(new_n524), .A3(new_n525), .A4(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n511), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n521), .A2(G52), .B1(new_n532), .B2(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n523), .A2(G90), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  NAND2_X1  g111(.A1(new_n523), .A2(G81), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n521), .A2(G43), .ZN(new_n538));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n511), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n537), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(G176));
  XOR2_X1   g122(.A(KEYINPUT70), .B(KEYINPUT8), .Z(new_n548));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n546), .A2(new_n550), .ZN(G188));
  NAND3_X1  g126(.A1(new_n504), .A2(new_n512), .A3(G91), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n508), .A2(new_n510), .A3(G65), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(G651), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(KEYINPUT71), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n504), .A2(KEYINPUT9), .A3(G543), .A4(new_n559), .ZN(new_n560));
  OAI211_X1 g135(.A(G543), .B(new_n559), .C1(new_n518), .C2(new_n519), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT72), .B1(new_n557), .B2(new_n564), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G299));
  XNOR2_X1  g145(.A(G166), .B(KEYINPUT73), .ZN(G303));
  NAND2_X1  g146(.A1(new_n521), .A2(G49), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n523), .A2(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  AOI22_X1  g150(.A1(G48), .A2(new_n521), .B1(new_n523), .B2(G86), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n511), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT74), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n579), .A2(new_n582), .A3(G651), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n576), .A2(new_n581), .A3(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(G72), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G60), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n511), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(KEYINPUT75), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(KEYINPUT75), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n588), .A2(G651), .A3(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(G47), .A2(new_n521), .B1(new_n523), .B2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n511), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n521), .A2(G54), .B1(new_n596), .B2(G651), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT10), .B1(new_n514), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n523), .A2(new_n600), .A3(G92), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n597), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT76), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n593), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n593), .B1(new_n606), .B2(G868), .ZN(G321));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NOR2_X1   g184(.A1(G286), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n569), .B2(new_n609), .ZN(G297));
  XNOR2_X1  g186(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n543), .A2(new_n609), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n605), .A2(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n609), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n461), .A2(new_n482), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n476), .A2(G135), .ZN(new_n623));
  INV_X1    g198(.A(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(new_n460), .B2(G111), .ZN(new_n626));
  OAI221_X1 g201(.A(new_n623), .B1(new_n624), .B2(new_n469), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G2096), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n622), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2435), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2438), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT14), .ZN(new_n635));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  OR3_X1    g218(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n643), .B1(new_n640), .B2(new_n641), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT79), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT79), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n644), .A2(new_n648), .A3(G14), .A4(new_n645), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(G401));
  XNOR2_X1  g226(.A(G2072), .B(G2078), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT17), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n656), .B1(new_n654), .B2(new_n652), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT81), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n653), .A2(new_n654), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n655), .A2(new_n654), .A3(new_n652), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT80), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n628), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(G2100), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT20), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  INV_X1    g251(.A(new_n673), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n676), .B1(new_n670), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n670), .A2(KEYINPUT82), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT83), .B(G1981), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1986), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n685), .B(new_n687), .Z(G229));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G32), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n470), .A2(G129), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n692));
  NAND3_X1  g267(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n482), .A2(G105), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT90), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n476), .A2(G141), .ZN(new_n698));
  AND4_X1   g273(.A1(new_n691), .A2(new_n694), .A3(new_n697), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT92), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n690), .B1(new_n701), .B2(new_n689), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT27), .B(G1996), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT93), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G1966), .ZN(new_n706));
  NAND2_X1  g281(.A1(G168), .A2(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G16), .B2(G21), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n705), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(G164), .A2(new_n689), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G27), .B2(new_n689), .ZN(new_n711));
  INV_X1    g286(.A(G2078), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n708), .A2(new_n706), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n476), .A2(G140), .ZN(new_n715));
  INV_X1    g290(.A(G128), .ZN(new_n716));
  NOR2_X1   g291(.A1(G104), .A2(G2105), .ZN(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(new_n460), .B2(G116), .ZN(new_n718));
  OAI221_X1 g293(.A(new_n715), .B1(new_n716), .B2(new_n469), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n689), .A2(G26), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT86), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT87), .B(G2067), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n544), .A2(G16), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G16), .B2(G19), .ZN(new_n728));
  INV_X1    g303(.A(G1341), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n713), .A2(new_n714), .A3(new_n726), .A4(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n709), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n461), .A2(G127), .ZN(new_n733));
  NAND2_X1  g308(.A1(G115), .A2(G2104), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n460), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT89), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n476), .A2(G139), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n482), .A2(G103), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n736), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  MUX2_X1   g316(.A(G33), .B(new_n741), .S(G29), .Z(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(G2072), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n732), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n605), .A2(G16), .ZN(new_n746));
  INV_X1    g321(.A(G1348), .ZN(new_n747));
  INV_X1    g322(.A(G4), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n746), .B(new_n747), .C1(new_n748), .C2(G16), .ZN(new_n749));
  INV_X1    g324(.A(G16), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n750), .A2(KEYINPUT23), .A3(G20), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT23), .ZN(new_n752));
  INV_X1    g327(.A(G20), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G16), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n751), .B(new_n754), .C1(new_n569), .C2(new_n750), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G1956), .Z(new_n756));
  NAND2_X1  g331(.A1(G171), .A2(G16), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G5), .B2(G16), .ZN(new_n758));
  INV_X1    g333(.A(G1961), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n711), .A2(new_n712), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n749), .A2(new_n756), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n758), .A2(new_n759), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n728), .A2(new_n729), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n746), .B1(new_n748), .B2(G16), .ZN(new_n766));
  AOI211_X1 g341(.A(new_n764), .B(new_n765), .C1(new_n766), .C2(G1348), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n689), .A2(G35), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G162), .B2(new_n689), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT29), .B(G2090), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n745), .A2(new_n763), .A3(new_n767), .A4(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT85), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(KEYINPUT36), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n750), .A2(G6), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G305), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT84), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT32), .B(G1981), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G16), .A2(G23), .ZN(new_n780));
  INV_X1    g355(.A(G288), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(G16), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT33), .B(G1976), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n750), .A2(G22), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G166), .B2(new_n750), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1971), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n779), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT34), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n779), .A2(KEYINPUT34), .A3(new_n788), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n689), .A2(G25), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n470), .A2(G119), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n476), .A2(G131), .ZN(new_n796));
  OR2_X1    g371(.A1(G95), .A2(G2105), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n797), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n795), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n794), .B1(new_n800), .B2(new_n689), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT35), .B(G1991), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G1986), .ZN(new_n804));
  INV_X1    g379(.A(G290), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(new_n750), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n750), .B2(G24), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n803), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n804), .B2(new_n807), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n774), .B1(new_n793), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n793), .A2(new_n774), .A3(new_n809), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n772), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT31), .B(G11), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT94), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT30), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n689), .B1(new_n816), .B2(G28), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(KEYINPUT95), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(G28), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(KEYINPUT95), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n815), .B(new_n821), .C1(new_n627), .C2(new_n689), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT96), .Z(new_n823));
  OR2_X1    g398(.A1(KEYINPUT24), .A2(G34), .ZN(new_n824));
  NAND2_X1  g399(.A1(KEYINPUT24), .A2(G34), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n824), .A2(new_n689), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G160), .B2(new_n689), .ZN(new_n827));
  INV_X1    g402(.A(G2084), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n702), .A2(new_n704), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n813), .A2(new_n823), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(G311));
  INV_X1    g407(.A(KEYINPUT97), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n765), .B1(new_n766), .B2(G1348), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n835), .B(new_n771), .C1(new_n759), .C2(new_n758), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n836), .A2(new_n744), .A3(new_n762), .ZN(new_n837));
  INV_X1    g412(.A(new_n812), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n837), .B(new_n830), .C1(new_n838), .C2(new_n810), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n840), .A2(KEYINPUT97), .A3(new_n823), .A4(new_n829), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n834), .A2(new_n841), .ZN(G150));
  NAND2_X1  g417(.A1(G80), .A2(G543), .ZN(new_n843));
  INV_X1    g418(.A(G67), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n511), .B2(new_n844), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n521), .A2(G55), .B1(new_n845), .B2(G651), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT99), .B(G93), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n523), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT101), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n606), .A2(G559), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n544), .A2(new_n849), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n543), .A2(new_n846), .A3(new_n848), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n855), .B(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT100), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(G860), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n852), .B1(new_n862), .B2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(new_n480), .B(KEYINPUT102), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G160), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n627), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n473), .A2(new_n475), .A3(G126), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n460), .B1(new_n869), .B2(new_n484), .ZN(new_n870));
  INV_X1    g445(.A(new_n483), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT103), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n873), .B(new_n483), .C1(new_n486), .C2(new_n460), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  AND4_X1   g450(.A1(G138), .A2(new_n473), .A3(new_n475), .A4(new_n460), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT68), .B1(new_n876), .B2(new_n488), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n491), .A2(new_n490), .A3(new_n494), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n500), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n799), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n868), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n741), .A2(new_n699), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n701), .B2(new_n741), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n868), .A2(new_n881), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n884), .B1(new_n882), .B2(new_n885), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n476), .A2(G142), .ZN(new_n888));
  INV_X1    g463(.A(G130), .ZN(new_n889));
  NOR2_X1   g464(.A1(G106), .A2(G2105), .ZN(new_n890));
  OAI21_X1  g465(.A(G2104), .B1(new_n460), .B2(G118), .ZN(new_n891));
  OAI221_X1 g466(.A(new_n888), .B1(new_n889), .B2(new_n469), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n620), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n719), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  OR3_X1    g470(.A1(new_n886), .A2(new_n887), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n895), .B1(new_n886), .B2(new_n887), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g475(.A1(new_n805), .A2(G288), .ZN(new_n901));
  NAND2_X1  g476(.A1(G290), .A2(new_n781), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT108), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(KEYINPUT108), .A3(new_n902), .ZN(new_n905));
  XNOR2_X1  g480(.A(G305), .B(G166), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n903), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(KEYINPUT110), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n907), .A2(new_n909), .A3(KEYINPUT109), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n912), .B1(new_n918), .B2(new_n911), .ZN(new_n919));
  INV_X1    g494(.A(new_n602), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n567), .A2(new_n920), .A3(new_n568), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT104), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n567), .A2(new_n920), .A3(new_n923), .A4(new_n568), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT106), .B1(new_n569), .B2(new_n602), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n569), .A2(KEYINPUT106), .A3(new_n602), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT107), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT105), .B1(new_n922), .B2(new_n924), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n569), .A2(new_n602), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n922), .A2(KEYINPUT105), .A3(new_n924), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n932), .A2(KEYINPUT41), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n934), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n937), .A2(new_n931), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n938), .A2(KEYINPUT107), .A3(KEYINPUT41), .A4(new_n933), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n616), .B(new_n858), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n919), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n919), .B1(new_n945), .B2(new_n942), .ZN(new_n947));
  OAI21_X1  g522(.A(G868), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n849), .A2(new_n609), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(G295));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n949), .ZN(G331));
  NAND2_X1  g526(.A1(G168), .A2(G301), .ZN(new_n952));
  NAND2_X1  g527(.A1(G171), .A2(G286), .ZN(new_n953));
  AND4_X1   g528(.A1(new_n856), .A2(new_n952), .A3(new_n953), .A4(new_n857), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n952), .A2(new_n953), .B1(new_n856), .B2(new_n857), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n936), .A2(new_n939), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT111), .B1(new_n954), .B2(new_n955), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n955), .A2(KEYINPUT111), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n943), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n916), .A2(new_n957), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n914), .A2(new_n915), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n928), .A2(KEYINPUT41), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n960), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n943), .B1(new_n965), .B2(new_n956), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n929), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n962), .A2(new_n968), .A3(new_n897), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n957), .A2(new_n961), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n963), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n972), .A2(new_n897), .A3(new_n962), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT43), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n972), .A2(new_n974), .A3(new_n897), .A4(new_n962), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n979), .A3(KEYINPUT44), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n977), .B1(new_n982), .B2(new_n983), .ZN(G397));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n872), .A2(new_n874), .B1(new_n496), .B2(new_n500), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n985), .B1(new_n986), .B2(G1384), .ZN(new_n987));
  NAND2_X1  g562(.A1(G160), .A2(G40), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  XOR2_X1   g565(.A(new_n719), .B(G2067), .Z(new_n991));
  AOI21_X1  g566(.A(new_n990), .B1(new_n699), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1996), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n989), .A2(KEYINPUT46), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT46), .B1(new_n989), .B2(new_n993), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT47), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n989), .A2(new_n804), .A3(new_n805), .ZN(new_n998));
  XOR2_X1   g573(.A(new_n998), .B(KEYINPUT48), .Z(new_n999));
  NAND2_X1  g574(.A1(new_n701), .A2(new_n993), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n1000), .B(new_n991), .C1(new_n993), .C2(new_n699), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n799), .B(new_n802), .Z(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n999), .B1(new_n1004), .B2(new_n989), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n800), .A2(new_n802), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n719), .A2(G2067), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n990), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n997), .A2(new_n1005), .A3(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(G305), .A2(G1981), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n576), .A2(new_n580), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(G1981), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT49), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1384), .B1(new_n875), .B2(new_n879), .ZN(new_n1017));
  INV_X1    g592(.A(new_n988), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1976), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1019), .B1(new_n1021), .B2(G288), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT52), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  AOI211_X1 g599(.A(KEYINPUT52), .B(new_n1022), .C1(new_n1021), .C2(G288), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G303), .A2(G8), .ZN(new_n1027));
  XOR2_X1   g602(.A(new_n1027), .B(KEYINPUT55), .Z(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  INV_X1    g604(.A(G1384), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n880), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n1018), .A3(new_n1032), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1033), .A2(G2090), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1017), .A2(KEYINPUT45), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n985), .B1(G164), .B2(G1384), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n1018), .ZN(new_n1037));
  INV_X1    g612(.A(G1971), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1016), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1028), .A2(new_n1040), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n1028), .A2(new_n1040), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1026), .A2(KEYINPUT63), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1031), .A2(new_n1032), .A3(new_n828), .A4(new_n1018), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1018), .B1(new_n1017), .B2(KEYINPUT45), .ZN(new_n1047));
  NOR3_X1   g622(.A1(G164), .A2(new_n985), .A3(G1384), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n706), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n988), .B1(new_n1017), .B2(new_n1029), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1050), .A2(KEYINPUT113), .A3(new_n828), .A4(new_n1032), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1046), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(G8), .A3(G168), .ZN(new_n1053));
  XOR2_X1   g628(.A(new_n1053), .B(KEYINPUT114), .Z(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT63), .B1(new_n1043), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1041), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1026), .A2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g632(.A(G1976), .B(G288), .C1(new_n1015), .C2(new_n1019), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1011), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1019), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1055), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1052), .A2(G8), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1062), .B1(new_n1063), .B2(KEYINPUT122), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1052), .A2(G286), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1046), .A2(new_n1049), .A3(new_n1051), .A4(G168), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(G8), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1069), .B1(new_n1052), .B2(G8), .ZN(new_n1070));
  OAI211_X1 g645(.A(G8), .B(new_n1066), .C1(new_n1070), .C2(new_n1062), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT62), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT125), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1068), .A2(new_n1075), .A3(new_n1071), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n987), .A2(KEYINPUT53), .A3(new_n712), .A4(new_n1018), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1077), .A2(new_n1048), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1035), .A2(new_n712), .A3(new_n1036), .A4(new_n1018), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1079), .A2(new_n1080), .B1(new_n1033), .B2(new_n759), .ZN(new_n1081));
  AOI21_X1  g656(.A(G301), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1076), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1072), .A2(new_n1084), .A3(KEYINPUT62), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1074), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1035), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1077), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1077), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1081), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1087), .B1(new_n1093), .B2(G171), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1078), .A2(new_n1081), .A3(G301), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT124), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1077), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(KEYINPUT123), .A3(new_n1035), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n1090), .ZN(new_n1100));
  AOI21_X1  g675(.A(G301), .B1(new_n1100), .B2(new_n1081), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n1102));
  NOR4_X1   g677(.A1(new_n1101), .A2(new_n1102), .A3(new_n1095), .A4(new_n1087), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1097), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT56), .B(G2072), .ZN(new_n1105));
  AND4_X1   g680(.A1(new_n1036), .A2(new_n1035), .A3(new_n1018), .A4(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT115), .B(G1956), .ZN(new_n1107));
  NOR2_X1   g682(.A1(G164), .A2(G1384), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n988), .B1(new_n1108), .B2(new_n1029), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT50), .B1(new_n986), .B2(G1384), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1107), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G91), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n520), .A2(new_n1113), .A3(new_n511), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n556), .B1(new_n553), .B2(new_n554), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT117), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n560), .A2(new_n563), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n552), .B(new_n1118), .C1(new_n555), .C2(new_n556), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1116), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(KEYINPUT116), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT116), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n565), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1122), .B1(new_n1124), .B2(new_n1121), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT118), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(new_n1122), .C1(new_n1124), .C2(new_n1121), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1112), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1126), .B(new_n1128), .C1(new_n1106), .C2(new_n1111), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1348), .B1(new_n1050), .B2(new_n1032), .ZN(new_n1135));
  INV_X1    g710(.A(new_n603), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(G2067), .ZN(new_n1138));
  NOR4_X1   g713(.A1(new_n1135), .A2(new_n1136), .A3(new_n1138), .A4(KEYINPUT60), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1033), .A2(new_n747), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1140), .B(new_n1136), .C1(G2067), .C2(new_n1137), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n603), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1139), .B1(new_n1143), .B2(KEYINPUT60), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1035), .A2(new_n993), .A3(new_n1036), .A4(new_n1018), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT121), .B(G1341), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT58), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1137), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n543), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(new_n1149), .B(KEYINPUT59), .Z(new_n1150));
  NAND3_X1  g725(.A1(new_n1130), .A2(KEYINPUT61), .A3(new_n1131), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1134), .A2(new_n1144), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1142), .A2(KEYINPUT119), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1154), .B(new_n603), .C1(new_n1135), .C2(new_n1138), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1153), .A2(new_n1131), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1130), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(KEYINPUT120), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1156), .A2(new_n1159), .A3(new_n1130), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1152), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1093), .A2(G171), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1087), .B1(new_n1162), .B2(new_n1082), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1104), .A2(new_n1161), .A3(new_n1163), .A4(new_n1072), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1054), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1043), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1086), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1039), .B1(G2090), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1028), .B1(G8), .B2(new_n1169), .ZN(new_n1170));
  NOR4_X1   g745(.A1(new_n1170), .A2(new_n1056), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1061), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(G290), .B(new_n804), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n990), .B1(new_n1003), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1010), .B1(new_n1172), .B2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g750(.A(G229), .ZN(new_n1177));
  NAND3_X1  g751(.A1(new_n650), .A2(G319), .A3(new_n667), .ZN(new_n1178));
  XNOR2_X1  g752(.A(new_n1178), .B(KEYINPUT126), .ZN(new_n1179));
  NAND4_X1  g753(.A1(new_n975), .A2(new_n1177), .A3(new_n899), .A4(new_n1179), .ZN(G225));
  INV_X1    g754(.A(G225), .ZN(G308));
endmodule


