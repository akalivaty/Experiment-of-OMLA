

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U550 ( .A(n870), .Z(n516) );
  XNOR2_X1 U551 ( .A(KEYINPUT17), .B(n518), .ZN(n870) );
  XNOR2_X1 U552 ( .A(n585), .B(n584), .ZN(n606) );
  NAND2_X1 U553 ( .A1(n658), .A2(n657), .ZN(n660) );
  INV_X1 U554 ( .A(KEYINPUT29), .ZN(n659) );
  XNOR2_X1 U555 ( .A(n660), .B(n659), .ZN(n661) );
  INV_X1 U556 ( .A(KEYINPUT84), .ZN(n584) );
  NOR2_X1 U557 ( .A1(G651), .A2(n562), .ZN(n790) );
  INV_X1 U558 ( .A(G2105), .ZN(n521) );
  AND2_X1 U559 ( .A1(n521), .A2(G2104), .ZN(n869) );
  NAND2_X1 U560 ( .A1(n869), .A2(G102), .ZN(n520) );
  NOR2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  XOR2_X1 U562 ( .A(KEYINPUT66), .B(n517), .Z(n518) );
  NAND2_X1 U563 ( .A1(G138), .A2(n516), .ZN(n519) );
  NAND2_X1 U564 ( .A1(n520), .A2(n519), .ZN(n525) );
  NOR2_X1 U565 ( .A1(G2104), .A2(n521), .ZN(n873) );
  NAND2_X1 U566 ( .A1(G126), .A2(n873), .ZN(n523) );
  AND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n875) );
  NAND2_X1 U568 ( .A1(G114), .A2(n875), .ZN(n522) );
  NAND2_X1 U569 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U570 ( .A1(n525), .A2(n524), .ZN(G164) );
  INV_X1 U571 ( .A(G651), .ZN(n528) );
  NOR2_X1 U572 ( .A1(G543), .A2(n528), .ZN(n526) );
  XOR2_X1 U573 ( .A(KEYINPUT68), .B(n526), .Z(n527) );
  XNOR2_X1 U574 ( .A(KEYINPUT1), .B(n527), .ZN(n786) );
  AND2_X1 U575 ( .A1(G60), .A2(n786), .ZN(n533) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n562) );
  NOR2_X1 U577 ( .A1(n562), .A2(n528), .ZN(n782) );
  NAND2_X1 U578 ( .A1(n782), .A2(G72), .ZN(n531) );
  NOR2_X1 U579 ( .A1(G543), .A2(G651), .ZN(n529) );
  XNOR2_X1 U580 ( .A(n529), .B(KEYINPUT64), .ZN(n783) );
  NAND2_X1 U581 ( .A1(G85), .A2(n783), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U583 ( .A1(n533), .A2(n532), .ZN(n535) );
  NAND2_X1 U584 ( .A1(n790), .A2(G47), .ZN(n534) );
  NAND2_X1 U585 ( .A1(n535), .A2(n534), .ZN(G290) );
  NAND2_X1 U586 ( .A1(G89), .A2(n783), .ZN(n536) );
  XNOR2_X1 U587 ( .A(n536), .B(KEYINPUT4), .ZN(n538) );
  NAND2_X1 U588 ( .A1(G76), .A2(n782), .ZN(n537) );
  NAND2_X1 U589 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U590 ( .A(n539), .B(KEYINPUT5), .ZN(n545) );
  XNOR2_X1 U591 ( .A(KEYINPUT73), .B(KEYINPUT6), .ZN(n543) );
  NAND2_X1 U592 ( .A1(n790), .A2(G51), .ZN(n541) );
  NAND2_X1 U593 ( .A1(G63), .A2(n786), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U595 ( .A(n543), .B(n542), .ZN(n544) );
  NAND2_X1 U596 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U597 ( .A(KEYINPUT7), .B(n546), .ZN(G168) );
  XOR2_X1 U598 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U599 ( .A1(n790), .A2(G52), .ZN(n548) );
  NAND2_X1 U600 ( .A1(G64), .A2(n786), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n548), .A2(n547), .ZN(n554) );
  NAND2_X1 U602 ( .A1(G90), .A2(n783), .ZN(n549) );
  XOR2_X1 U603 ( .A(KEYINPUT69), .B(n549), .Z(n551) );
  NAND2_X1 U604 ( .A1(n782), .A2(G77), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U606 ( .A(KEYINPUT9), .B(n552), .Z(n553) );
  NOR2_X1 U607 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U608 ( .A(KEYINPUT70), .B(n555), .ZN(G171) );
  INV_X1 U609 ( .A(G171), .ZN(G301) );
  NAND2_X1 U610 ( .A1(n782), .A2(G75), .ZN(n557) );
  NAND2_X1 U611 ( .A1(G88), .A2(n783), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U613 ( .A1(n790), .A2(G50), .ZN(n559) );
  NAND2_X1 U614 ( .A1(G62), .A2(n786), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U616 ( .A1(n561), .A2(n560), .ZN(G166) );
  NAND2_X1 U617 ( .A1(G87), .A2(n562), .ZN(n564) );
  NAND2_X1 U618 ( .A1(G74), .A2(G651), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U620 ( .A1(n786), .A2(n565), .ZN(n567) );
  NAND2_X1 U621 ( .A1(n790), .A2(G49), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n567), .A2(n566), .ZN(G288) );
  INV_X1 U623 ( .A(G166), .ZN(G303) );
  NAND2_X1 U624 ( .A1(G73), .A2(n782), .ZN(n568) );
  XOR2_X1 U625 ( .A(KEYINPUT2), .B(n568), .Z(n573) );
  NAND2_X1 U626 ( .A1(G61), .A2(n786), .ZN(n570) );
  NAND2_X1 U627 ( .A1(G86), .A2(n783), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U629 ( .A(KEYINPUT81), .B(n571), .Z(n572) );
  NOR2_X1 U630 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U631 ( .A1(n790), .A2(G48), .ZN(n574) );
  NAND2_X1 U632 ( .A1(n575), .A2(n574), .ZN(G305) );
  NOR2_X1 U633 ( .A1(G164), .A2(G1384), .ZN(n607) );
  NAND2_X1 U634 ( .A1(G125), .A2(n873), .ZN(n581) );
  NAND2_X1 U635 ( .A1(G137), .A2(n870), .ZN(n578) );
  NAND2_X1 U636 ( .A1(n875), .A2(G113), .ZN(n576) );
  XOR2_X1 U637 ( .A(KEYINPUT65), .B(n576), .Z(n577) );
  NAND2_X1 U638 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U639 ( .A(n579), .B(KEYINPUT67), .ZN(n580) );
  AND2_X1 U640 ( .A1(n581), .A2(n580), .ZN(n753) );
  NAND2_X1 U641 ( .A1(G101), .A2(n869), .ZN(n582) );
  XOR2_X1 U642 ( .A(KEYINPUT23), .B(n582), .Z(n752) );
  AND2_X1 U643 ( .A1(G40), .A2(n752), .ZN(n583) );
  NAND2_X1 U644 ( .A1(n753), .A2(n583), .ZN(n585) );
  INV_X1 U645 ( .A(n606), .ZN(n586) );
  NOR2_X1 U646 ( .A1(n607), .A2(n586), .ZN(n748) );
  NAND2_X1 U647 ( .A1(n873), .A2(G129), .ZN(n588) );
  NAND2_X1 U648 ( .A1(G141), .A2(n516), .ZN(n587) );
  NAND2_X1 U649 ( .A1(n588), .A2(n587), .ZN(n593) );
  XOR2_X1 U650 ( .A(KEYINPUT38), .B(KEYINPUT90), .Z(n590) );
  NAND2_X1 U651 ( .A1(G105), .A2(n869), .ZN(n589) );
  XNOR2_X1 U652 ( .A(n590), .B(n589), .ZN(n591) );
  XOR2_X1 U653 ( .A(KEYINPUT89), .B(n591), .Z(n592) );
  NOR2_X1 U654 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U655 ( .A1(n875), .A2(G117), .ZN(n594) );
  NAND2_X1 U656 ( .A1(n595), .A2(n594), .ZN(n881) );
  NAND2_X1 U657 ( .A1(G1996), .A2(n881), .ZN(n604) );
  NAND2_X1 U658 ( .A1(G119), .A2(n873), .ZN(n597) );
  NAND2_X1 U659 ( .A1(G107), .A2(n875), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U661 ( .A1(n516), .A2(G131), .ZN(n598) );
  XOR2_X1 U662 ( .A(KEYINPUT88), .B(n598), .Z(n599) );
  NOR2_X1 U663 ( .A1(n600), .A2(n599), .ZN(n602) );
  NAND2_X1 U664 ( .A1(n869), .A2(G95), .ZN(n601) );
  NAND2_X1 U665 ( .A1(n602), .A2(n601), .ZN(n886) );
  NAND2_X1 U666 ( .A1(G1991), .A2(n886), .ZN(n603) );
  NAND2_X1 U667 ( .A1(n604), .A2(n603), .ZN(n972) );
  NAND2_X1 U668 ( .A1(n748), .A2(n972), .ZN(n736) );
  XNOR2_X1 U669 ( .A(G1986), .B(G290), .ZN(n1006) );
  NAND2_X1 U670 ( .A1(n748), .A2(n1006), .ZN(n605) );
  NAND2_X1 U671 ( .A1(n736), .A2(n605), .ZN(n721) );
  XOR2_X1 U672 ( .A(KEYINPUT25), .B(G2078), .Z(n918) );
  NAND2_X1 U673 ( .A1(n607), .A2(n606), .ZN(n674) );
  NOR2_X1 U674 ( .A1(n918), .A2(n674), .ZN(n609) );
  INV_X1 U675 ( .A(n674), .ZN(n646) );
  NOR2_X1 U676 ( .A1(n646), .A2(G1961), .ZN(n608) );
  NOR2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U678 ( .A(KEYINPUT92), .B(n610), .ZN(n668) );
  NOR2_X1 U679 ( .A1(G301), .A2(n668), .ZN(n611) );
  XNOR2_X1 U680 ( .A(n611), .B(KEYINPUT93), .ZN(n662) );
  NAND2_X1 U681 ( .A1(n646), .A2(G2072), .ZN(n612) );
  XNOR2_X1 U682 ( .A(KEYINPUT27), .B(n612), .ZN(n615) );
  NAND2_X1 U683 ( .A1(G1956), .A2(n674), .ZN(n613) );
  XOR2_X1 U684 ( .A(n613), .B(KEYINPUT94), .Z(n614) );
  NOR2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n654) );
  NAND2_X1 U686 ( .A1(n790), .A2(G53), .ZN(n617) );
  NAND2_X1 U687 ( .A1(G65), .A2(n786), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U689 ( .A1(n782), .A2(G78), .ZN(n619) );
  NAND2_X1 U690 ( .A1(G91), .A2(n783), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U692 ( .A1(n621), .A2(n620), .ZN(n996) );
  NOR2_X1 U693 ( .A1(n654), .A2(n996), .ZN(n623) );
  XNOR2_X1 U694 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n623), .B(n622), .ZN(n658) );
  INV_X1 U696 ( .A(G1996), .ZN(n624) );
  NOR2_X1 U697 ( .A1(n674), .A2(n624), .ZN(n625) );
  XNOR2_X1 U698 ( .A(n625), .B(KEYINPUT26), .ZN(n637) );
  NAND2_X1 U699 ( .A1(n674), .A2(G1341), .ZN(n635) );
  NAND2_X1 U700 ( .A1(n786), .A2(G56), .ZN(n626) );
  XOR2_X1 U701 ( .A(KEYINPUT14), .B(n626), .Z(n632) );
  NAND2_X1 U702 ( .A1(G81), .A2(n783), .ZN(n627) );
  XNOR2_X1 U703 ( .A(n627), .B(KEYINPUT12), .ZN(n629) );
  NAND2_X1 U704 ( .A1(G68), .A2(n782), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U706 ( .A(KEYINPUT13), .B(n630), .Z(n631) );
  NOR2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n790), .A2(G43), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n1014) );
  INV_X1 U710 ( .A(n1014), .ZN(n756) );
  NAND2_X1 U711 ( .A1(n635), .A2(n756), .ZN(n636) );
  NOR2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n650) );
  NAND2_X1 U713 ( .A1(n790), .A2(G54), .ZN(n644) );
  NAND2_X1 U714 ( .A1(n782), .A2(G79), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G66), .A2(n786), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n783), .A2(G92), .ZN(n640) );
  XOR2_X1 U718 ( .A(KEYINPUT72), .B(n640), .Z(n641) );
  NOR2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U721 ( .A(KEYINPUT15), .B(n645), .Z(n999) );
  NAND2_X1 U722 ( .A1(G1348), .A2(n674), .ZN(n648) );
  NAND2_X1 U723 ( .A1(G2067), .A2(n646), .ZN(n647) );
  NAND2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n651) );
  NOR2_X1 U725 ( .A1(n999), .A2(n651), .ZN(n649) );
  OR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U727 ( .A1(n999), .A2(n651), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U729 ( .A1(n996), .A2(n654), .ZN(n655) );
  NAND2_X1 U730 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n673) );
  NOR2_X1 U732 ( .A1(G2084), .A2(n674), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(KEYINPUT91), .ZN(n684) );
  NAND2_X1 U734 ( .A1(G8), .A2(n684), .ZN(n664) );
  NAND2_X1 U735 ( .A1(G8), .A2(n674), .ZN(n715) );
  NOR2_X1 U736 ( .A1(G1966), .A2(n715), .ZN(n688) );
  NOR2_X1 U737 ( .A1(n664), .A2(n688), .ZN(n666) );
  XOR2_X1 U738 ( .A(KEYINPUT30), .B(KEYINPUT96), .Z(n665) );
  XNOR2_X1 U739 ( .A(n666), .B(n665), .ZN(n667) );
  NOR2_X1 U740 ( .A1(n667), .A2(G168), .ZN(n670) );
  AND2_X1 U741 ( .A1(n668), .A2(G301), .ZN(n669) );
  NOR2_X1 U742 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U743 ( .A(KEYINPUT31), .B(n671), .Z(n672) );
  NAND2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n686) );
  NAND2_X1 U745 ( .A1(G286), .A2(n686), .ZN(n681) );
  NOR2_X1 U746 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U747 ( .A(KEYINPUT97), .B(n675), .ZN(n678) );
  NOR2_X1 U748 ( .A1(G1971), .A2(n715), .ZN(n676) );
  NOR2_X1 U749 ( .A1(G166), .A2(n676), .ZN(n677) );
  NAND2_X1 U750 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U751 ( .A(n679), .B(KEYINPUT98), .ZN(n680) );
  NAND2_X1 U752 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U753 ( .A1(n682), .A2(G8), .ZN(n683) );
  XNOR2_X1 U754 ( .A(n683), .B(KEYINPUT32), .ZN(n692) );
  INV_X1 U755 ( .A(n684), .ZN(n685) );
  NAND2_X1 U756 ( .A1(G8), .A2(n685), .ZN(n690) );
  INV_X1 U757 ( .A(n686), .ZN(n687) );
  NOR2_X1 U758 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n711) );
  NOR2_X1 U761 ( .A1(G1976), .A2(G288), .ZN(n700) );
  NOR2_X1 U762 ( .A1(G1971), .A2(G303), .ZN(n693) );
  NOR2_X1 U763 ( .A1(n700), .A2(n693), .ZN(n997) );
  INV_X1 U764 ( .A(KEYINPUT33), .ZN(n694) );
  AND2_X1 U765 ( .A1(n997), .A2(n694), .ZN(n695) );
  NAND2_X1 U766 ( .A1(n711), .A2(n695), .ZN(n699) );
  NAND2_X1 U767 ( .A1(G1976), .A2(G288), .ZN(n1004) );
  INV_X1 U768 ( .A(n1004), .ZN(n696) );
  NOR2_X1 U769 ( .A1(n696), .A2(n715), .ZN(n697) );
  OR2_X1 U770 ( .A1(KEYINPUT33), .A2(n697), .ZN(n698) );
  AND2_X1 U771 ( .A1(n699), .A2(n698), .ZN(n708) );
  NAND2_X1 U772 ( .A1(KEYINPUT33), .A2(n700), .ZN(n701) );
  XOR2_X1 U773 ( .A(KEYINPUT99), .B(n701), .Z(n702) );
  NOR2_X1 U774 ( .A1(n715), .A2(n702), .ZN(n703) );
  XNOR2_X1 U775 ( .A(n703), .B(KEYINPUT100), .ZN(n706) );
  XNOR2_X1 U776 ( .A(G1981), .B(KEYINPUT101), .ZN(n704) );
  XNOR2_X1 U777 ( .A(n704), .B(G305), .ZN(n993) );
  INV_X1 U778 ( .A(n993), .ZN(n705) );
  NOR2_X1 U779 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U780 ( .A1(n708), .A2(n707), .ZN(n719) );
  NOR2_X1 U781 ( .A1(G2090), .A2(G303), .ZN(n709) );
  NAND2_X1 U782 ( .A1(G8), .A2(n709), .ZN(n710) );
  NAND2_X1 U783 ( .A1(n711), .A2(n710), .ZN(n712) );
  AND2_X1 U784 ( .A1(n712), .A2(n715), .ZN(n717) );
  NOR2_X1 U785 ( .A1(G1981), .A2(G305), .ZN(n713) );
  XOR2_X1 U786 ( .A(n713), .B(KEYINPUT24), .Z(n714) );
  NOR2_X1 U787 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U788 ( .A1(n717), .A2(n716), .ZN(n718) );
  AND2_X1 U789 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U790 ( .A1(n721), .A2(n720), .ZN(n734) );
  NAND2_X1 U791 ( .A1(n869), .A2(G104), .ZN(n723) );
  NAND2_X1 U792 ( .A1(G140), .A2(n516), .ZN(n722) );
  NAND2_X1 U793 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U794 ( .A(KEYINPUT34), .B(n724), .ZN(n731) );
  XNOR2_X1 U795 ( .A(KEYINPUT86), .B(KEYINPUT35), .ZN(n729) );
  NAND2_X1 U796 ( .A1(n875), .A2(G116), .ZN(n727) );
  NAND2_X1 U797 ( .A1(n873), .A2(G128), .ZN(n725) );
  XOR2_X1 U798 ( .A(KEYINPUT85), .B(n725), .Z(n726) );
  NAND2_X1 U799 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U800 ( .A(n729), .B(n728), .Z(n730) );
  NOR2_X1 U801 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U802 ( .A(n732), .B(KEYINPUT36), .Z(n733) );
  XNOR2_X1 U803 ( .A(KEYINPUT87), .B(n733), .ZN(n889) );
  XNOR2_X1 U804 ( .A(G2067), .B(KEYINPUT37), .ZN(n745) );
  NOR2_X1 U805 ( .A1(n889), .A2(n745), .ZN(n973) );
  NAND2_X1 U806 ( .A1(n748), .A2(n973), .ZN(n743) );
  NAND2_X1 U807 ( .A1(n734), .A2(n743), .ZN(n735) );
  XNOR2_X1 U808 ( .A(n735), .B(KEYINPUT102), .ZN(n750) );
  XOR2_X1 U809 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n742) );
  NOR2_X1 U810 ( .A1(G1996), .A2(n881), .ZN(n977) );
  INV_X1 U811 ( .A(n736), .ZN(n739) );
  NOR2_X1 U812 ( .A1(G1986), .A2(G290), .ZN(n737) );
  NOR2_X1 U813 ( .A1(G1991), .A2(n886), .ZN(n963) );
  NOR2_X1 U814 ( .A1(n737), .A2(n963), .ZN(n738) );
  NOR2_X1 U815 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U816 ( .A1(n977), .A2(n740), .ZN(n741) );
  XNOR2_X1 U817 ( .A(n742), .B(n741), .ZN(n744) );
  NAND2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n746) );
  NAND2_X1 U819 ( .A1(n889), .A2(n745), .ZN(n966) );
  NAND2_X1 U820 ( .A1(n746), .A2(n966), .ZN(n747) );
  NAND2_X1 U821 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U822 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U823 ( .A(n751), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U824 ( .A1(n753), .A2(n752), .ZN(G160) );
  AND2_X1 U825 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U826 ( .A(G132), .ZN(G219) );
  INV_X1 U827 ( .A(G82), .ZN(G220) );
  NAND2_X1 U828 ( .A1(G7), .A2(G661), .ZN(n754) );
  XNOR2_X1 U829 ( .A(n754), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U830 ( .A(G223), .ZN(n821) );
  NAND2_X1 U831 ( .A1(n821), .A2(G567), .ZN(n755) );
  XOR2_X1 U832 ( .A(KEYINPUT11), .B(n755), .Z(G234) );
  NAND2_X1 U833 ( .A1(n756), .A2(G860), .ZN(G153) );
  NAND2_X1 U834 ( .A1(G301), .A2(G868), .ZN(n758) );
  INV_X1 U835 ( .A(G868), .ZN(n803) );
  NAND2_X1 U836 ( .A1(n999), .A2(n803), .ZN(n757) );
  NAND2_X1 U837 ( .A1(n758), .A2(n757), .ZN(G284) );
  INV_X1 U838 ( .A(n996), .ZN(G299) );
  NOR2_X1 U839 ( .A1(G868), .A2(G299), .ZN(n759) );
  XNOR2_X1 U840 ( .A(n759), .B(KEYINPUT74), .ZN(n761) );
  NOR2_X1 U841 ( .A1(n803), .A2(G286), .ZN(n760) );
  NOR2_X1 U842 ( .A1(n761), .A2(n760), .ZN(G297) );
  INV_X1 U843 ( .A(G559), .ZN(n762) );
  NOR2_X1 U844 ( .A1(G860), .A2(n762), .ZN(n763) );
  XNOR2_X1 U845 ( .A(KEYINPUT75), .B(n763), .ZN(n764) );
  INV_X1 U846 ( .A(n999), .ZN(n780) );
  NAND2_X1 U847 ( .A1(n764), .A2(n780), .ZN(n765) );
  XNOR2_X1 U848 ( .A(n765), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U849 ( .A1(n780), .A2(G868), .ZN(n766) );
  NOR2_X1 U850 ( .A1(G559), .A2(n766), .ZN(n767) );
  XNOR2_X1 U851 ( .A(n767), .B(KEYINPUT76), .ZN(n769) );
  NOR2_X1 U852 ( .A1(n1014), .A2(G868), .ZN(n768) );
  NOR2_X1 U853 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U854 ( .A(KEYINPUT77), .B(n770), .Z(G282) );
  NAND2_X1 U855 ( .A1(n873), .A2(G123), .ZN(n771) );
  XNOR2_X1 U856 ( .A(n771), .B(KEYINPUT18), .ZN(n773) );
  NAND2_X1 U857 ( .A1(G111), .A2(n875), .ZN(n772) );
  NAND2_X1 U858 ( .A1(n773), .A2(n772), .ZN(n777) );
  NAND2_X1 U859 ( .A1(n869), .A2(G99), .ZN(n775) );
  NAND2_X1 U860 ( .A1(G135), .A2(n516), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n962) );
  XOR2_X1 U863 ( .A(G2096), .B(n962), .Z(n778) );
  NOR2_X1 U864 ( .A1(G2100), .A2(n778), .ZN(n779) );
  XOR2_X1 U865 ( .A(KEYINPUT78), .B(n779), .Z(G156) );
  NAND2_X1 U866 ( .A1(n780), .A2(G559), .ZN(n801) );
  XNOR2_X1 U867 ( .A(n1014), .B(n801), .ZN(n781) );
  NOR2_X1 U868 ( .A1(n781), .A2(G860), .ZN(n794) );
  NAND2_X1 U869 ( .A1(n782), .A2(G80), .ZN(n785) );
  NAND2_X1 U870 ( .A1(G93), .A2(n783), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n789) );
  NAND2_X1 U872 ( .A1(G67), .A2(n786), .ZN(n787) );
  XNOR2_X1 U873 ( .A(KEYINPUT79), .B(n787), .ZN(n788) );
  NOR2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U875 ( .A1(n790), .A2(G55), .ZN(n791) );
  NAND2_X1 U876 ( .A1(n792), .A2(n791), .ZN(n804) );
  XOR2_X1 U877 ( .A(n804), .B(KEYINPUT80), .Z(n793) );
  XNOR2_X1 U878 ( .A(n794), .B(n793), .ZN(G145) );
  XNOR2_X1 U879 ( .A(n1014), .B(G305), .ZN(n800) );
  XNOR2_X1 U880 ( .A(G288), .B(KEYINPUT19), .ZN(n796) );
  XNOR2_X1 U881 ( .A(n996), .B(G166), .ZN(n795) );
  XNOR2_X1 U882 ( .A(n796), .B(n795), .ZN(n797) );
  XOR2_X1 U883 ( .A(n797), .B(G290), .Z(n798) );
  XNOR2_X1 U884 ( .A(n804), .B(n798), .ZN(n799) );
  XNOR2_X1 U885 ( .A(n800), .B(n799), .ZN(n892) );
  XNOR2_X1 U886 ( .A(n801), .B(n892), .ZN(n802) );
  NAND2_X1 U887 ( .A1(n802), .A2(G868), .ZN(n806) );
  NAND2_X1 U888 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U889 ( .A1(n806), .A2(n805), .ZN(G295) );
  NAND2_X1 U890 ( .A1(G2078), .A2(G2084), .ZN(n807) );
  XOR2_X1 U891 ( .A(KEYINPUT20), .B(n807), .Z(n808) );
  NAND2_X1 U892 ( .A1(G2090), .A2(n808), .ZN(n810) );
  XNOR2_X1 U893 ( .A(KEYINPUT21), .B(KEYINPUT82), .ZN(n809) );
  XNOR2_X1 U894 ( .A(n810), .B(n809), .ZN(n811) );
  NAND2_X1 U895 ( .A1(G2072), .A2(n811), .ZN(G158) );
  XNOR2_X1 U896 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  XNOR2_X1 U897 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U898 ( .A1(G108), .A2(G120), .ZN(n812) );
  NOR2_X1 U899 ( .A1(G237), .A2(n812), .ZN(n813) );
  NAND2_X1 U900 ( .A1(G69), .A2(n813), .ZN(n826) );
  NAND2_X1 U901 ( .A1(n826), .A2(G567), .ZN(n819) );
  NOR2_X1 U902 ( .A1(G220), .A2(G219), .ZN(n814) );
  XOR2_X1 U903 ( .A(KEYINPUT22), .B(n814), .Z(n815) );
  NOR2_X1 U904 ( .A1(G218), .A2(n815), .ZN(n816) );
  XOR2_X1 U905 ( .A(KEYINPUT83), .B(n816), .Z(n817) );
  NAND2_X1 U906 ( .A1(G96), .A2(n817), .ZN(n827) );
  NAND2_X1 U907 ( .A1(n827), .A2(G2106), .ZN(n818) );
  NAND2_X1 U908 ( .A1(n819), .A2(n818), .ZN(n847) );
  NAND2_X1 U909 ( .A1(G661), .A2(G483), .ZN(n820) );
  NOR2_X1 U910 ( .A1(n847), .A2(n820), .ZN(n823) );
  NAND2_X1 U911 ( .A1(n823), .A2(G36), .ZN(G176) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U914 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G1), .A2(G3), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U917 ( .A(n825), .B(KEYINPUT106), .ZN(G188) );
  INV_X1 U919 ( .A(G120), .ZN(G236) );
  INV_X1 U920 ( .A(G108), .ZN(G238) );
  INV_X1 U921 ( .A(G96), .ZN(G221) );
  INV_X1 U922 ( .A(G69), .ZN(G235) );
  NOR2_X1 U923 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U924 ( .A(G325), .ZN(G261) );
  XOR2_X1 U925 ( .A(KEYINPUT41), .B(G1986), .Z(n829) );
  XNOR2_X1 U926 ( .A(G1996), .B(G1991), .ZN(n828) );
  XNOR2_X1 U927 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U928 ( .A(n830), .B(G2474), .Z(n832) );
  XNOR2_X1 U929 ( .A(G1966), .B(G1981), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U931 ( .A(G1976), .B(G1971), .Z(n834) );
  XNOR2_X1 U932 ( .A(G1961), .B(G1956), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U934 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U935 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(G229) );
  XOR2_X1 U937 ( .A(G2100), .B(G2096), .Z(n840) );
  XNOR2_X1 U938 ( .A(KEYINPUT42), .B(G2678), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U940 ( .A(KEYINPUT43), .B(G2090), .Z(n842) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(G227) );
  INV_X1 U946 ( .A(n847), .ZN(G319) );
  NAND2_X1 U947 ( .A1(G100), .A2(n869), .ZN(n849) );
  NAND2_X1 U948 ( .A1(G112), .A2(n875), .ZN(n848) );
  NAND2_X1 U949 ( .A1(n849), .A2(n848), .ZN(n856) );
  NAND2_X1 U950 ( .A1(G136), .A2(n516), .ZN(n850) );
  XNOR2_X1 U951 ( .A(KEYINPUT109), .B(n850), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n873), .A2(G124), .ZN(n851) );
  XOR2_X1 U953 ( .A(KEYINPUT44), .B(n851), .Z(n852) );
  NOR2_X1 U954 ( .A1(n853), .A2(n852), .ZN(n854) );
  XOR2_X1 U955 ( .A(KEYINPUT110), .B(n854), .Z(n855) );
  NOR2_X1 U956 ( .A1(n856), .A2(n855), .ZN(G162) );
  NAND2_X1 U957 ( .A1(n869), .A2(G106), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G142), .A2(n516), .ZN(n857) );
  NAND2_X1 U959 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n859), .B(KEYINPUT45), .ZN(n861) );
  NAND2_X1 U961 ( .A1(G118), .A2(n875), .ZN(n860) );
  NAND2_X1 U962 ( .A1(n861), .A2(n860), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G130), .A2(n873), .ZN(n862) );
  XNOR2_X1 U964 ( .A(KEYINPUT111), .B(n862), .ZN(n863) );
  NOR2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U966 ( .A(G160), .B(n865), .ZN(n888) );
  XOR2_X1 U967 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n867) );
  XNOR2_X1 U968 ( .A(G164), .B(KEYINPUT46), .ZN(n866) );
  XNOR2_X1 U969 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n962), .B(n868), .ZN(n883) );
  NAND2_X1 U971 ( .A1(n869), .A2(G103), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G139), .A2(n516), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n880) );
  NAND2_X1 U974 ( .A1(n873), .A2(G127), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n874), .B(KEYINPUT112), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G115), .A2(n875), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U978 ( .A(KEYINPUT47), .B(n878), .Z(n879) );
  NOR2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n967) );
  XNOR2_X1 U980 ( .A(n881), .B(n967), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U982 ( .A(G162), .B(n884), .Z(n885) );
  XNOR2_X1 U983 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n890) );
  XOR2_X1 U985 ( .A(n890), .B(n889), .Z(n891) );
  NOR2_X1 U986 ( .A1(G37), .A2(n891), .ZN(G395) );
  XNOR2_X1 U987 ( .A(G286), .B(n999), .ZN(n893) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n894), .B(G171), .ZN(n895) );
  NOR2_X1 U990 ( .A1(G37), .A2(n895), .ZN(G397) );
  XNOR2_X1 U991 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n897) );
  NOR2_X1 U992 ( .A1(G229), .A2(G227), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n910) );
  XNOR2_X1 U994 ( .A(G2446), .B(KEYINPUT104), .ZN(n907) );
  XOR2_X1 U995 ( .A(G2430), .B(G2427), .Z(n899) );
  XNOR2_X1 U996 ( .A(KEYINPUT105), .B(G2438), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n903) );
  XOR2_X1 U998 ( .A(G2435), .B(G2454), .Z(n901) );
  XNOR2_X1 U999 ( .A(G1341), .B(G1348), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1001 ( .A(n903), .B(n902), .Z(n905) );
  XNOR2_X1 U1002 ( .A(G2443), .B(G2451), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  NAND2_X1 U1005 ( .A1(n908), .A2(G14), .ZN(n913) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n913), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(n913), .ZN(G401) );
  XNOR2_X1 U1012 ( .A(G29), .B(KEYINPUT119), .ZN(n934) );
  XNOR2_X1 U1013 ( .A(G2084), .B(G34), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(n914), .B(KEYINPUT54), .ZN(n930) );
  XNOR2_X1 U1015 ( .A(G2090), .B(G35), .ZN(n927) );
  XOR2_X1 U1016 ( .A(G1991), .B(G25), .Z(n915) );
  NAND2_X1 U1017 ( .A1(n915), .A2(G28), .ZN(n924) );
  XNOR2_X1 U1018 ( .A(G1996), .B(G32), .ZN(n917) );
  XNOR2_X1 U1019 ( .A(G33), .B(G2072), .ZN(n916) );
  NOR2_X1 U1020 ( .A1(n917), .A2(n916), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(G2067), .B(G26), .ZN(n920) );
  XNOR2_X1 U1022 ( .A(G27), .B(n918), .ZN(n919) );
  NOR2_X1 U1023 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(KEYINPUT53), .B(n925), .ZN(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(n928), .B(KEYINPUT117), .ZN(n929) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(n931), .B(KEYINPUT118), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(n932), .B(KEYINPUT55), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1033 ( .A(n935), .B(KEYINPUT120), .ZN(n992) );
  XOR2_X1 U1034 ( .A(G16), .B(KEYINPUT124), .Z(n960) );
  XNOR2_X1 U1035 ( .A(KEYINPUT125), .B(G1961), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(n936), .B(G5), .ZN(n955) );
  XNOR2_X1 U1037 ( .A(G1971), .B(G22), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(G1976), .B(G23), .ZN(n937) );
  NOR2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1040 ( .A(KEYINPUT126), .B(n939), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(G1986), .B(KEYINPUT127), .ZN(n940) );
  XNOR2_X1 U1042 ( .A(n940), .B(G24), .ZN(n941) );
  NAND2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1044 ( .A(n943), .B(KEYINPUT58), .ZN(n953) );
  XOR2_X1 U1045 ( .A(G1348), .B(KEYINPUT59), .Z(n944) );
  XNOR2_X1 U1046 ( .A(G4), .B(n944), .ZN(n946) );
  XNOR2_X1 U1047 ( .A(G20), .B(G1956), .ZN(n945) );
  NOR2_X1 U1048 ( .A1(n946), .A2(n945), .ZN(n950) );
  XNOR2_X1 U1049 ( .A(G1341), .B(G19), .ZN(n948) );
  XNOR2_X1 U1050 ( .A(G1981), .B(G6), .ZN(n947) );
  NOR2_X1 U1051 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1052 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1053 ( .A(KEYINPUT60), .B(n951), .ZN(n952) );
  NOR2_X1 U1054 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n957) );
  XNOR2_X1 U1056 ( .A(G21), .B(G1966), .ZN(n956) );
  NOR2_X1 U1057 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1058 ( .A(n958), .B(KEYINPUT61), .ZN(n959) );
  NAND2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n961), .ZN(n990) );
  NOR2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1062 ( .A(KEYINPUT115), .B(n964), .Z(n965) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n984) );
  XOR2_X1 U1064 ( .A(G2072), .B(n967), .Z(n969) );
  XOR2_X1 U1065 ( .A(G164), .B(G2078), .Z(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1067 ( .A(KEYINPUT50), .B(n970), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(n971), .B(KEYINPUT116), .ZN(n982) );
  XNOR2_X1 U1069 ( .A(G160), .B(G2084), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n980) );
  XOR2_X1 U1072 ( .A(G2090), .B(G162), .Z(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(n978), .B(KEYINPUT51), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1078 ( .A(KEYINPUT52), .B(n985), .Z(n986) );
  NOR2_X1 U1079 ( .A1(KEYINPUT55), .A2(n986), .ZN(n988) );
  INV_X1 U1080 ( .A(G29), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n1021) );
  XNOR2_X1 U1084 ( .A(G1966), .B(G168), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(n995), .B(KEYINPUT57), .ZN(n1013) );
  XNOR2_X1 U1087 ( .A(n996), .B(G1956), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1002) );
  XOR2_X1 U1089 ( .A(G1348), .B(n999), .Z(n1000) );
  XNOR2_X1 U1090 ( .A(KEYINPUT121), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1008) );
  NAND2_X1 U1092 ( .A1(G1971), .A2(G303), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1096 ( .A(G1961), .B(G171), .Z(n1009) );
  XNOR2_X1 U1097 ( .A(KEYINPUT122), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1016) );
  XNOR2_X1 U1100 ( .A(G1341), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XOR2_X1 U1102 ( .A(KEYINPUT56), .B(G16), .Z(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1104 ( .A(KEYINPUT123), .B(n1019), .Z(n1020) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(n1022), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

