//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G116), .B(G119), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(KEYINPUT69), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT2), .B(G113), .Z(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n196), .A2(KEYINPUT3), .A3(G107), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT81), .B(G104), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G107), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G101), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n195), .B1(KEYINPUT4), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n199), .B(new_n205), .C1(new_n200), .C2(new_n201), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT82), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n206), .A2(KEYINPUT4), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT82), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(new_n203), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n204), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT83), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n196), .A2(G107), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n198), .B2(G107), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n213), .B1(new_n215), .B2(G101), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n206), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n213), .A3(G101), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n191), .A2(KEYINPUT5), .ZN(new_n220));
  INV_X1    g034(.A(G116), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n221), .A2(KEYINPUT5), .A3(G119), .ZN(new_n222));
  INV_X1    g036(.A(G113), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n220), .A2(new_n224), .B1(new_n193), .B2(new_n191), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n219), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n190), .B1(new_n212), .B2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n203), .A2(KEYINPUT4), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(new_n194), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n210), .B1(new_n209), .B2(new_n203), .ZN(new_n231));
  AND4_X1   g045(.A1(new_n210), .A2(new_n203), .A3(KEYINPUT4), .A4(new_n206), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(new_n226), .A3(new_n189), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT85), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n228), .A2(new_n234), .A3(new_n235), .A4(KEYINPUT6), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n228), .A2(new_n234), .A3(KEYINPUT6), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT6), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n238), .B(new_n190), .C1(new_n212), .C2(new_n227), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT85), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n236), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G128), .ZN(new_n242));
  INV_X1    g056(.A(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G143), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n242), .B1(new_n244), .B2(KEYINPUT1), .ZN(new_n245));
  XNOR2_X1  g059(.A(G143), .B(G146), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G125), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT76), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT76), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G125), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT88), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n246), .A2(KEYINPUT0), .A3(G128), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT0), .B(G128), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n256), .B1(new_n246), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT86), .A3(new_n252), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT86), .B1(new_n258), .B2(new_n252), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT87), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT87), .B1(new_n260), .B2(new_n261), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n255), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G224), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(G953), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n266), .B(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n241), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n268), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT7), .B1(new_n272), .B2(KEYINPUT90), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(KEYINPUT90), .B2(new_n272), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n253), .B(KEYINPUT88), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n262), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n272), .A2(KEYINPUT7), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n266), .A2(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n189), .B(KEYINPUT8), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n219), .A2(new_n225), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n279), .B1(new_n227), .B2(new_n280), .ZN(new_n281));
  OR2_X1    g095(.A1(new_n281), .A2(KEYINPUT89), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(KEYINPUT89), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n278), .A2(new_n282), .A3(new_n234), .A4(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G210), .B1(G237), .B2(G902), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n271), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n287), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n228), .A2(new_n234), .A3(KEYINPUT6), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(KEYINPUT85), .A3(new_n239), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n269), .B1(new_n291), .B2(new_n236), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n284), .A2(new_n285), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n188), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT20), .ZN(new_n296));
  XNOR2_X1  g110(.A(G113), .B(G122), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(new_n196), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT71), .B(G237), .Z(new_n300));
  INV_X1    g114(.A(G953), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(G214), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G143), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT71), .B(G237), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(G953), .ZN(new_n306));
  AOI21_X1  g120(.A(G143), .B1(new_n306), .B2(G214), .ZN(new_n307));
  OAI211_X1 g121(.A(KEYINPUT18), .B(G131), .C1(new_n304), .C2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G125), .B(G140), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n243), .ZN(new_n310));
  INV_X1    g124(.A(G140), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G125), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT76), .B(G125), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(G140), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n310), .B1(new_n315), .B2(new_n243), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n302), .A2(new_n303), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n306), .A2(G143), .A3(G214), .ZN(new_n318));
  NAND2_X1  g132(.A1(KEYINPUT18), .A2(G131), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n308), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n249), .A2(new_n251), .A3(G140), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT16), .A3(new_n312), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT16), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n252), .A2(new_n325), .A3(new_n311), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(G146), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT19), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n309), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n315), .B2(new_n328), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n327), .B1(new_n330), .B2(G146), .ZN(new_n331));
  OAI21_X1  g145(.A(G131), .B1(new_n304), .B2(new_n307), .ZN(new_n332));
  INV_X1    g146(.A(G131), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n317), .A2(new_n333), .A3(new_n318), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n331), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n299), .B1(new_n322), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT17), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n332), .A2(new_n337), .A3(new_n334), .ZN(new_n338));
  INV_X1    g152(.A(new_n327), .ZN(new_n339));
  AOI21_X1  g153(.A(G146), .B1(new_n324), .B2(new_n326), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n332), .B2(new_n337), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n298), .B(new_n321), .C1(new_n338), .C2(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n336), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(G475), .A2(G902), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n296), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n336), .A2(new_n343), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(KEYINPUT20), .A3(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n321), .B1(new_n338), .B2(new_n342), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n299), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n343), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n285), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT92), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT91), .B(G475), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(G902), .B1(new_n352), .B2(new_n343), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n358), .B1(new_n359), .B2(KEYINPUT92), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n350), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G134), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT95), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n242), .B2(G143), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n303), .A2(KEYINPUT95), .A3(G128), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n303), .A2(G128), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n363), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(KEYINPUT13), .B2(new_n367), .ZN(new_n371));
  NAND2_X1  g185(.A1(KEYINPUT13), .A2(G134), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT94), .ZN(new_n374));
  INV_X1    g188(.A(G122), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n374), .B1(new_n375), .B2(G116), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n221), .A2(KEYINPUT94), .A3(G122), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(KEYINPUT93), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT93), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G122), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n221), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G107), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n384), .A2(new_n385), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n371), .B(new_n373), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT9), .B(G234), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT80), .ZN(new_n391));
  INV_X1    g205(.A(G217), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n391), .A2(new_n392), .A3(G953), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n383), .B1(KEYINPUT14), .B2(new_n378), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT96), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n378), .A2(KEYINPUT14), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n397), .A2(KEYINPUT97), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n395), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(KEYINPUT97), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n396), .A2(new_n398), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n401), .A2(G107), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n368), .A2(new_n363), .A3(new_n369), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n386), .B1(new_n403), .B2(new_n370), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n389), .B(new_n393), .C1(new_n402), .C2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n393), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n404), .B1(new_n401), .B2(G107), .ZN(new_n407));
  INV_X1    g221(.A(new_n389), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(G902), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G478), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(KEYINPUT15), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n410), .B(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n362), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(G234), .A2(G237), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n416), .A2(G902), .A3(G953), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT21), .B(G898), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n416), .A2(G952), .A3(new_n301), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n295), .A2(new_n415), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT68), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT64), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT11), .ZN(new_n426));
  INV_X1    g240(.A(G137), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n425), .A2(new_n426), .A3(new_n427), .A4(G134), .ZN(new_n428));
  OAI22_X1  g242(.A1(new_n363), .A2(G137), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n427), .B2(G134), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(KEYINPUT66), .A3(G131), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT66), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n432), .B1(new_n429), .B2(new_n428), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n436), .B1(new_n437), .B2(new_n333), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n430), .A2(new_n433), .A3(new_n333), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT65), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n437), .A2(KEYINPUT65), .A3(new_n333), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n258), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n247), .ZN(new_n446));
  XOR2_X1   g260(.A(G134), .B(G137), .Z(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G131), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n440), .A2(new_n441), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT65), .B1(new_n437), .B2(new_n333), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT67), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n446), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n442), .A2(new_n443), .B1(G131), .B2(new_n447), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT67), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n445), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n424), .B1(new_n456), .B2(KEYINPUT30), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n439), .A2(new_n444), .ZN(new_n458));
  INV_X1    g272(.A(new_n258), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n247), .B1(new_n454), .B2(KEYINPUT67), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n451), .A2(new_n452), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT30), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(KEYINPUT68), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT70), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n454), .A2(new_n247), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n445), .A2(KEYINPUT70), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n467), .A2(KEYINPUT30), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n457), .A2(new_n465), .A3(new_n195), .A4(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n467), .A2(new_n194), .A3(new_n468), .A4(new_n469), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n306), .A2(G210), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT27), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT26), .B(G101), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT29), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n469), .A2(new_n468), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT73), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n481), .A2(new_n482), .A3(new_n194), .A4(new_n467), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n472), .A2(KEYINPUT73), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n195), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT28), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n460), .A2(new_n194), .A3(new_n468), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT28), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT74), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n491), .B(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n479), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n463), .A2(new_n195), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n497), .B1(new_n498), .B2(new_n472), .ZN(new_n499));
  INV_X1    g313(.A(new_n491), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n477), .B1(new_n501), .B2(KEYINPUT29), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n480), .B(new_n285), .C1(new_n495), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G472), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT32), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n472), .A2(new_n477), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n471), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT31), .ZN(new_n508));
  INV_X1    g322(.A(new_n477), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n499), .B2(new_n500), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT31), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n471), .A2(new_n511), .A3(new_n506), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(G472), .A2(G902), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n505), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n514), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(KEYINPUT32), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n504), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n392), .B1(G234), .B2(new_n285), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT78), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n327), .A2(new_n310), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT24), .B(G110), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT75), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n242), .A2(G119), .ZN(new_n525));
  INV_X1    g339(.A(G119), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(G128), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(G128), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n242), .A2(G119), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT75), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n523), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT23), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n526), .B2(G128), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n242), .A2(KEYINPUT23), .A3(G119), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n529), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(G110), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT77), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT75), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT75), .B1(new_n529), .B2(new_n530), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n522), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n534), .A2(new_n529), .A3(new_n535), .ZN(new_n542));
  INV_X1    g356(.A(G110), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT77), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n541), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n521), .B1(new_n538), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n528), .A2(new_n523), .A3(new_n531), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n543), .B2(new_n542), .ZN(new_n549));
  INV_X1    g363(.A(new_n340), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n550), .B2(new_n327), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n520), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n327), .A2(new_n310), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n532), .A2(new_n537), .A3(KEYINPUT77), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n545), .B1(new_n541), .B2(new_n544), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n536), .A2(G110), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n548), .B(new_n557), .C1(new_n339), .C2(new_n340), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(KEYINPUT78), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT22), .B(G137), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n301), .A2(G221), .A3(G234), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n560), .B(new_n561), .Z(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n552), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n556), .A2(new_n558), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(new_n520), .A3(new_n562), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT25), .B1(new_n567), .B2(new_n285), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT25), .ZN(new_n569));
  AOI211_X1 g383(.A(new_n569), .B(G902), .C1(new_n564), .C2(new_n566), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n519), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT79), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(KEYINPUT79), .B(new_n519), .C1(new_n568), .C2(new_n570), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n519), .A2(G902), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n567), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G221), .ZN(new_n580));
  INV_X1    g394(.A(new_n391), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n581), .B2(new_n285), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n219), .A2(new_n247), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n446), .B1(new_n217), .B2(new_n218), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n458), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT12), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n218), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n206), .B2(new_n216), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n446), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n219), .A2(new_n247), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(KEYINPUT12), .A3(new_n458), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n229), .A2(new_n258), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n231), .B2(new_n232), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT10), .B1(new_n589), .B2(new_n446), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n584), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n458), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n596), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n594), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(G110), .B(G140), .ZN(new_n604));
  INV_X1    g418(.A(G227), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(G953), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n604), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT84), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n601), .B1(new_n596), .B2(new_n600), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n607), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n602), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n608), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n596), .A2(new_n600), .A3(new_n601), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n615), .A2(new_n610), .A3(new_n607), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n612), .B1(new_n594), .B2(new_n602), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT84), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n614), .A2(new_n618), .A3(G469), .ZN(new_n619));
  INV_X1    g433(.A(G469), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n285), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n607), .B1(new_n615), .B2(new_n610), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n594), .A2(new_n602), .A3(new_n612), .ZN(new_n623));
  AOI21_X1  g437(.A(G902), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n621), .B1(new_n624), .B2(new_n620), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n582), .B1(new_n619), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n423), .A2(new_n518), .A3(new_n579), .A4(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT98), .B(G101), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G3));
  AND4_X1   g443(.A1(new_n575), .A2(new_n295), .A3(new_n577), .A4(new_n422), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n513), .A2(new_n285), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(G472), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n626), .A2(new_n632), .A3(new_n516), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n405), .A2(new_n409), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT33), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n405), .A2(new_n409), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(G478), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n410), .A2(new_n411), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n411), .A2(new_n285), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n362), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n634), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT34), .B(G104), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NAND2_X1  g462(.A1(new_n361), .A2(new_n414), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n634), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT35), .B(G107), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  NOR2_X1   g466(.A1(new_n563), .A2(KEYINPUT36), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n565), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n576), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n573), .A2(new_n574), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n573), .A2(KEYINPUT99), .A3(new_n574), .A4(new_n655), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n423), .A2(new_n633), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT37), .B(G110), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT100), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n661), .B(new_n663), .ZN(G12));
  AND2_X1   g478(.A1(new_n295), .A2(new_n626), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n356), .A2(new_n360), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n347), .A2(new_n349), .ZN(new_n667));
  INV_X1    g481(.A(new_n417), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n421), .B1(new_n668), .B2(G900), .ZN(new_n669));
  AND4_X1   g483(.A1(new_n414), .A2(new_n666), .A3(new_n667), .A4(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n665), .A2(new_n518), .A3(new_n660), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  XNOR2_X1  g486(.A(new_n669), .B(KEYINPUT39), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n626), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT40), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n285), .B1(new_n487), .B2(new_n477), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n509), .B1(new_n471), .B2(new_n472), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n678), .B1(new_n517), .B2(new_n515), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n288), .A2(new_n294), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n410), .B(new_n412), .ZN(new_n683));
  NOR4_X1   g497(.A1(new_n660), .A2(new_n683), .A3(new_n361), .A4(new_n188), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n675), .A2(new_n679), .A3(new_n682), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G143), .ZN(G45));
  NAND3_X1  g500(.A1(new_n362), .A2(new_n644), .A3(new_n669), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n658), .B2(new_n659), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n665), .A2(new_n518), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G146), .ZN(G48));
  NOR2_X1   g504(.A1(new_n624), .A2(new_n620), .ZN(new_n691));
  AOI211_X1 g505(.A(G469), .B(G902), .C1(new_n622), .C2(new_n623), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n691), .A2(new_n692), .A3(new_n582), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n295), .A2(new_n422), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n361), .A2(new_n643), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n694), .A2(new_n518), .A3(new_n579), .A4(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT41), .B(G113), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT102), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n696), .B(new_n698), .ZN(G15));
  INV_X1    g513(.A(new_n649), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n694), .A2(new_n518), .A3(new_n579), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  NAND4_X1  g516(.A1(new_n423), .A2(new_n518), .A3(new_n660), .A4(new_n693), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT103), .B(G119), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G21));
  AOI21_X1  g519(.A(new_n493), .B1(new_n487), .B2(KEYINPUT28), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n508), .B(new_n512), .C1(new_n706), .C2(new_n477), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n514), .B(KEYINPUT104), .Z(new_n708));
  AOI22_X1  g522(.A1(new_n631), .A2(G472), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n579), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n693), .A2(new_n422), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n361), .A2(new_n683), .ZN(new_n712));
  AND4_X1   g526(.A1(KEYINPUT105), .A2(new_n680), .A3(new_n187), .A4(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT105), .B1(new_n295), .B2(new_n712), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n710), .B(new_n711), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  NAND2_X1  g530(.A1(new_n295), .A2(new_n693), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n687), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n660), .A2(KEYINPUT106), .A3(new_n709), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT106), .B1(new_n660), .B2(new_n709), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(KEYINPUT107), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  NAND3_X1  g540(.A1(new_n288), .A2(new_n294), .A3(new_n187), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n687), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n616), .A2(new_n617), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n621), .B1(new_n729), .B2(G469), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n624), .A2(new_n620), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n582), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n518), .A2(new_n579), .A3(new_n728), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT42), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n333), .ZN(G33));
  INV_X1    g549(.A(new_n670), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n727), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n518), .A2(new_n579), .A3(new_n732), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G134), .ZN(G36));
  NOR2_X1   g553(.A1(new_n362), .A2(new_n643), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT43), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n632), .A2(new_n516), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n742), .A3(new_n660), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n727), .B1(new_n743), .B2(new_n744), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n582), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n729), .A2(KEYINPUT45), .ZN(new_n749));
  XOR2_X1   g563(.A(new_n749), .B(KEYINPUT108), .Z(new_n750));
  AOI21_X1  g564(.A(KEYINPUT45), .B1(new_n614), .B2(new_n618), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n620), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n621), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT46), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n731), .B1(new_n753), .B2(KEYINPUT46), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n748), .B(new_n673), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n747), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g572(.A(KEYINPUT109), .B(G137), .Z(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT110), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n758), .B(new_n760), .ZN(G39));
  NOR4_X1   g575(.A1(new_n518), .A2(new_n579), .A3(new_n687), .A4(new_n727), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n750), .A2(new_n752), .ZN(new_n763));
  INV_X1    g577(.A(new_n621), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n692), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n582), .B1(new_n767), .B2(new_n754), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(KEYINPUT47), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n770));
  AOI211_X1 g584(.A(new_n770), .B(new_n582), .C1(new_n767), .C2(new_n754), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n762), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  NOR2_X1   g587(.A1(G952), .A2(G953), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT118), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n741), .A2(new_n420), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n710), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n727), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n769), .A2(new_n771), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n691), .A2(new_n692), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n582), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n782), .B(KEYINPUT116), .Z(new_n783));
  OAI21_X1  g597(.A(new_n778), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n693), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n682), .A2(new_n187), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n710), .A3(new_n776), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n660), .A2(new_n709), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT106), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n660), .A2(KEYINPUT106), .A3(new_n709), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n785), .A2(new_n727), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n776), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n679), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n579), .A3(new_n420), .A4(new_n795), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n361), .A3(new_n643), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n789), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT51), .B1(new_n784), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n789), .A2(KEYINPUT51), .A3(new_n796), .A4(new_n800), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n779), .A2(new_n782), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n803), .B1(new_n804), .B2(new_n778), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n518), .A2(new_n575), .A3(new_n577), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n776), .A2(new_n806), .A3(new_n795), .ZN(new_n807));
  NAND2_X1  g621(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g623(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n810));
  AOI21_X1  g624(.A(new_n809), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(G952), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n812), .B(G953), .C1(new_n799), .C2(new_n695), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n811), .B(new_n813), .C1(new_n717), .C2(new_n777), .ZN(new_n814));
  OR3_X1    g628(.A1(new_n802), .A2(new_n805), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n671), .A2(new_n689), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n713), .A2(new_n714), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n575), .A2(new_n732), .A3(new_n655), .A4(new_n669), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n679), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT107), .B1(new_n794), .B2(new_n718), .ZN(new_n823));
  INV_X1    g637(.A(new_n724), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n817), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n816), .B1(new_n723), .B2(new_n724), .ZN(new_n827));
  INV_X1    g641(.A(new_n818), .ZN(new_n828));
  INV_X1    g642(.A(new_n820), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n825), .A2(new_n826), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n361), .A2(new_n832), .A3(new_n683), .A4(new_n669), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n666), .A2(new_n683), .A3(new_n667), .A4(new_n669), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT113), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n626), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n727), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n518), .A2(new_n836), .A3(new_n660), .A4(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n838), .A2(new_n738), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n728), .B(new_n732), .C1(new_n719), .C2(new_n720), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n645), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n695), .A2(KEYINPUT112), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n649), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n630), .A2(new_n633), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n627), .A3(new_n661), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n715), .A2(new_n696), .A3(new_n701), .A4(new_n703), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n734), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT53), .B1(new_n831), .B2(new_n851), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n830), .B(new_n817), .C1(new_n823), .C2(new_n824), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n827), .A2(KEYINPUT114), .A3(new_n830), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n855), .A2(new_n856), .B1(new_n826), .B2(new_n825), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n848), .A2(new_n850), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n852), .B(KEYINPUT54), .C1(new_n857), .C2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n859), .B1(new_n831), .B2(new_n851), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT115), .B1(new_n841), .B2(new_n847), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n846), .A2(new_n627), .A3(new_n661), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n866), .A3(new_n840), .A4(new_n839), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n864), .A2(KEYINPUT53), .A3(new_n850), .A4(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n862), .B(new_n863), .C1(new_n857), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n861), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n775), .B1(new_n815), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n579), .A2(new_n748), .A3(new_n187), .A4(new_n740), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT111), .Z(new_n873));
  XOR2_X1   g687(.A(new_n781), .B(KEYINPUT49), .Z(new_n874));
  OR4_X1    g688(.A1(new_n679), .A2(new_n873), .A3(new_n682), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n871), .A2(new_n875), .ZN(G75));
  NOR2_X1   g690(.A1(new_n301), .A2(G952), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n855), .A2(new_n856), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n825), .A2(new_n826), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n868), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n821), .B(new_n816), .C1(new_n723), .C2(new_n724), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n853), .B1(new_n882), .B2(KEYINPUT52), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT53), .B1(new_n883), .B2(new_n858), .ZN(new_n884));
  OAI211_X1 g698(.A(G210), .B(G902), .C1(new_n881), .C2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n241), .B(new_n269), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n885), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n886), .B1(new_n885), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n878), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT56), .B1(new_n885), .B2(KEYINPUT119), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n862), .B1(new_n857), .B2(new_n868), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n895), .A2(new_n896), .A3(G210), .A4(G902), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n888), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n893), .A2(new_n898), .ZN(G51));
  NAND2_X1  g713(.A1(new_n895), .A2(KEYINPUT54), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n869), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n621), .B(KEYINPUT57), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n622), .A2(new_n623), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n895), .A2(G902), .A3(new_n750), .A4(new_n752), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n877), .B1(new_n905), .B2(new_n906), .ZN(G54));
  NAND4_X1  g721(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n908), .A2(new_n344), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n344), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n877), .ZN(G60));
  XNOR2_X1  g725(.A(new_n641), .B(KEYINPUT59), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n870), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n636), .A2(new_n638), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(KEYINPUT121), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n912), .B1(new_n861), .B2(new_n869), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n919), .B2(new_n915), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n916), .A2(new_n912), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n877), .B1(new_n901), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n917), .A2(new_n920), .A3(new_n922), .ZN(G63));
  XNOR2_X1  g737(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n392), .A2(new_n285), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n895), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n927), .A2(new_n566), .A3(new_n564), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n895), .A2(new_n654), .A3(new_n926), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n928), .A2(new_n878), .A3(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n928), .A2(KEYINPUT61), .A3(new_n878), .A4(new_n929), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(G66));
  OAI21_X1  g748(.A(G953), .B1(new_n418), .B2(new_n267), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n849), .A2(new_n847), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(G953), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n291), .B(new_n236), .C1(G898), .C2(new_n301), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT123), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n937), .B(new_n939), .ZN(G69));
  OR2_X1    g754(.A1(new_n747), .A2(new_n757), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n772), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n827), .A2(new_n685), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n806), .A2(new_n674), .A3(new_n837), .A4(new_n845), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n942), .A2(new_n944), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n457), .A2(new_n465), .A3(new_n470), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT124), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(new_n330), .Z(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(G953), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n301), .A2(G900), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n828), .A2(new_n806), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n738), .B1(new_n757), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(new_n734), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n956), .A2(new_n772), .A3(new_n941), .A4(new_n827), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n953), .B1(new_n957), .B2(new_n301), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n958), .A2(KEYINPUT125), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n950), .B1(new_n958), .B2(KEYINPUT125), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n952), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(G900), .ZN(new_n962));
  OAI21_X1  g776(.A(G953), .B1(new_n605), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n963), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n952), .B(new_n965), .C1(new_n959), .C2(new_n960), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(G72));
  XNOR2_X1  g781(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n968));
  NAND2_X1  g782(.A1(G472), .A2(G902), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n936), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n970), .B1(new_n947), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n677), .ZN(new_n973));
  INV_X1    g787(.A(new_n478), .ZN(new_n974));
  INV_X1    g788(.A(new_n677), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n975), .A3(new_n970), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT127), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n852), .B(new_n977), .C1(new_n857), .C2(new_n860), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n970), .B1(new_n957), .B2(new_n971), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n877), .B1(new_n979), .B2(new_n478), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n973), .A2(new_n978), .A3(new_n980), .ZN(G57));
endmodule


