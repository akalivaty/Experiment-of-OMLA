//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT26), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT26), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n203), .B(new_n204), .C1(new_n207), .C2(new_n202), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT27), .B(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT28), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(KEYINPUT28), .A3(new_n210), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n208), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217));
  AND2_X1   g016(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n204), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n220), .B1(new_n204), .B2(new_n221), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n219), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n219), .B(new_n226), .C1(new_n222), .C2(new_n223), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT23), .B1(new_n202), .B2(KEYINPUT64), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n229), .B(new_n230), .C1(G169gat), .C2(G176gat), .ZN(new_n231));
  AND4_X1   g030(.A1(KEYINPUT25), .A2(new_n228), .A3(new_n231), .A4(new_n205), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n225), .A2(new_n227), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n204), .A2(new_n221), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n219), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n228), .A2(new_n231), .A3(new_n205), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n233), .A2(KEYINPUT67), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT67), .B1(new_n233), .B2(new_n238), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n216), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G134gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G127gat), .ZN(new_n243));
  INV_X1    g042(.A(G127gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G134gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(KEYINPUT1), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n248));
  INV_X1    g047(.A(G113gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n248), .B1(new_n249), .B2(G120gat), .ZN(new_n250));
  INV_X1    g049(.A(G120gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n250), .B(new_n252), .C1(G113gat), .C2(new_n251), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n249), .A2(G120gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n251), .A2(G113gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n247), .A2(new_n253), .B1(new_n257), .B2(new_n246), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n258), .A2(KEYINPUT69), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(KEYINPUT69), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G227gat), .ZN(new_n263));
  INV_X1    g062(.A(G233gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n216), .B(new_n259), .C1(new_n239), .C2(new_n240), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n262), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT34), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G15gat), .B(G43gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT71), .ZN(new_n272));
  XNOR2_X1  g071(.A(G71gat), .B(G99gat), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n272), .B(new_n273), .Z(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n233), .A2(new_n238), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n233), .A2(KEYINPUT67), .A3(new_n238), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n215), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n261), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n267), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n265), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT33), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n275), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT70), .B1(new_n283), .B2(KEYINPUT32), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT32), .ZN(new_n288));
  AOI211_X1 g087(.A(new_n287), .B(new_n288), .C1(new_n282), .C2(new_n265), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n285), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(KEYINPUT72), .B(new_n285), .C1(new_n286), .C2(new_n289), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n266), .B1(new_n262), .B2(new_n267), .ZN(new_n295));
  AOI211_X1 g094(.A(new_n288), .B(new_n295), .C1(KEYINPUT33), .C2(new_n274), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n270), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  AOI211_X1 g097(.A(new_n269), .B(new_n296), .C1(new_n292), .C2(new_n293), .ZN(new_n299));
  XNOR2_X1  g098(.A(G78gat), .B(G106gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(G22gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G197gat), .B(G204gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT22), .ZN(new_n304));
  INV_X1    g103(.A(G211gat), .ZN(new_n305));
  INV_X1    g104(.A(G218gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G211gat), .B(G218gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT3), .ZN(new_n313));
  NAND2_X1  g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G141gat), .ZN(new_n317));
  INV_X1    g116(.A(G148gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G141gat), .A2(G148gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n314), .B(new_n316), .C1(new_n321), .C2(KEYINPUT2), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT78), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n316), .A2(new_n323), .A3(new_n314), .ZN(new_n324));
  AND2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT78), .B1(new_n325), .B2(new_n315), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n319), .A2(new_n327), .A3(new_n320), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n324), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT2), .ZN(new_n330));
  AND2_X1   g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n330), .B1(new_n333), .B2(new_n327), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n313), .B(new_n322), .C1(new_n329), .C2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n311), .B1(new_n312), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(G228gat), .A2(G233gat), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n309), .A2(new_n303), .A3(KEYINPUT82), .A4(new_n307), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n339), .B(new_n312), .C1(new_n311), .C2(KEYINPUT82), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n322), .B1(new_n329), .B2(new_n334), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT80), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n343), .B(new_n322), .C1(new_n329), .C2(new_n334), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n340), .A2(new_n313), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  OR2_X1    g144(.A1(new_n338), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n313), .B1(new_n310), .B2(KEYINPUT29), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n347), .A2(new_n341), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n337), .B1(new_n348), .B2(new_n336), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT31), .B(G50gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n346), .B2(new_n349), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n302), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n354), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n356), .A2(new_n301), .A3(new_n352), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n298), .A2(new_n299), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT85), .B(KEYINPUT35), .ZN(new_n360));
  XNOR2_X1  g159(.A(G8gat), .B(G36gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(G64gat), .B(G92gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT74), .ZN(new_n364));
  AND2_X1   g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n276), .A2(new_n365), .A3(new_n216), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(KEYINPUT29), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n311), .B(new_n366), .C1(new_n241), .C2(new_n367), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n365), .B(new_n216), .C1(new_n239), .C2(new_n240), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n215), .B1(new_n233), .B2(new_n238), .ZN(new_n370));
  INV_X1    g169(.A(new_n367), .ZN(new_n371));
  OR2_X1    g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n310), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n364), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT75), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n369), .A2(new_n372), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n311), .ZN(new_n378));
  INV_X1    g177(.A(new_n366), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n379), .B(new_n310), .C1(new_n280), .C2(new_n371), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(KEYINPUT75), .A3(new_n364), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n378), .A2(new_n380), .A3(new_n363), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT76), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT30), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n378), .A2(new_n380), .A3(new_n387), .A4(new_n363), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n384), .A2(new_n386), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n383), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(G1gat), .B(G29gat), .Z(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(KEYINPUT0), .ZN(new_n393));
  XNOR2_X1  g192(.A(G57gat), .B(G85gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n342), .A2(KEYINPUT4), .A3(new_n258), .A4(new_n344), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n341), .A2(KEYINPUT3), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n247), .A2(new_n253), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n257), .A2(new_n246), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(new_n400), .A3(new_n335), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n321), .A2(KEYINPUT77), .B1(KEYINPUT2), .B2(new_n314), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n402), .A2(new_n324), .A3(new_n328), .A4(new_n326), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n258), .A3(new_n322), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(G225gat), .A2(G233gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n407), .B(KEYINPUT79), .Z(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n396), .A2(new_n401), .A3(new_n406), .A4(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT5), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n341), .A2(new_n400), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n404), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n413), .B2(new_n408), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n342), .A2(new_n405), .A3(new_n258), .A4(new_n344), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n404), .A2(KEYINPUT4), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n258), .B1(new_n341), .B2(KEYINPUT3), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n408), .B1(new_n419), .B2(new_n335), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n411), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n395), .B1(new_n415), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT6), .ZN(new_n423));
  INV_X1    g222(.A(new_n422), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n415), .A2(new_n395), .A3(new_n421), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI211_X1 g226(.A(new_n360), .B(new_n391), .C1(new_n423), .C2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n293), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n287), .B1(new_n295), .B2(new_n288), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n283), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT72), .B1(new_n432), .B2(new_n285), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n297), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n269), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n425), .B(new_n426), .C1(new_n422), .C2(KEYINPUT81), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n422), .A2(KEYINPUT81), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n423), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n383), .A2(new_n438), .A3(new_n389), .A4(new_n390), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n270), .B(new_n297), .C1(new_n429), .C2(new_n433), .ZN(new_n441));
  INV_X1    g240(.A(new_n358), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n435), .A2(new_n440), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n359), .A2(new_n428), .B1(new_n443), .B2(KEYINPUT35), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n427), .A2(new_n385), .A3(new_n423), .A4(new_n388), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT38), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n378), .A2(new_n380), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n377), .A2(new_n310), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n379), .B(new_n311), .C1(new_n280), .C2(new_n371), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(KEYINPUT37), .A3(new_n450), .ZN(new_n451));
  AND4_X1   g250(.A1(new_n446), .A2(new_n448), .A3(new_n451), .A4(new_n364), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n445), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n363), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n447), .B1(new_n378), .B2(new_n380), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT38), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n358), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n409), .B1(new_n418), .B2(new_n401), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT39), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT39), .B1(new_n413), .B2(new_n408), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n461), .B(new_n395), .C1(new_n459), .C2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT40), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT84), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n463), .A2(new_n464), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n466), .A2(new_n391), .A3(new_n424), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n458), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT73), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n471), .B(KEYINPUT36), .C1(new_n298), .C2(new_n299), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT36), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n294), .A2(new_n471), .A3(new_n270), .A4(new_n297), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n473), .B(new_n474), .C1(new_n435), .C2(KEYINPUT73), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n439), .A2(new_n358), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n470), .B1(new_n477), .B2(KEYINPUT83), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n472), .A2(new_n475), .A3(new_n479), .A4(new_n476), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n444), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT87), .B1(G29gat), .B2(G36gat), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT14), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n483), .A2(new_n484), .B1(G29gat), .B2(G36gat), .ZN(new_n485));
  OR3_X1    g284(.A1(KEYINPUT87), .A2(G29gat), .A3(G36gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(KEYINPUT14), .A3(new_n482), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(G43gat), .B(G50gat), .Z(new_n489));
  AND2_X1   g288(.A1(new_n489), .A2(KEYINPUT88), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT15), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(new_n488), .B2(new_n489), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n492), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT17), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n494), .A2(new_n491), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT89), .B(KEYINPUT17), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n492), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G1gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT16), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n501), .B(KEYINPUT90), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n504), .ZN(new_n508));
  INV_X1    g307(.A(G8gat), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n509), .B1(new_n506), .B2(new_n508), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n500), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT91), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n497), .B(new_n492), .C1(new_n510), .C2(new_n511), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n513), .A2(KEYINPUT18), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT18), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n512), .A2(new_n495), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n516), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n515), .B(KEYINPUT13), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(G169gat), .B(G197gat), .Z(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT12), .ZN(new_n531));
  AND4_X1   g330(.A1(new_n517), .A2(new_n520), .A3(new_n525), .A4(new_n531), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n518), .A2(new_n519), .B1(new_n522), .B2(new_n524), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n531), .B1(new_n533), .B2(new_n517), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT98), .ZN(new_n536));
  INV_X1    g335(.A(G57gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT92), .ZN(new_n538));
  INV_X1    g337(.A(G64gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(KEYINPUT92), .A2(G64gat), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n542), .A2(new_n543), .B1(new_n537), .B2(G64gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n541), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(G57gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT93), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G71gat), .B(G78gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT94), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n550), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT9), .ZN(new_n553));
  INV_X1    g352(.A(G71gat), .ZN(new_n554));
  INV_X1    g353(.A(G78gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n548), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G57gat), .B(G64gat), .Z(new_n559));
  AOI21_X1  g358(.A(new_n549), .B1(new_n559), .B2(KEYINPUT9), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G85gat), .A2(G92gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT7), .ZN(new_n564));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  INV_X1    g364(.A(G85gat), .ZN(new_n566));
  INV_X1    g365(.A(G92gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(KEYINPUT8), .A2(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G99gat), .B(G106gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT96), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n564), .A2(new_n570), .A3(new_n568), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n570), .B1(new_n564), .B2(new_n568), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT96), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n574), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n558), .B(new_n561), .C1(new_n576), .C2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT10), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n578), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT10), .ZN(new_n584));
  NOR3_X1   g383(.A1(new_n583), .A2(new_n562), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n536), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n551), .A2(new_n556), .A3(new_n552), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n547), .B2(new_n544), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n580), .A2(new_n576), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n588), .A2(new_n589), .A3(new_n560), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n558), .A2(new_n561), .B1(new_n575), .B2(new_n577), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n584), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n588), .A2(new_n560), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(new_n578), .A3(KEYINPUT10), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(KEYINPUT98), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n586), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n590), .A2(new_n591), .A3(new_n596), .ZN(new_n598));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT99), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n597), .A2(KEYINPUT99), .A3(new_n603), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n582), .A2(new_n585), .ZN(new_n609));
  INV_X1    g408(.A(new_n596), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n602), .B1(new_n611), .B2(new_n598), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT100), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n597), .A2(KEYINPUT99), .A3(new_n603), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT99), .B1(new_n597), .B2(new_n603), .ZN(new_n615));
  OAI211_X1 g414(.A(KEYINPUT100), .B(new_n612), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(G231gat), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT21), .ZN(new_n620));
  AOI211_X1 g419(.A(new_n619), .B(new_n264), .C1(new_n562), .C2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n619), .A2(new_n264), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n593), .A2(KEYINPUT21), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(G127gat), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G183gat), .B(G211gat), .Z(new_n626));
  NOR3_X1   g425(.A1(new_n621), .A2(new_n623), .A3(G127gat), .ZN(new_n627));
  OR3_X1    g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n626), .B1(new_n625), .B2(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n631));
  INV_X1    g430(.A(G155gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n512), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n562), .A2(new_n620), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT95), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n634), .A2(KEYINPUT95), .A3(new_n635), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n638), .ZN(new_n640));
  INV_X1    g439(.A(new_n633), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n636), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n630), .A2(new_n643), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n628), .A2(new_n629), .B1(new_n642), .B2(new_n639), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n583), .A2(new_n495), .ZN(new_n646));
  AND3_X1   g445(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n496), .A2(new_n500), .A3(new_n583), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(G190gat), .B(G218gat), .Z(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n651), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n648), .A2(new_n653), .A3(new_n649), .ZN(new_n654));
  XNOR2_X1  g453(.A(G134gat), .B(G162gat), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(KEYINPUT97), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n657), .A2(KEYINPUT97), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n652), .B(new_n654), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n652), .A2(new_n654), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n660), .B1(new_n661), .B2(new_n659), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n644), .A2(new_n645), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n618), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n481), .A2(new_n535), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n438), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(new_n391), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n665), .ZN(new_n671));
  INV_X1    g470(.A(new_n391), .ZN(new_n672));
  OAI21_X1  g471(.A(G8gat), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n670), .ZN(new_n674));
  MUX2_X1   g473(.A(new_n670), .B(new_n674), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g474(.A1(new_n472), .A2(new_n475), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G15gat), .B1(new_n671), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(G15gat), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n298), .A2(new_n299), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n681), .ZN(G1326gat));
  NAND2_X1  g481(.A1(new_n665), .A2(new_n358), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT43), .B(G22gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  INV_X1    g484(.A(KEYINPUT45), .ZN(new_n686));
  INV_X1    g485(.A(new_n662), .ZN(new_n687));
  INV_X1    g486(.A(new_n618), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n644), .A2(new_n645), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n535), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n481), .A2(new_n687), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(G29gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n694), .A3(new_n666), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT101), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n695), .A2(KEYINPUT101), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n686), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n698), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(KEYINPUT45), .A3(new_n696), .ZN(new_n701));
  INV_X1    g500(.A(new_n692), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n476), .A2(KEYINPUT102), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n439), .A2(new_n705), .A3(new_n358), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n704), .A2(new_n706), .B1(new_n468), .B2(new_n458), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n707), .A2(new_n472), .A3(new_n475), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n703), .B(new_n662), .C1(new_n708), .C2(new_n444), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT103), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n680), .A2(new_n442), .A3(new_n428), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n443), .A2(KEYINPUT35), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n707), .A2(new_n472), .A3(new_n475), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n687), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n716), .A3(new_n703), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n477), .A2(KEYINPUT83), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n480), .A3(new_n469), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n713), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n703), .B1(new_n721), .B2(new_n662), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n702), .B1(new_n718), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723), .B2(new_n438), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n699), .A2(new_n701), .A3(new_n724), .ZN(G1328gat));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n672), .A2(G36gat), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n721), .A2(new_n662), .A3(new_n702), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT104), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n687), .B1(new_n720), .B2(new_n713), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n730), .A2(new_n731), .A3(new_n702), .A4(new_n727), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n729), .A2(KEYINPUT46), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT44), .B1(new_n481), .B2(new_n687), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n710), .A2(new_n717), .ZN(new_n735));
  AOI211_X1 g534(.A(new_n672), .B(new_n692), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(G36gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n733), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT46), .B1(new_n729), .B2(new_n732), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n726), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n739), .ZN(new_n741));
  OAI21_X1  g540(.A(G36gat), .B1(new_n723), .B2(new_n672), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n741), .A2(new_n742), .A3(KEYINPUT105), .A4(new_n733), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(G1329gat));
  NOR2_X1   g543(.A1(new_n481), .A2(new_n535), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n745), .A2(new_n680), .A3(new_n662), .A4(new_n690), .ZN(new_n746));
  INV_X1    g545(.A(G43gat), .ZN(new_n747));
  AOI22_X1  g546(.A1(new_n746), .A2(new_n747), .B1(KEYINPUT106), .B2(KEYINPUT47), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n677), .A2(new_n747), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n702), .B(new_n749), .C1(new_n718), .C2(new_n722), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  OR2_X1    g550(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1330gat));
  NAND2_X1  g552(.A1(new_n358), .A2(G50gat), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n693), .A2(new_n358), .ZN(new_n755));
  OAI22_X1  g554(.A1(new_n723), .A2(new_n754), .B1(new_n755), .B2(G50gat), .ZN(new_n756));
  XNOR2_X1  g555(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n756), .B(new_n758), .ZN(G1331gat));
  NAND2_X1  g558(.A1(new_n713), .A2(new_n714), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n688), .A2(new_n535), .A3(new_n663), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n666), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g563(.A(new_n391), .B(KEYINPUT108), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  AND2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n767), .B2(new_n768), .ZN(G1333gat));
  AOI21_X1  g570(.A(new_n554), .B1(new_n762), .B2(new_n676), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n298), .A2(new_n299), .A3(G71gat), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(new_n762), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n762), .A2(new_n358), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g576(.A1(new_n689), .A2(new_n691), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT109), .Z(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n715), .A2(KEYINPUT51), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT51), .B1(new_n715), .B2(new_n780), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n783), .A2(new_n688), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(new_n566), .A3(new_n666), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n779), .A2(new_n618), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n734), .B2(new_n735), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G85gat), .B1(new_n789), .B2(new_n438), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n785), .A2(new_n790), .ZN(G1336gat));
  AOI21_X1  g590(.A(new_n567), .B1(new_n788), .B2(new_n391), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n766), .A2(new_n567), .A3(new_n688), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT110), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n781), .B2(new_n782), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT52), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n766), .B(new_n786), .C1(new_n718), .C2(new_n722), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G92gat), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT111), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n804), .B(new_n801), .C1(new_n798), .C2(G92gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n797), .B1(new_n803), .B2(new_n805), .ZN(G1337gat));
  XNOR2_X1  g605(.A(KEYINPUT112), .B(G99gat), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n784), .A2(new_n680), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n789), .A2(new_n677), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n807), .ZN(G1338gat));
  INV_X1    g609(.A(G106gat), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n788), .B2(new_n358), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n442), .A2(G106gat), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n783), .A2(new_n688), .A3(new_n813), .ZN(new_n814));
  OR3_X1    g613(.A1(new_n812), .A2(new_n814), .A3(KEYINPUT53), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT53), .B1(new_n812), .B2(new_n814), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1339gat));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n533), .A2(new_n517), .A3(new_n531), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n522), .A2(new_n524), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n515), .B1(new_n513), .B2(new_n516), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n530), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n613), .B2(new_n617), .ZN(new_n825));
  INV_X1    g624(.A(new_n534), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n609), .B2(new_n610), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n597), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g628(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n596), .B(new_n830), .C1(new_n582), .C2(new_n585), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(new_n602), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n826), .A2(new_n819), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n602), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n835), .B1(new_n828), .B2(new_n597), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT114), .B1(new_n836), .B2(KEYINPUT55), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(KEYINPUT114), .A3(KEYINPUT55), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n834), .A2(new_n608), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n662), .B1(new_n825), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n608), .A3(new_n839), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n824), .B(new_n662), .C1(KEYINPUT55), .C2(new_n836), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n818), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n689), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT100), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n823), .B1(new_n849), .B2(new_n616), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n839), .A2(new_n608), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n532), .A2(new_n534), .B1(new_n836), .B2(KEYINPUT55), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n851), .A2(new_n852), .A3(new_n837), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n687), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n844), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(KEYINPUT115), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n845), .A2(new_n846), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n618), .A2(new_n663), .A3(new_n535), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n666), .A3(new_n359), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n765), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n862), .A2(new_n249), .A3(new_n535), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n860), .A2(KEYINPUT116), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(KEYINPUT116), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n691), .A3(new_n765), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n863), .B1(new_n867), .B2(new_n249), .ZN(G1340gat));
  OAI21_X1  g667(.A(G120gat), .B1(new_n862), .B2(new_n618), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n765), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n618), .A2(G120gat), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT117), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n869), .B1(new_n870), .B2(new_n872), .ZN(G1341gat));
  NOR3_X1   g672(.A1(new_n862), .A2(new_n244), .A3(new_n846), .ZN(new_n874));
  AOI211_X1 g673(.A(new_n846), .B(new_n766), .C1(new_n864), .C2(new_n865), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n876));
  AOI21_X1  g675(.A(G127gat), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT118), .B1(new_n870), .B2(new_n846), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(G1342gat));
  NAND2_X1  g678(.A1(new_n672), .A2(new_n662), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n880), .B(KEYINPUT119), .Z(new_n881));
  AOI211_X1 g680(.A(G134gat), .B(new_n881), .C1(new_n864), .C2(new_n865), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT56), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n861), .A2(new_n662), .A3(new_n765), .ZN(new_n884));
  AOI22_X1  g683(.A1(new_n882), .A2(new_n883), .B1(G134gat), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n881), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n866), .A2(new_n242), .A3(new_n886), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n887), .A2(KEYINPUT120), .A3(KEYINPUT56), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT120), .B1(new_n887), .B2(KEYINPUT56), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(G1343gat));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n442), .B1(new_n857), .B2(new_n858), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(KEYINPUT57), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  INV_X1    g693(.A(new_n858), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n854), .A2(new_n855), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n689), .B1(new_n896), .B2(new_n818), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n897), .B2(new_n856), .ZN(new_n898));
  OAI211_X1 g697(.A(KEYINPUT121), .B(new_n894), .C1(new_n898), .C2(new_n442), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n442), .A2(new_n894), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n841), .A2(new_n844), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n689), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n900), .B1(new_n902), .B2(new_n895), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n893), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n676), .A2(new_n438), .A3(new_n766), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n691), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G141gat), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n892), .A2(new_n905), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n317), .A3(new_n691), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT58), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n907), .A2(new_n912), .A3(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1344gat));
  NOR2_X1   g713(.A1(new_n318), .A2(KEYINPUT59), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n904), .A2(new_n905), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(new_n618), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n858), .B(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n358), .B1(new_n902), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n894), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n859), .A2(new_n900), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n923), .A2(new_n688), .A3(new_n905), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT59), .B1(new_n924), .B2(new_n318), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n917), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n908), .A2(new_n318), .A3(new_n688), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1345gat));
  OAI21_X1  g727(.A(G155gat), .B1(new_n916), .B2(new_n846), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n908), .A2(new_n632), .A3(new_n689), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1346gat));
  OAI21_X1  g730(.A(G162gat), .B1(new_n916), .B2(new_n687), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n881), .A2(G162gat), .A3(new_n438), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n892), .A2(new_n677), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1347gat));
  NOR2_X1   g734(.A1(new_n898), .A2(new_n666), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n359), .A2(new_n766), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT123), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(G169gat), .B1(new_n940), .B2(new_n691), .ZN(new_n941));
  INV_X1    g740(.A(new_n359), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n898), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n672), .A2(new_n666), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(KEYINPUT124), .A3(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT124), .B1(new_n943), .B2(new_n944), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n691), .A2(G169gat), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n941), .B1(new_n948), .B2(new_n949), .ZN(G1348gat));
  INV_X1    g749(.A(G176gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n940), .A2(new_n951), .A3(new_n688), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n946), .A2(new_n947), .A3(new_n618), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n953), .B2(new_n951), .ZN(G1349gat));
  INV_X1    g753(.A(G183gat), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n955), .B1(new_n948), .B2(new_n689), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n689), .A2(new_n209), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n939), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT60), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT60), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n946), .A2(new_n947), .A3(new_n846), .ZN(new_n961));
  OAI221_X1 g760(.A(new_n960), .B1(new_n939), .B2(new_n957), .C1(new_n961), .C2(new_n955), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n959), .A2(new_n962), .ZN(G1350gat));
  NAND3_X1  g762(.A1(new_n940), .A2(new_n210), .A3(new_n662), .ZN(new_n964));
  INV_X1    g763(.A(new_n947), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n965), .A2(new_n662), .A3(new_n945), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n966), .A2(new_n967), .A3(G190gat), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n967), .B1(new_n966), .B2(G190gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(G1351gat));
  AND2_X1   g769(.A1(new_n859), .A2(new_n900), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n858), .B(KEYINPUT122), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n972), .B1(new_n689), .B2(new_n901), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT57), .B1(new_n973), .B2(new_n358), .ZN(new_n974));
  OAI21_X1  g773(.A(KEYINPUT125), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n676), .A2(new_n666), .A3(new_n672), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n921), .A2(new_n922), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(G197gat), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n979), .A2(new_n980), .A3(new_n535), .ZN(new_n981));
  AND4_X1   g780(.A1(new_n358), .A2(new_n936), .A3(new_n677), .A4(new_n766), .ZN(new_n982));
  AOI21_X1  g781(.A(G197gat), .B1(new_n982), .B2(new_n691), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n981), .A2(new_n983), .ZN(G1352gat));
  XNOR2_X1  g783(.A(KEYINPUT126), .B(G204gat), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n618), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT62), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n987), .B(new_n988), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n985), .B1(new_n979), .B2(new_n618), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1353gat));
  NAND3_X1  g790(.A1(new_n923), .A2(new_n689), .A3(new_n976), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(G211gat), .ZN(new_n993));
  XOR2_X1   g792(.A(new_n993), .B(KEYINPUT63), .Z(new_n994));
  NAND3_X1  g793(.A1(new_n982), .A2(new_n305), .A3(new_n689), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(G1354gat));
  NAND3_X1  g795(.A1(new_n982), .A2(new_n306), .A3(new_n662), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n975), .A2(new_n999), .A3(new_n976), .A4(new_n978), .ZN(new_n1000));
  AND3_X1   g799(.A1(new_n998), .A2(new_n662), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n997), .B1(new_n1001), .B2(new_n306), .ZN(G1355gat));
endmodule


