//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT75), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(G211gat), .A2(G218gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G211gat), .A2(G218gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT71), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G211gat), .ZN(new_n210));
  INV_X1    g009(.A(G218gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT71), .ZN(new_n213));
  NAND2_X1  g012(.A1(G211gat), .A2(G218gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(KEYINPUT70), .A2(KEYINPUT22), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT70), .A2(KEYINPUT22), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n214), .A3(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G197gat), .B(G204gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n209), .A2(new_n219), .A3(new_n215), .A4(new_n220), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G183gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT27), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT27), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT28), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT27), .B(G183gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(KEYINPUT28), .A3(new_n230), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT65), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(new_n241), .A3(new_n238), .ZN(new_n242));
  NOR2_X1   g041(.A1(G169gat), .A2(G176gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT26), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n240), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G183gat), .A2(G190gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n236), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n250));
  AND2_X1   g049(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n247), .A2(new_n250), .B1(new_n251), .B2(G190gat), .ZN(new_n252));
  INV_X1    g051(.A(G169gat), .ZN(new_n253));
  INV_X1    g052(.A(G176gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT23), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT23), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(G169gat), .B2(G176gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n257), .A3(new_n238), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n249), .B1(new_n252), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n250), .A2(new_n247), .ZN(new_n260));
  NAND3_X1  g059(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n253), .A2(new_n254), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n263), .A2(new_n256), .B1(KEYINPUT64), .B2(new_n238), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n249), .B1(new_n243), .B2(KEYINPUT23), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n238), .A2(KEYINPUT64), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n262), .A2(new_n264), .A3(new_n265), .A4(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n248), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT29), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n248), .A2(new_n268), .A3(KEYINPUT72), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT73), .ZN(new_n275));
  NAND2_X1  g074(.A1(G226gat), .A2(G233gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n269), .A2(G226gat), .A3(G233gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n275), .B1(new_n274), .B2(new_n276), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n225), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n269), .A2(new_n272), .A3(new_n276), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n271), .A2(new_n273), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(new_n276), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n224), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT74), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n281), .A2(new_n288), .A3(new_n285), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n206), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n281), .A2(new_n206), .A3(new_n285), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT30), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n281), .A2(KEYINPUT30), .A3(new_n206), .A4(new_n285), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G1gat), .B(G29gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT0), .ZN(new_n297));
  XNOR2_X1  g096(.A(G57gat), .B(G85gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G225gat), .A2(G233gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT2), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT78), .ZN(new_n306));
  AND2_X1   g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(G141gat), .A2(G148gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G141gat), .ZN(new_n310));
  INV_X1    g109(.A(G148gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(KEYINPUT78), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n305), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G155gat), .ZN(new_n316));
  INV_X1    g115(.A(G162gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT77), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT77), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(G155gat), .B2(G162gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n303), .A2(KEYINPUT76), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT76), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(G155gat), .A3(G162gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT2), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT79), .B(G155gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT80), .B(G162gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n316), .A2(new_n317), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n303), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(new_n312), .A3(new_n313), .ZN(new_n333));
  OAI22_X1  g132(.A1(new_n315), .A2(new_n326), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G113gat), .ZN(new_n335));
  INV_X1    g134(.A(G120gat), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT1), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G134gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G127gat), .ZN(new_n339));
  INV_X1    g138(.A(G127gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G134gat), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n337), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT66), .B(G113gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G120gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n337), .B1(new_n335), .B2(new_n336), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n339), .A2(new_n341), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n334), .A2(new_n349), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n342), .A2(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n307), .A2(new_n308), .A3(new_n306), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT78), .B1(new_n312), .B2(new_n313), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n304), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n326), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n328), .A2(new_n329), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT2), .ZN(new_n358));
  AOI211_X1 g157(.A(new_n308), .B(new_n307), .C1(new_n303), .C2(new_n331), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n351), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n302), .B1(new_n350), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n356), .A2(new_n360), .A3(new_n351), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT82), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n354), .A2(new_n355), .B1(new_n358), .B2(new_n359), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n369), .A2(new_n370), .A3(new_n366), .A4(new_n351), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT4), .B1(new_n334), .B2(new_n349), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n368), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(new_n334), .B2(KEYINPUT3), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT3), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n356), .A2(new_n360), .A3(KEYINPUT81), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n351), .B1(new_n334), .B2(KEYINPUT3), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n302), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n365), .B1(new_n373), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n379), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n372), .A2(new_n367), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n364), .A2(new_n302), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n300), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n382), .A2(new_n373), .A3(new_n301), .ZN(new_n388));
  INV_X1    g187(.A(new_n365), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(new_n299), .A3(new_n385), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT6), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n387), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(KEYINPUT6), .B(new_n300), .C1(new_n381), .C2(new_n386), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n290), .A2(new_n295), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n222), .A2(new_n272), .A3(new_n223), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n397), .A2(new_n376), .B1(new_n356), .B2(new_n360), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT29), .B1(new_n375), .B2(new_n377), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(new_n224), .ZN(new_n401));
  OAI211_X1 g200(.A(G228gat), .B(G233gat), .C1(new_n398), .C2(KEYINPUT84), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n402), .B(new_n399), .C1(new_n224), .C2(new_n400), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(G22gat), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT85), .ZN(new_n407));
  XOR2_X1   g206(.A(G78gat), .B(G106gat), .Z(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT31), .B(G50gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n404), .A2(new_n405), .ZN(new_n412));
  INV_X1    g211(.A(G22gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n406), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n407), .A2(new_n414), .A3(new_n406), .A4(new_n410), .ZN(new_n417));
  XOR2_X1   g216(.A(G15gat), .B(G43gat), .Z(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT67), .ZN(new_n419));
  XNOR2_X1  g218(.A(G71gat), .B(G99gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n269), .A2(new_n351), .ZN(new_n422));
  NAND2_X1  g221(.A1(G227gat), .A2(G233gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n248), .A2(new_n268), .A3(new_n349), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n422), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT33), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n421), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(KEYINPUT32), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n426), .B(KEYINPUT32), .C1(new_n427), .C2(new_n421), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n248), .A2(new_n268), .A3(new_n349), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n349), .B1(new_n248), .B2(new_n268), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n423), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT68), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n436), .A2(KEYINPUT34), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(KEYINPUT34), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n425), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n440), .A2(new_n436), .A3(KEYINPUT34), .A4(new_n423), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n432), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT69), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n430), .A2(new_n442), .A3(new_n431), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT69), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n442), .B1(new_n430), .B2(new_n431), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n416), .A2(new_n417), .A3(new_n445), .A4(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT90), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n448), .A2(new_n447), .ZN(new_n453));
  INV_X1    g252(.A(new_n446), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n445), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n455), .A2(KEYINPUT90), .A3(new_n417), .A4(new_n416), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n396), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT35), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT91), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT91), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n460), .A3(KEYINPUT35), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT35), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n416), .A2(new_n417), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n446), .A2(new_n448), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n396), .A2(new_n462), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n459), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n445), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT36), .ZN(new_n469));
  INV_X1    g268(.A(new_n465), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n470), .A2(KEYINPUT36), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n463), .B(KEYINPUT86), .ZN(new_n473));
  INV_X1    g272(.A(new_n396), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n476), .B1(new_n287), .B2(new_n289), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n205), .B1(new_n286), .B2(KEYINPUT37), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT38), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT89), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g280(.A(KEYINPUT89), .B(KEYINPUT38), .C1(new_n477), .C2(new_n478), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n478), .A2(KEYINPUT38), .ZN(new_n483));
  OR3_X1    g282(.A1(new_n279), .A2(new_n225), .A3(new_n280), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT88), .ZN(new_n485));
  OR4_X1    g284(.A1(KEYINPUT88), .A2(new_n279), .A3(new_n225), .A4(new_n280), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n284), .A2(new_n224), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n483), .B1(new_n488), .B2(new_n476), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n395), .A2(new_n291), .ZN(new_n490));
  AND4_X1   g289(.A1(new_n481), .A2(new_n482), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n382), .A2(new_n383), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT39), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n493), .A3(new_n302), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n494), .A2(new_n299), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n302), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n350), .A2(new_n361), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n496), .B(KEYINPUT39), .C1(new_n302), .C2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(new_n498), .A3(KEYINPUT40), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n387), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT40), .B1(new_n495), .B2(new_n498), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(new_n290), .B2(new_n295), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n463), .B1(new_n503), .B2(KEYINPUT87), .ZN(new_n504));
  INV_X1    g303(.A(new_n290), .ZN(new_n505));
  INV_X1    g304(.A(new_n295), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT87), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n508), .A3(new_n502), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n475), .B1(new_n491), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n467), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT16), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(G1gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(G1gat), .B2(new_n513), .ZN(new_n516));
  INV_X1    g315(.A(G8gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(KEYINPUT94), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT93), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n522), .A2(KEYINPUT15), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n521), .B(new_n523), .ZN(new_n524));
  NOR3_X1   g323(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT95), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n527), .A2(new_n528), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G29gat), .A2(G36gat), .ZN(new_n531));
  INV_X1    g330(.A(new_n528), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n531), .B1(new_n532), .B2(new_n525), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n524), .A2(new_n522), .A3(new_n529), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n519), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT96), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n538), .A2(new_n543), .A3(KEYINPUT17), .A4(new_n539), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n533), .B1(new_n524), .B2(new_n529), .ZN(new_n545));
  OAI211_X1 g344(.A(KEYINPUT17), .B(new_n539), .C1(new_n545), .C2(new_n536), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT96), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n542), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n540), .A2(new_n519), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n549), .A2(KEYINPUT18), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n530), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n535), .A2(new_n537), .B1(new_n553), .B2(new_n522), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n518), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n551), .A2(KEYINPUT97), .A3(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n550), .B(KEYINPUT13), .Z(new_n557));
  INV_X1    g356(.A(KEYINPUT97), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n558), .A3(new_n519), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n552), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n554), .A2(new_n518), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(new_n542), .B2(new_n548), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT18), .B1(new_n563), .B2(new_n550), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G169gat), .B(G197gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT12), .Z(new_n571));
  AOI21_X1  g370(.A(KEYINPUT98), .B1(new_n565), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT98), .ZN(new_n573));
  INV_X1    g372(.A(new_n571), .ZN(new_n574));
  NOR4_X1   g373(.A1(new_n561), .A2(new_n564), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  OAI22_X1  g374(.A1(new_n572), .A2(new_n575), .B1(new_n565), .B2(new_n571), .ZN(new_n576));
  XOR2_X1   g375(.A(G99gat), .B(G106gat), .Z(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT102), .B(KEYINPUT7), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(G85gat), .A3(G92gat), .ZN(new_n579));
  OR2_X1    g378(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n580));
  NAND2_X1  g379(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n581));
  INV_X1    g380(.A(G85gat), .ZN(new_n582));
  INV_X1    g381(.A(G92gat), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT8), .A2(new_n585), .B1(new_n582), .B2(new_n583), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n579), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT103), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT103), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n579), .A2(new_n589), .A3(new_n584), .A4(new_n586), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n577), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n577), .A3(new_n590), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n540), .A2(new_n594), .B1(KEYINPUT41), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n594), .B1(new_n540), .B2(new_n541), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT104), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n597), .A2(new_n548), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n597), .B2(new_n548), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G190gat), .B(G218gat), .Z(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n602), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n604), .B(new_n596), .C1(new_n599), .C2(new_n600), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n595), .A2(KEYINPUT41), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT101), .ZN(new_n608));
  XNOR2_X1  g407(.A(G134gat), .B(G162gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n606), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G57gat), .B(G64gat), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G71gat), .B(G78gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT99), .B(KEYINPUT21), .Z(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G127gat), .B(G155gat), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n620), .B(new_n621), .Z(new_n622));
  AOI21_X1  g421(.A(new_n519), .B1(KEYINPUT21), .B2(new_n617), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT100), .ZN(new_n626));
  XOR2_X1   g425(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G183gat), .B(G211gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n624), .B(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n612), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n593), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n617), .B1(new_n636), .B2(new_n591), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n592), .A2(new_n618), .A3(new_n593), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n594), .A2(KEYINPUT10), .A3(new_n617), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n635), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT105), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n634), .B1(new_n637), .B2(new_n638), .ZN(new_n644));
  XNOR2_X1  g443(.A(G120gat), .B(G148gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n642), .B2(new_n644), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n633), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n512), .A2(new_n576), .A3(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n654), .A2(KEYINPUT106), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(KEYINPUT106), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n395), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g458(.A(new_n517), .B1(new_n657), .B2(new_n507), .ZN(new_n660));
  INV_X1    g459(.A(new_n507), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT16), .B(G8gat), .Z(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AOI211_X1 g462(.A(new_n661), .B(new_n663), .C1(new_n655), .C2(new_n656), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT42), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n657), .A2(new_n507), .A3(new_n662), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(G1325gat));
  INV_X1    g468(.A(G15gat), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n657), .A2(new_n670), .A3(new_n465), .ZN(new_n671));
  INV_X1    g470(.A(new_n472), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n655), .B2(new_n656), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n673), .B2(new_n670), .ZN(G1326gat));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n473), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT43), .B(G22gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  AOI21_X1  g476(.A(new_n460), .B1(new_n457), .B2(KEYINPUT35), .ZN(new_n678));
  INV_X1    g477(.A(new_n466), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n481), .A2(new_n482), .A3(new_n489), .A4(new_n490), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(new_n509), .A3(new_n504), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n680), .A2(new_n461), .B1(new_n682), .B2(new_n475), .ZN(new_n683));
  INV_X1    g482(.A(new_n652), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n612), .A2(new_n631), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT107), .ZN(new_n686));
  INV_X1    g485(.A(new_n561), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n563), .A2(new_n550), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT18), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n571), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n690), .A2(new_n552), .A3(new_n560), .A4(new_n571), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n573), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n565), .A2(KEYINPUT98), .A3(new_n571), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OR3_X1    g494(.A1(new_n683), .A2(new_n686), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n395), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n696), .A2(G29gat), .A3(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT45), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n606), .B(new_n610), .ZN(new_n700));
  OAI22_X1  g499(.A1(new_n683), .A2(new_n700), .B1(KEYINPUT109), .B2(KEYINPUT44), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n512), .A2(new_n612), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n652), .B(KEYINPUT108), .ZN(new_n706));
  INV_X1    g505(.A(new_n631), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n706), .A2(new_n695), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(KEYINPUT110), .A3(new_n395), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n709), .B2(new_n697), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(G29gat), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n714), .ZN(G1328gat));
  NOR3_X1   g514(.A1(new_n696), .A2(G36gat), .A3(new_n661), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT46), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT111), .B1(new_n709), .B2(new_n661), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G36gat), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n709), .A2(KEYINPUT111), .A3(new_n661), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n717), .B1(new_n719), .B2(new_n720), .ZN(G1329gat));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n472), .A3(new_n708), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n683), .A2(new_n686), .A3(new_n695), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n470), .A2(G43gat), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n722), .A2(G43gat), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g525(.A(G50gat), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n710), .B2(new_n463), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n723), .A2(KEYINPUT112), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT86), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n463), .B(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(G50gat), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n733), .B1(new_n723), .B2(KEYINPUT112), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT48), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n705), .A2(new_n473), .A3(new_n708), .ZN(new_n737));
  AOI22_X1  g536(.A1(new_n737), .A2(G50gat), .B1(new_n729), .B2(new_n734), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n728), .A2(new_n736), .B1(new_n738), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g538(.A1(new_n632), .A2(new_n695), .A3(new_n706), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT113), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n512), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n395), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g544(.A(new_n661), .B(new_n742), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1333gat));
  NOR3_X1   g547(.A1(new_n742), .A2(G71gat), .A3(new_n470), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n743), .A2(new_n472), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(G71gat), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n743), .A2(new_n473), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g553(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n755), .B1(new_n512), .B2(new_n612), .ZN(new_n756));
  AOI211_X1 g555(.A(new_n700), .B(new_n702), .C1(new_n467), .C2(new_n511), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n695), .A2(new_n631), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT114), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n652), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n758), .A2(new_n697), .A3(new_n761), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n457), .A2(new_n460), .A3(KEYINPUT35), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n763), .A2(new_n678), .A3(new_n679), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n672), .B1(new_n731), .B2(new_n396), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n504), .A2(new_n509), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n766), .B2(new_n681), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n612), .B(new_n760), .C1(new_n764), .C2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n512), .A2(KEYINPUT51), .A3(new_n612), .A4(new_n760), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n652), .A2(new_n582), .A3(new_n395), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n762), .A2(new_n582), .B1(new_n773), .B2(new_n774), .ZN(G1336gat));
  NAND4_X1  g574(.A1(new_n772), .A2(new_n583), .A3(new_n507), .A4(new_n706), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n758), .A2(new_n661), .A3(new_n761), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(new_n583), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT52), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n780), .B(new_n776), .C1(new_n777), .C2(new_n583), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(G1337gat));
  NOR3_X1   g581(.A1(new_n758), .A2(new_n672), .A3(new_n761), .ZN(new_n783));
  INV_X1    g582(.A(G99gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n652), .A2(new_n784), .A3(new_n465), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n783), .A2(new_n784), .B1(new_n773), .B2(new_n785), .ZN(G1338gat));
  INV_X1    g585(.A(new_n761), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n473), .B(new_n787), .C1(new_n756), .C2(new_n757), .ZN(new_n788));
  INV_X1    g587(.A(new_n706), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n789), .A2(G106gat), .A3(new_n464), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n788), .A2(G106gat), .B1(new_n772), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT115), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794));
  INV_X1    g593(.A(G106gat), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n761), .B1(new_n701), .B2(new_n704), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(new_n473), .ZN(new_n797));
  INV_X1    g596(.A(new_n790), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n770), .B2(new_n771), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n794), .B(KEYINPUT53), .C1(new_n797), .C2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT53), .B1(new_n772), .B2(new_n790), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n463), .B(new_n787), .C1(new_n756), .C2(new_n757), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G106gat), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n801), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n801), .B2(new_n803), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n793), .B(new_n800), .C1(new_n805), .C2(new_n806), .ZN(G1339gat));
  INV_X1    g606(.A(new_n642), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT105), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n640), .A2(new_n641), .A3(new_n635), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(KEYINPUT54), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT105), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n642), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n809), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n647), .B1(new_n642), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n817), .A2(new_n818), .B1(new_n643), .B2(new_n649), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820));
  INV_X1    g619(.A(new_n816), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n643), .B2(new_n811), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n820), .B1(new_n822), .B2(KEYINPUT55), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n814), .A2(new_n816), .A3(KEYINPUT55), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(KEYINPUT117), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n819), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n695), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n556), .A2(new_n559), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n828), .A2(new_n557), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n563), .A2(new_n550), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n570), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n831), .B(new_n684), .C1(new_n693), .C2(new_n694), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n700), .B1(new_n827), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n650), .B1(new_n822), .B2(KEYINPUT55), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n824), .A2(KEYINPUT117), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n822), .A2(new_n820), .A3(KEYINPUT55), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n831), .B1(new_n693), .B2(new_n694), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n612), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n707), .B1(new_n833), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n700), .A2(new_n695), .A3(new_n707), .A4(new_n684), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n697), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n452), .A2(new_n456), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n507), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n695), .A2(new_n343), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n731), .A2(new_n465), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n507), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n844), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n695), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT118), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n849), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(G1340gat));
  AOI21_X1  g657(.A(G120gat), .B1(new_n847), .B2(new_n652), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n852), .A2(new_n336), .A3(new_n789), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(G1341gat));
  NAND3_X1  g660(.A1(new_n847), .A2(new_n340), .A3(new_n707), .ZN(new_n862));
  OAI21_X1  g661(.A(G127gat), .B1(new_n852), .B2(new_n631), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1342gat));
  AND4_X1   g663(.A1(new_n338), .A2(new_n844), .A3(new_n612), .A4(new_n846), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT56), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(G134gat), .B1(new_n852), .B2(new_n700), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n865), .A2(new_n869), .A3(new_n866), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n865), .B2(new_n866), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n867), .B(new_n868), .C1(new_n870), .C2(new_n871), .ZN(G1343gat));
  NOR3_X1   g671(.A1(new_n472), .A2(new_n507), .A3(new_n697), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n878), .B1(new_n843), .B2(new_n464), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n837), .A2(new_n576), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n838), .A2(new_n652), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n612), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n839), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n631), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n841), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n731), .A2(new_n878), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n877), .B1(new_n879), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n310), .B1(new_n888), .B2(new_n576), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n672), .A2(new_n463), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n507), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n844), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n576), .A2(new_n310), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT58), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n877), .ZN(new_n896));
  INV_X1    g695(.A(new_n887), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT57), .B1(new_n885), .B2(new_n463), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G141gat), .B1(new_n899), .B2(new_n695), .ZN(new_n900));
  INV_X1    g699(.A(new_n894), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT58), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n895), .A2(new_n903), .ZN(G1344gat));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n905), .B(G148gat), .C1(new_n899), .C2(new_n684), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n731), .A2(KEYINPUT57), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n632), .A2(KEYINPUT121), .A3(new_n695), .A4(new_n684), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n841), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n908), .B1(new_n840), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n877), .A2(new_n684), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n464), .B1(new_n884), .B2(new_n841), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n913), .B(new_n914), .C1(new_n915), .C2(new_n878), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G148gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n907), .B1(new_n917), .B2(KEYINPUT59), .ZN(new_n918));
  AOI211_X1 g717(.A(KEYINPUT122), .B(new_n905), .C1(new_n916), .C2(G148gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n906), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n892), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n311), .A3(new_n652), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1345gat));
  AOI21_X1  g722(.A(new_n328), .B1(new_n921), .B2(new_n707), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n707), .A2(new_n328), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT123), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n924), .B1(new_n888), .B2(new_n926), .ZN(G1346gat));
  OR3_X1    g726(.A1(new_n892), .A2(new_n329), .A3(new_n700), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n888), .A2(KEYINPUT124), .A3(new_n612), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n329), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT124), .B1(new_n888), .B2(new_n612), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1347gat));
  NAND2_X1  g731(.A1(new_n507), .A2(new_n697), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n850), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n885), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n935), .A2(new_n253), .A3(new_n695), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n843), .A2(new_n395), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n845), .A2(new_n661), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n939), .A2(KEYINPUT125), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(KEYINPUT125), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n940), .A2(new_n576), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n936), .B1(new_n942), .B2(new_n253), .ZN(G1348gat));
  OAI21_X1  g742(.A(G176gat), .B1(new_n935), .B2(new_n789), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n940), .A2(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n652), .A2(new_n254), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(G1349gat));
  OAI21_X1  g746(.A(G183gat), .B1(new_n935), .B2(new_n631), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n707), .A2(new_n234), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n939), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g750(.A(G190gat), .B1(new_n935), .B2(new_n700), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n952), .A2(KEYINPUT126), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(KEYINPUT126), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(KEYINPUT61), .A3(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n952), .A2(KEYINPUT126), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n612), .A2(new_n230), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n955), .B(new_n957), .C1(new_n945), .C2(new_n958), .ZN(G1351gat));
  NOR2_X1   g758(.A1(new_n890), .A2(new_n661), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n695), .A2(G197gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n937), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT127), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT57), .B1(new_n843), .B2(new_n464), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n933), .A2(new_n472), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(new_n913), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(G197gat), .B1(new_n966), .B2(new_n695), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n963), .A2(new_n967), .ZN(G1352gat));
  NOR2_X1   g767(.A1(new_n684), .A2(G204gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n937), .A2(new_n960), .A3(new_n969), .ZN(new_n970));
  XOR2_X1   g769(.A(new_n970), .B(KEYINPUT62), .Z(new_n971));
  OAI21_X1  g770(.A(G204gat), .B1(new_n966), .B2(new_n789), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1353gat));
  AND2_X1   g772(.A1(new_n937), .A2(new_n960), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n974), .A2(new_n210), .A3(new_n707), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n964), .A2(new_n707), .A3(new_n913), .A4(new_n965), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n976), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT63), .B1(new_n976), .B2(G211gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(G1354gat));
  OAI21_X1  g778(.A(G218gat), .B1(new_n966), .B2(new_n700), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n974), .A2(new_n211), .A3(new_n612), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1355gat));
endmodule


