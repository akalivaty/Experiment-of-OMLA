//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n566,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  XNOR2_X1  g032(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n463), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n472), .A2(KEYINPUT69), .A3(G137), .A4(new_n469), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n465), .A2(G2105), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n471), .A2(new_n473), .B1(G101), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n477), .B1(new_n466), .B2(new_n467), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n472), .A2(new_n479), .A3(G125), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(G2105), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n475), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  AND2_X1   g060(.A1(new_n472), .A2(KEYINPUT70), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n472), .A2(KEYINPUT70), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n469), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  OAI21_X1  g065(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n469), .A2(G112), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n490), .B(new_n493), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n496), .B(new_n497), .ZN(G162));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n472), .A2(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(new_n469), .A2(G114), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n469), .A2(G138), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT4), .B1(new_n468), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n472), .A2(new_n508), .A3(G138), .A4(new_n469), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(new_n507), .B2(new_n509), .ZN(G164));
  NAND2_X1  g085(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(KEYINPUT73), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n514), .B1(KEYINPUT72), .B2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  OAI21_X1  g091(.A(G543), .B1(new_n516), .B2(KEYINPUT73), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n513), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(new_n512), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G50), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n522), .A2(new_n523), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n518), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G88), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n521), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  NAND3_X1  g107(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT74), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n518), .A2(new_n535), .A3(G63), .A4(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  OAI211_X1 g114(.A(G51), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n511), .A2(KEYINPUT73), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n542), .A2(G543), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n524), .B1(new_n544), .B2(new_n513), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n541), .B1(G89), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n537), .A2(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  AOI22_X1  g123(.A1(new_n545), .A2(G90), .B1(G52), .B2(new_n525), .ZN(new_n549));
  AND2_X1   g124(.A1(G77), .A2(G543), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n518), .B2(G64), .ZN(new_n551));
  OAI21_X1  g126(.A(G651), .B1(new_n551), .B2(KEYINPUT75), .ZN(new_n552));
  INV_X1    g127(.A(G64), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n544), .B2(new_n513), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n555));
  NOR3_X1   g130(.A1(new_n554), .A2(new_n555), .A3(new_n550), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n549), .B1(new_n552), .B2(new_n556), .ZN(G301));
  INV_X1    g132(.A(G301), .ZN(G171));
  NAND2_X1  g133(.A1(new_n525), .A2(G43), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n518), .A2(G81), .A3(new_n527), .ZN(new_n560));
  AND2_X1   g135(.A1(G68), .A2(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n518), .B2(G56), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n559), .B(new_n560), .C1(new_n562), .C2(new_n520), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n566), .B(KEYINPUT76), .Z(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n544), .B2(new_n513), .ZN(new_n572));
  AND2_X1   g147(.A1(G78), .A2(G543), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n527), .A2(KEYINPUT77), .A3(G53), .A4(G543), .ZN(new_n575));
  OAI211_X1 g150(.A(G53), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n575), .A2(KEYINPUT9), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n545), .A2(G91), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT9), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n576), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n574), .A2(new_n579), .A3(new_n580), .A4(new_n582), .ZN(G299));
  INV_X1    g158(.A(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n544), .A2(new_n584), .A3(new_n513), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(new_n525), .B2(G49), .ZN(new_n586));
  AOI21_X1  g161(.A(KEYINPUT78), .B1(new_n545), .B2(G87), .ZN(new_n587));
  AND4_X1   g162(.A1(KEYINPUT78), .A2(new_n518), .A3(G87), .A4(new_n527), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n525), .A2(G48), .ZN(new_n590));
  INV_X1    g165(.A(G86), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  OAI221_X1 g167(.A(new_n590), .B1(new_n528), .B2(new_n591), .C1(new_n592), .C2(new_n520), .ZN(G305));
  AOI22_X1  g168(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n520), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n525), .A2(G47), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n528), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n528), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n545), .A2(KEYINPUT10), .A3(G92), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n525), .A2(G54), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(new_n544), .B2(new_n513), .ZN(new_n609));
  AND2_X1   g184(.A1(G79), .A2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(G651), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n606), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n601), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n601), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  AND4_X1   g191(.A1(new_n574), .A2(new_n579), .A3(new_n580), .A4(new_n582), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(G868), .B2(new_n617), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(G868), .B2(new_n617), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n472), .A2(new_n474), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n630), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n631));
  INV_X1    g206(.A(G135), .ZN(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  OAI221_X1 g208(.A(new_n631), .B1(new_n488), .B2(new_n632), .C1(new_n633), .C2(new_n491), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(G2096), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n635), .A3(new_n636), .ZN(G156));
  XOR2_X1   g212(.A(KEYINPUT79), .B(KEYINPUT14), .Z(new_n638));
  XOR2_X1   g213(.A(KEYINPUT15), .B(G2435), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2438), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2430), .Z(new_n641));
  AOI21_X1  g216(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n640), .B2(new_n641), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n645), .B(new_n646), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(G14), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n650), .B2(new_n648), .ZN(G401));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT80), .ZN(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  XNOR2_X1  g230(.A(G2084), .B(G2090), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n655), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n655), .B(KEYINPUT17), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n659), .B(new_n656), .C1(new_n654), .C2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n656), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n660), .A2(new_n654), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n658), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2096), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT81), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n669), .A2(new_n674), .A3(new_n672), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n669), .A2(new_n674), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n677));
  AOI211_X1 g252(.A(new_n673), .B(new_n675), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(new_n676), .B2(new_n677), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT84), .Z(new_n680));
  XOR2_X1   g255(.A(G1991), .B(G1996), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT83), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n680), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G229));
  NOR2_X1   g263(.A1(G6), .A2(G16), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n592), .A2(new_n520), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n590), .B1(new_n528), .B2(new_n591), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n689), .B1(new_n692), .B2(G16), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT32), .B(G1981), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(KEYINPUT87), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(KEYINPUT87), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(G1971), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  AND3_X1   g277(.A1(new_n696), .A2(new_n697), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(G16), .A2(G23), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT88), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT78), .ZN(new_n706));
  INV_X1    g281(.A(G87), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n528), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n545), .A2(KEYINPUT78), .A3(G87), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n705), .B1(new_n710), .B2(new_n586), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n705), .B(new_n586), .C1(new_n587), .C2(new_n588), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n704), .B1(new_n714), .B2(G16), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT33), .B(G1976), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n703), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n703), .A2(KEYINPUT89), .A3(new_n717), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n720), .A2(KEYINPUT34), .A3(new_n721), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n698), .A2(G24), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n599), .B2(new_n698), .ZN(new_n727));
  INV_X1    g302(.A(G1986), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G25), .A2(G29), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n489), .A2(G131), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n492), .A2(G119), .ZN(new_n732));
  OR2_X1    g307(.A1(G95), .A2(G2105), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n733), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n734));
  AND3_X1   g309(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n730), .B1(new_n735), .B2(G29), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT85), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT35), .B(G1991), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n729), .B1(new_n739), .B2(KEYINPUT86), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(KEYINPUT86), .B2(new_n739), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n724), .A2(new_n725), .A3(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(KEYINPUT36), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT91), .Z(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n724), .A2(new_n741), .A3(new_n745), .A4(new_n725), .ZN(new_n748));
  INV_X1    g323(.A(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G32), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n489), .A2(G141), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n492), .A2(G129), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT26), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n755), .A2(new_n756), .B1(G105), .B2(new_n474), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n751), .A2(new_n752), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n750), .B1(new_n759), .B2(new_n749), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT27), .ZN(new_n761));
  INV_X1    g336(.A(G1996), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NOR2_X1   g339(.A1(G171), .A2(new_n698), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G5), .B2(new_n698), .ZN(new_n766));
  INV_X1    g341(.A(G1961), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT24), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n749), .B1(new_n769), .B2(G34), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n769), .B2(G34), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G160), .B2(G29), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G2084), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT94), .Z(new_n774));
  NAND4_X1  g349(.A1(new_n763), .A2(new_n764), .A3(new_n768), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n766), .A2(new_n767), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n749), .A2(G33), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT25), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n489), .B2(G139), .ZN(new_n780));
  NAND2_X1  g355(.A1(G115), .A2(G2104), .ZN(new_n781));
  INV_X1    g356(.A(G127), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n468), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n469), .B1(new_n783), .B2(KEYINPUT93), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(KEYINPUT93), .B2(new_n783), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n777), .B1(new_n786), .B2(G29), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n787), .A2(new_n442), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n442), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n749), .A2(G27), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G164), .B2(new_n749), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(new_n443), .ZN(new_n792));
  INV_X1    g367(.A(G28), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(KEYINPUT30), .ZN(new_n794));
  AOI21_X1  g369(.A(G29), .B1(new_n793), .B2(KEYINPUT30), .ZN(new_n795));
  OR2_X1    g370(.A1(KEYINPUT31), .A2(G11), .ZN(new_n796));
  NAND2_X1  g371(.A1(KEYINPUT31), .A2(G11), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n794), .A2(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n792), .B(new_n798), .C1(new_n749), .C2(new_n634), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n776), .A2(new_n788), .A3(new_n789), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n772), .A2(G2084), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(KEYINPUT95), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n698), .A2(G21), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G168), .B2(new_n698), .ZN(new_n804));
  INV_X1    g379(.A(G1966), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n801), .A2(KEYINPUT95), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n800), .A2(new_n802), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n775), .A2(new_n808), .A3(KEYINPUT96), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT96), .B1(new_n775), .B2(new_n808), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n749), .A2(G26), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT28), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n813));
  INV_X1    g388(.A(G116), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G2105), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n492), .B2(G128), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n489), .A2(G140), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G29), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n819), .A2(KEYINPUT92), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(KEYINPUT92), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n812), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(G2067), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(G2067), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n613), .A2(G16), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G4), .B2(G16), .ZN(new_n826));
  INV_X1    g401(.A(G1348), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n698), .A2(G19), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n564), .B2(new_n698), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(G1341), .Z(new_n831));
  NAND4_X1  g406(.A1(new_n823), .A2(new_n824), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(G29), .A2(G35), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(G162), .B2(G29), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT29), .B(G2090), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n698), .A2(G20), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT23), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n617), .B2(new_n698), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(G1956), .Z(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n827), .B2(new_n826), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n832), .A2(new_n836), .A3(new_n841), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n809), .A2(new_n810), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n747), .A2(new_n748), .A3(new_n843), .ZN(G150));
  INV_X1    g419(.A(G150), .ZN(G311));
  NAND2_X1  g420(.A1(new_n613), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n525), .A2(G55), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT97), .B(G93), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n518), .A2(new_n527), .A3(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(G80), .A2(G543), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n518), .B2(G67), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n848), .B(new_n850), .C1(new_n852), .C2(new_n520), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n563), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n560), .A2(new_n559), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n545), .A2(new_n849), .B1(G55), .B2(new_n525), .ZN(new_n856));
  INV_X1    g431(.A(G56), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(new_n544), .B2(new_n513), .ZN(new_n858));
  OAI21_X1  g433(.A(G651), .B1(new_n858), .B2(new_n561), .ZN(new_n859));
  INV_X1    g434(.A(G67), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(new_n544), .B2(new_n513), .ZN(new_n861));
  OAI21_X1  g436(.A(G651), .B1(new_n861), .B2(new_n851), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n855), .A2(new_n856), .A3(new_n859), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n854), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n847), .B(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT98), .ZN(new_n868));
  AOI21_X1  g443(.A(G860), .B1(new_n866), .B2(KEYINPUT39), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n853), .A2(G860), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT37), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(G145));
  OR2_X1    g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n874), .B(G2104), .C1(G118), .C2(new_n469), .ZN(new_n875));
  INV_X1    g450(.A(G142), .ZN(new_n876));
  INV_X1    g451(.A(G130), .ZN(new_n877));
  OAI221_X1 g452(.A(new_n875), .B1(new_n488), .B2(new_n876), .C1(new_n877), .C2(new_n491), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n627), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n879), .A2(new_n735), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n735), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n507), .A2(new_n509), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n505), .A2(new_n884), .ZN(new_n885));
  AOI22_X1  g460(.A1(new_n472), .A2(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT99), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n883), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n816), .B2(new_n817), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n816), .A2(new_n889), .A3(new_n817), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n758), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n759), .B1(new_n894), .B2(new_n890), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n786), .A2(KEYINPUT100), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n895), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n786), .B(KEYINPUT100), .Z(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n882), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n882), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n897), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n902), .B2(new_n903), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(G162), .B(new_n634), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n908), .A2(new_n484), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n484), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n909), .A2(new_n910), .B1(new_n901), .B2(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n901), .A2(new_n913), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n914), .B(new_n915), .C1(new_n906), .C2(new_n905), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT40), .ZN(G395));
  AND2_X1   g493(.A1(new_n611), .A2(new_n607), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n617), .B1(new_n606), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n612), .A2(G299), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT103), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n622), .B(new_n864), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n612), .A2(G299), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n617), .A2(new_n606), .A3(new_n919), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT41), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT41), .B1(new_n926), .B2(new_n927), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n925), .B1(new_n924), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT42), .ZN(new_n932));
  NAND2_X1  g507(.A1(G288), .A2(KEYINPUT88), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n933), .A2(new_n599), .A3(new_n712), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n599), .B1(new_n933), .B2(new_n712), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT104), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(G290), .B1(new_n711), .B2(new_n713), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n933), .A2(new_n599), .A3(new_n712), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(G303), .B(new_n692), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n941), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n943), .A2(new_n938), .A3(new_n937), .A4(new_n939), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT105), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT106), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n932), .B(new_n947), .ZN(new_n948));
  MUX2_X1   g523(.A(new_n853), .B(new_n948), .S(G868), .Z(G295));
  MUX2_X1   g524(.A(new_n853), .B(new_n948), .S(G868), .Z(G331));
  NOR2_X1   g525(.A1(G301), .A2(G286), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n555), .B1(new_n554), .B2(new_n550), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n518), .A2(G64), .ZN(new_n953));
  INV_X1    g528(.A(new_n550), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(KEYINPUT75), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n952), .A2(new_n955), .A3(G651), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n956), .A2(new_n549), .B1(new_n537), .B2(new_n546), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n864), .B1(new_n951), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(G301), .A2(G286), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n956), .A2(new_n537), .A3(new_n546), .A4(new_n549), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n959), .A2(new_n854), .A3(new_n960), .A4(new_n863), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT107), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n961), .A2(KEYINPUT107), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n930), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT108), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n942), .A2(new_n944), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n958), .A2(new_n961), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n967), .A2(new_n920), .A3(new_n921), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n930), .B(new_n970), .C1(new_n962), .C2(new_n963), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n965), .A2(new_n966), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G37), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n923), .A2(new_n963), .A3(new_n962), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n930), .A2(new_n967), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n945), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT110), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n980), .B(new_n945), .C1(new_n976), .C2(new_n977), .ZN(new_n981));
  AND4_X1   g556(.A1(KEYINPUT43), .A2(new_n975), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT41), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n920), .B2(new_n921), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT41), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n951), .A2(new_n864), .A3(new_n957), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n959), .A2(new_n960), .B1(new_n854), .B2(new_n863), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n961), .A2(KEYINPUT107), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n986), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n968), .B1(new_n992), .B2(new_n970), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n966), .B1(new_n993), .B2(new_n965), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT43), .B1(new_n975), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT44), .B1(new_n982), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT43), .B1(new_n974), .B2(new_n994), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT109), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n1000), .B(KEYINPUT43), .C1(new_n974), .C2(new_n994), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT43), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n975), .A2(new_n979), .A3(new_n1002), .A4(new_n981), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n997), .B1(new_n1005), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g581(.A(KEYINPUT123), .ZN(new_n1007));
  INV_X1    g582(.A(G1384), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n888), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g584(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT112), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n883), .A2(new_n886), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n1008), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n888), .A2(new_n1016), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1012), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G2084), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n475), .A2(new_n483), .A3(G40), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1018), .A2(KEYINPUT118), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1012), .A2(new_n1021), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1023), .B1(new_n1024), .B2(G2084), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1020), .B1(new_n1009), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1013), .A2(KEYINPUT45), .A3(new_n1008), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1966), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1022), .A2(G168), .A3(new_n1025), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1031), .A2(new_n1032), .A3(G8), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1034), .A2(new_n1019), .A3(new_n1021), .A4(new_n1012), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1030), .B1(new_n1035), .B2(new_n1023), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1025), .ZN(new_n1037));
  OAI21_X1  g612(.A(G286), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1038), .A2(G8), .A3(new_n1031), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1033), .B1(new_n1039), .B2(KEYINPUT51), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1024), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1034), .A2(KEYINPUT120), .A3(new_n1021), .A4(new_n1012), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1042), .A2(new_n1043), .A3(new_n767), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n888), .A2(KEYINPUT45), .A3(new_n1008), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1026), .B1(G164), .B2(G1384), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1021), .A2(new_n1045), .A3(new_n443), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1047), .A2(KEYINPUT122), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT122), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1027), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1028), .ZN(new_n1052));
  XNOR2_X1  g627(.A(G301), .B(KEYINPUT54), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1044), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1027), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1045), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1044), .A2(new_n1051), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1054), .B1(new_n1056), .B2(new_n1053), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1020), .A2(G2090), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1012), .A2(new_n1015), .A3(new_n1017), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT113), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1034), .A2(new_n1061), .A3(new_n1012), .A4(new_n1058), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1021), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n701), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1060), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G303), .A2(G8), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1068), .B(KEYINPUT55), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1060), .A2(new_n1062), .A3(KEYINPUT114), .A4(new_n1064), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1067), .A2(G8), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  NOR3_X1   g647(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(new_n1020), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G2090), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1076), .A2(new_n1077), .B1(new_n701), .B2(new_n1063), .ZN(new_n1078));
  INV_X1    g653(.A(G8), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1069), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1009), .A2(new_n1020), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT115), .B1(new_n1081), .B2(new_n1079), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1083), .B(G8), .C1(new_n1009), .C2(new_n1020), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n714), .A2(G1976), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT52), .ZN(new_n1088));
  NAND2_X1  g663(.A1(G305), .A2(G1981), .ZN(new_n1089));
  NOR3_X1   g664(.A1(G305), .A2(KEYINPUT117), .A3(G1981), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n1091));
  INV_X1    g666(.A(G1981), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n692), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1089), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT49), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(KEYINPUT49), .B(new_n1089), .C1(new_n1090), .C2(new_n1093), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(new_n1085), .A3(new_n1097), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT116), .B(G1976), .Z(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT52), .B1(G288), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1085), .A2(new_n1086), .A3(new_n1100), .ZN(new_n1101));
  AND4_X1   g676(.A1(new_n1080), .A2(new_n1088), .A3(new_n1098), .A4(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1057), .A2(new_n1072), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1007), .B1(new_n1040), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1031), .A2(G8), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1024), .A2(G2084), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1029), .B1(new_n1106), .B2(KEYINPUT118), .ZN(new_n1107));
  AOI21_X1  g682(.A(G168), .B1(new_n1107), .B2(new_n1025), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT51), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1031), .A2(new_n1032), .A3(G8), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1102), .A2(new_n1072), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1111), .A2(KEYINPUT123), .A3(new_n1112), .A4(new_n1057), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n617), .B(KEYINPUT57), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1021), .A2(new_n1045), .A3(new_n1046), .A4(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1114), .B(new_n1116), .C1(new_n1076), .C2(G1956), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1042), .A2(new_n1043), .A3(new_n827), .ZN(new_n1118));
  INV_X1    g693(.A(G2067), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1081), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n612), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1114), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1116), .ZN(new_n1123));
  AOI21_X1  g698(.A(G1956), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1117), .B1(new_n1121), .B2(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1118), .A2(KEYINPUT60), .A3(new_n1120), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT60), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n612), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1118), .A2(KEYINPUT60), .A3(new_n612), .A4(new_n1120), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT58), .B(G1341), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1063), .A2(G1996), .B1(new_n1081), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n564), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1136), .A3(new_n564), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1125), .A2(new_n1139), .A3(new_n1117), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1125), .B2(new_n1117), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1131), .B(new_n1138), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1127), .B1(new_n1130), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(KEYINPUT121), .B(new_n1127), .C1(new_n1130), .C2(new_n1142), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1104), .A2(new_n1113), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT63), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1102), .A2(new_n1072), .ZN(new_n1149));
  OAI211_X1 g724(.A(G8), .B(G168), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(KEYINPUT119), .B(new_n1148), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1088), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1150), .A2(new_n1155), .A3(new_n1148), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1067), .A2(G8), .A3(new_n1071), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1069), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1156), .A2(new_n1072), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1153), .A2(new_n1154), .A3(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1161));
  OR2_X1    g736(.A1(G288), .A2(G1976), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1161), .B1(new_n1098), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1085), .ZN(new_n1165));
  OAI22_X1  g740(.A1(new_n1072), .A2(new_n1155), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1044), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1102), .A2(new_n1072), .A3(G171), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1168), .B1(new_n1040), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1111), .A2(KEYINPUT62), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1166), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1147), .A2(new_n1160), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1009), .A2(new_n1026), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(new_n1020), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n735), .B(new_n738), .Z(new_n1176));
  XNOR2_X1  g751(.A(new_n818), .B(new_n1119), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n758), .B(new_n762), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n599), .B(new_n728), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1175), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1173), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1175), .A2(new_n762), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT46), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1175), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1177), .A2(new_n759), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  XOR2_X1   g762(.A(new_n1187), .B(KEYINPUT124), .Z(new_n1188));
  INV_X1    g763(.A(KEYINPUT47), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1187), .B(KEYINPUT124), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(KEYINPUT47), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1177), .A2(new_n1178), .A3(new_n738), .A4(new_n735), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n816), .A2(new_n1119), .A3(new_n817), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1185), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1179), .A2(new_n1175), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1175), .A2(new_n728), .A3(new_n599), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT48), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1195), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1190), .A2(new_n1192), .A3(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT125), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1182), .A2(new_n1201), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g777(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1204));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n1205));
  OR2_X1    g779(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1207));
  NAND3_X1  g781(.A1(new_n1206), .A2(new_n687), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g782(.A(new_n1208), .B1(new_n912), .B2(new_n916), .ZN(new_n1209));
  AND3_X1   g783(.A1(new_n1004), .A2(KEYINPUT127), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g784(.A(KEYINPUT127), .B1(new_n1004), .B2(new_n1209), .ZN(new_n1211));
  NOR2_X1   g785(.A1(new_n1210), .A2(new_n1211), .ZN(G308));
  NAND2_X1  g786(.A1(new_n1004), .A2(new_n1209), .ZN(G225));
endmodule


