//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n213, new_n214, new_n215,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1275, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(KEYINPUT65), .ZN(new_n207));
  INV_X1    g0007(.A(G50), .ZN(new_n208));
  NAND3_X1  g0008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n207), .B1(new_n206), .B2(new_n208), .ZN(new_n211));
  NOR3_X1   g0011(.A1(new_n210), .A2(G77), .A3(new_n211), .ZN(G353));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G107), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G87), .ZN(G355));
  NOR2_X1   g0016(.A1(new_n206), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT67), .B(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G238), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G87), .A2(G250), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n231));
  NAND4_X1  g0031(.A1(new_n228), .A2(new_n229), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  AOI22_X1  g0032(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n222), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n221), .B(new_n225), .C1(new_n235), .C2(KEYINPUT1), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n235), .ZN(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G226), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G250), .B(G257), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT69), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n208), .A2(G68), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n202), .A2(G50), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G58), .B(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n250), .B(new_n255), .ZN(G351));
  INV_X1    g0056(.A(KEYINPUT16), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n202), .A2(KEYINPUT67), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G68), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n201), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(G20), .B1(new_n261), .B2(new_n206), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G159), .ZN(new_n265));
  OAI21_X1  g0065(.A(KEYINPUT78), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT78), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n263), .A2(new_n267), .A3(G159), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT7), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n271), .B1(new_n272), .B2(G20), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n226), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n257), .B1(new_n270), .B2(new_n280), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n205), .B(new_n203), .C1(new_n226), .C2(new_n201), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n282), .A2(G20), .B1(new_n266), .B2(new_n268), .ZN(new_n283));
  AOI21_X1  g0083(.A(KEYINPUT7), .B1(new_n278), .B2(new_n219), .ZN(new_n284));
  AOI211_X1 g0084(.A(new_n271), .B(G20), .C1(new_n275), .C2(new_n277), .ZN(new_n285));
  OAI21_X1  g0085(.A(G68), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(new_n286), .A3(KEYINPUT16), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n218), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n281), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n288), .A2(new_n218), .ZN(new_n291));
  INV_X1    g0091(.A(G1), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G13), .A3(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT8), .B(G58), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n292), .B2(G20), .ZN(new_n297));
  INV_X1    g0097(.A(new_n293), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n295), .A2(new_n297), .B1(new_n298), .B2(new_n296), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n290), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n275), .A2(new_n277), .A3(G226), .A4(G1698), .ZN(new_n301));
  INV_X1    g0101(.A(G1698), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n275), .A2(new_n277), .A3(G223), .A4(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G87), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n301), .B(new_n303), .C1(new_n274), .C2(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(G1), .A2(G13), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G41), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n306), .A2(KEYINPUT73), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT73), .B1(new_n306), .B2(new_n307), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G232), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n307), .A2(G1), .A3(G13), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n292), .B1(G41), .B2(G45), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(G274), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n312), .A2(new_n315), .B1(new_n316), .B2(new_n314), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n311), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G169), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n317), .B1(new_n310), .B2(new_n305), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G179), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n300), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT18), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT18), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n300), .A2(new_n326), .A3(new_n323), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n311), .A2(new_n318), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n321), .B2(G200), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n290), .A2(new_n330), .A3(new_n299), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT17), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n290), .A2(new_n330), .A3(KEYINPUT17), .A4(new_n299), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n325), .A2(new_n327), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT79), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n300), .A2(new_n326), .A3(new_n323), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n326), .B1(new_n300), .B2(new_n323), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n333), .A2(new_n334), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT79), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n275), .A2(new_n277), .A3(G232), .A4(G1698), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n275), .A2(new_n277), .A3(G226), .A4(new_n302), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G97), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n310), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n313), .A2(new_n314), .ZN(new_n348));
  INV_X1    g0148(.A(G274), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n306), .B2(new_n307), .ZN(new_n350));
  INV_X1    g0150(.A(new_n314), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n348), .A2(G238), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT13), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n347), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n353), .B1(new_n347), .B2(new_n352), .ZN(new_n355));
  OAI21_X1  g0155(.A(G200), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n347), .A2(new_n352), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT13), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n347), .A2(new_n352), .A3(new_n353), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(G190), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n292), .A2(G20), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n295), .A2(G68), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT11), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n274), .A2(G20), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(G77), .B1(new_n263), .B2(G50), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n258), .A2(new_n260), .A3(G20), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n363), .B1(new_n367), .B2(new_n289), .ZN(new_n368));
  AOI211_X1 g0168(.A(KEYINPUT11), .B(new_n291), .C1(new_n365), .C2(new_n366), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n362), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n293), .A2(KEYINPUT12), .A3(G68), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n226), .A2(new_n298), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT12), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT76), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(KEYINPUT76), .A3(KEYINPUT12), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n371), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n356), .A2(new_n360), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT77), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT77), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n356), .A2(new_n360), .A3(new_n378), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n378), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n354), .A2(new_n355), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G179), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT14), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n387), .B(G169), .C1(new_n354), .C2(new_n355), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G169), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n358), .B2(new_n359), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(new_n387), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n384), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n383), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n296), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n219), .A2(G33), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT15), .B(G87), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n289), .ZN(new_n400));
  INV_X1    g0200(.A(G77), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(new_n292), .B2(G20), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n295), .A2(new_n402), .B1(new_n401), .B2(new_n298), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n275), .A2(new_n277), .A3(G1698), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G238), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n214), .B2(new_n272), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n278), .A2(new_n312), .A3(G1698), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n310), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n316), .A2(new_n314), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(G244), .B2(new_n348), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n404), .B1(new_n413), .B2(G190), .ZN(new_n414));
  INV_X1    g0214(.A(G200), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n413), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n390), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n417), .B(new_n404), .C1(G179), .C2(new_n412), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n336), .A2(new_n342), .A3(new_n394), .A4(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT75), .ZN(new_n422));
  INV_X1    g0222(.A(new_n211), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n219), .B1(new_n423), .B2(new_n209), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n395), .A2(new_n364), .B1(G150), .B2(new_n263), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n289), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n361), .A2(G50), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n294), .A2(new_n428), .B1(G50), .B2(new_n293), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n310), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n275), .A2(new_n277), .A3(G222), .A4(new_n302), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT71), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT71), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n272), .A2(new_n436), .A3(G222), .A4(new_n302), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n401), .B1(new_n275), .B2(new_n277), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(new_n405), .B2(G223), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT72), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT72), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n438), .A2(new_n443), .A3(new_n440), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n433), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  XOR2_X1   g0245(.A(KEYINPUT70), .B(G226), .Z(new_n446));
  AOI21_X1  g0246(.A(new_n410), .B1(new_n348), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT74), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n438), .A2(new_n443), .A3(new_n440), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n443), .B1(new_n438), .B2(new_n440), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n310), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT74), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(new_n447), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G179), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n432), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n449), .A2(new_n390), .A3(new_n454), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n422), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n445), .A2(KEYINPUT74), .A3(new_n448), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n453), .B1(new_n452), .B2(new_n447), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND4_X1   g0262(.A1(new_n422), .A2(new_n462), .A3(new_n431), .A4(new_n458), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n421), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n449), .A2(G200), .A3(new_n454), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n427), .A2(KEYINPUT9), .A3(new_n430), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT9), .B1(new_n427), .B2(new_n430), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n328), .B1(new_n449), .B2(new_n454), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT10), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n455), .A2(G190), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT10), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n473), .A2(new_n474), .A3(new_n466), .A4(new_n469), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n465), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n275), .A2(new_n277), .A3(G250), .A4(G1698), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n275), .A2(new_n277), .A3(G244), .A4(new_n302), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT4), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n478), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n480), .A2(new_n481), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n310), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n292), .A2(G45), .ZN(new_n485));
  OR2_X1    g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  NAND2_X1  g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n350), .ZN(new_n489));
  XNOR2_X1  g0289(.A(KEYINPUT5), .B(G41), .ZN(new_n490));
  INV_X1    g0290(.A(G45), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(G1), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n490), .A2(new_n492), .B1(new_n306), .B2(new_n307), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G257), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n484), .A2(new_n489), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n390), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n484), .A2(new_n456), .A3(new_n494), .A4(new_n489), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n214), .A2(KEYINPUT6), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT80), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n213), .ZN(new_n500));
  NAND2_X1  g0300(.A1(KEYINPUT80), .A2(G97), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G97), .A2(G107), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT6), .B1(new_n215), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(G20), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n263), .A2(G77), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n214), .B1(new_n273), .B2(new_n279), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n289), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n293), .A2(G97), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n291), .B(new_n293), .C1(G1), .C2(new_n274), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n510), .B1(new_n512), .B2(G97), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n496), .A2(new_n497), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT81), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n495), .A2(new_n390), .B1(new_n509), .B2(new_n513), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(KEYINPUT81), .A3(new_n497), .ZN(new_n519));
  INV_X1    g0319(.A(new_n398), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(new_n293), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n511), .A2(new_n304), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n275), .A2(new_n277), .A3(new_n219), .A4(G68), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT19), .ZN(new_n524));
  AND2_X1   g0324(.A1(KEYINPUT80), .A2(G97), .ZN(new_n525));
  NOR2_X1   g0325(.A1(KEYINPUT80), .A2(G97), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n524), .B1(new_n527), .B2(new_n397), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n500), .A2(new_n304), .A3(new_n214), .A4(new_n501), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n219), .B1(new_n345), .B2(new_n524), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n529), .A2(KEYINPUT82), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT82), .B1(new_n529), .B2(new_n530), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n523), .B(new_n528), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  AOI211_X1 g0333(.A(new_n521), .B(new_n522), .C1(new_n533), .C2(new_n289), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n313), .A2(G274), .A3(new_n492), .ZN(new_n535));
  AND2_X1   g0335(.A1(G33), .A2(G41), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n485), .B(G250), .C1(new_n536), .C2(new_n218), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n275), .A2(new_n277), .A3(G244), .A4(G1698), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n275), .A2(new_n277), .A3(G238), .A4(new_n302), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G116), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n538), .B1(new_n542), .B2(new_n310), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n543), .A2(new_n415), .ZN(new_n544));
  AOI211_X1 g0344(.A(new_n328), .B(new_n538), .C1(new_n310), .C2(new_n542), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI211_X1 g0346(.A(G179), .B(new_n538), .C1(new_n310), .C2(new_n542), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n542), .A2(new_n310), .ZN(new_n548));
  INV_X1    g0348(.A(new_n538), .ZN(new_n549));
  AOI21_X1  g0349(.A(G169), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n521), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n511), .A2(new_n398), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n397), .B1(new_n500), .B2(new_n501), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n523), .B1(new_n555), .B2(KEYINPUT19), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n529), .A2(new_n530), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT82), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n529), .A2(KEYINPUT82), .A3(new_n530), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n556), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n552), .B(new_n554), .C1(new_n561), .C2(new_n291), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n534), .A2(new_n546), .B1(new_n551), .B2(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n509), .A2(new_n513), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n495), .A2(G200), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n564), .B(new_n565), .C1(new_n328), .C2(new_n495), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n517), .A2(new_n519), .A3(new_n563), .A4(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n275), .A2(new_n277), .A3(G257), .A4(G1698), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n275), .A2(new_n277), .A3(G250), .A4(new_n302), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G294), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n310), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n493), .A2(G264), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n489), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n415), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n571), .A2(new_n310), .B1(new_n493), .B2(G264), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(new_n328), .A3(new_n489), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(KEYINPUT85), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT85), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n574), .A2(new_n579), .A3(new_n415), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n304), .A2(KEYINPUT84), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n581), .A2(new_n275), .A3(new_n277), .A4(new_n219), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT22), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT22), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n272), .A2(new_n584), .A3(new_n219), .A4(new_n581), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT24), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n541), .A2(G20), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT23), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n219), .B2(G107), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n214), .A2(KEYINPUT23), .A3(G20), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n586), .A2(new_n587), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n587), .B1(new_n586), .B2(new_n592), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n289), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT25), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n293), .B2(G107), .ZN(new_n598));
  NOR3_X1   g0398(.A1(new_n293), .A2(new_n597), .A3(G107), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n512), .A2(G107), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n578), .A2(new_n580), .A3(new_n596), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n574), .A2(new_n390), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n576), .A2(new_n456), .A3(new_n489), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n586), .A2(new_n592), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT24), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n291), .B1(new_n606), .B2(new_n593), .ZN(new_n607));
  INV_X1    g0407(.A(new_n601), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n603), .B(new_n604), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT21), .ZN(new_n611));
  INV_X1    g0411(.A(G116), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n298), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n511), .B2(new_n612), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n219), .B(new_n479), .C1(new_n527), .C2(G33), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT83), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n612), .A2(G20), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n289), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n289), .B2(new_n617), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n615), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT20), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n615), .B(KEYINPUT20), .C1(new_n619), .C2(new_n620), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n614), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n275), .A2(new_n277), .A3(G264), .A4(G1698), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n275), .A2(new_n277), .A3(G257), .A4(new_n302), .ZN(new_n627));
  INV_X1    g0427(.A(G303), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n272), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n310), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n493), .A2(G270), .B1(new_n488), .B2(new_n350), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G169), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n611), .B1(new_n625), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n614), .ZN(new_n635));
  INV_X1    g0435(.A(new_n624), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n289), .A2(new_n617), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT83), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n618), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT20), .B1(new_n639), .B2(new_n615), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n635), .B1(new_n636), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n390), .B1(new_n630), .B2(new_n631), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(KEYINPUT21), .A3(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n630), .A2(new_n631), .A3(G179), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n632), .A2(G200), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n630), .A2(new_n631), .A3(G190), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n625), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n634), .A2(new_n643), .A3(new_n645), .A4(new_n648), .ZN(new_n649));
  NOR4_X1   g0449(.A1(new_n477), .A2(new_n567), .A3(new_n610), .A4(new_n649), .ZN(G372));
  INV_X1    g0450(.A(new_n459), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n457), .A2(new_n422), .A3(new_n458), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT86), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n418), .B1(new_n380), .B2(new_n382), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n391), .A2(new_n387), .B1(new_n385), .B2(G179), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT14), .B1(new_n385), .B2(new_n390), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n378), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n340), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n339), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n472), .A2(new_n475), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n653), .B(new_n654), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n659), .A2(new_n339), .B1(new_n472), .B2(new_n475), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT86), .B1(new_n663), .B2(new_n464), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n562), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n543), .A2(new_n456), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(G169), .B2(new_n543), .ZN(new_n668));
  INV_X1    g0468(.A(new_n522), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n552), .B(new_n669), .C1(new_n561), .C2(new_n291), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n543), .A2(G190), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n415), .B2(new_n543), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n666), .A2(new_n668), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n673), .A2(KEYINPUT26), .A3(new_n515), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n515), .A2(new_n516), .ZN(new_n675));
  AOI21_X1  g0475(.A(KEYINPUT81), .B1(new_n518), .B2(new_n497), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n563), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n674), .B1(new_n677), .B2(KEYINPUT26), .ZN(new_n678));
  INV_X1    g0478(.A(new_n602), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n634), .A2(new_n643), .A3(new_n645), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n609), .ZN(new_n681));
  AND4_X1   g0481(.A1(new_n517), .A2(new_n519), .A3(new_n566), .A4(new_n563), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n551), .A2(new_n562), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n678), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n665), .B1(new_n477), .B2(new_n686), .ZN(G369));
  NAND3_X1  g0487(.A1(new_n292), .A2(new_n219), .A3(G13), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G343), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT87), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n625), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n649), .B2(KEYINPUT88), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(KEYINPUT88), .B2(new_n649), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n680), .A2(new_n696), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(KEYINPUT89), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT89), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n698), .B2(new_n699), .ZN(new_n703));
  OAI21_X1  g0503(.A(G330), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT90), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n606), .A2(new_n593), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n608), .B1(new_n706), .B2(new_n289), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n705), .B1(new_n707), .B2(new_n695), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n693), .B(KEYINPUT87), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n709), .B(KEYINPUT90), .C1(new_n607), .C2(new_n608), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n708), .A2(new_n602), .A3(new_n710), .A4(new_n609), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT91), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n603), .A2(new_n604), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n709), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n711), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n712), .B1(new_n711), .B2(new_n715), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n704), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n680), .A2(new_n709), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n716), .B2(new_n717), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n714), .A2(new_n695), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT92), .ZN(G399));
  INV_X1    g0526(.A(new_n223), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G41), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G1), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n529), .A2(G116), .ZN(new_n731));
  INV_X1    g0531(.A(new_n217), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n730), .A2(new_n731), .B1(new_n732), .B2(new_n729), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  INV_X1    g0534(.A(G330), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n576), .A2(new_n543), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT93), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n484), .A2(new_n494), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT93), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n576), .A2(new_n543), .A3(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n738), .A2(new_n739), .A3(new_n644), .A4(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n543), .A2(G179), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n744), .A2(new_n574), .A3(new_n632), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n742), .A2(new_n743), .B1(new_n745), .B2(new_n495), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n484), .A2(new_n494), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n747), .A2(new_n456), .A3(new_n632), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n748), .A2(KEYINPUT30), .A3(new_n741), .A4(new_n738), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n736), .B(new_n695), .C1(new_n746), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n742), .A2(new_n743), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n745), .A2(new_n495), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n751), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(KEYINPUT31), .B1(new_n753), .B2(new_n709), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n610), .A2(new_n649), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n682), .A2(new_n756), .A3(new_n695), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n735), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n634), .A2(new_n643), .A3(new_n645), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n602), .B1(new_n759), .B2(new_n714), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n684), .B1(new_n760), .B2(new_n567), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT26), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n563), .A2(new_n762), .A3(new_n497), .A4(new_n518), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n673), .B1(new_n517), .B2(new_n519), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(new_n764), .B2(new_n762), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n695), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT29), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(KEYINPUT26), .B1(new_n673), .B2(new_n515), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(new_n677), .B2(KEYINPUT26), .ZN(new_n770));
  OAI211_X1 g0570(.A(KEYINPUT29), .B(new_n695), .C1(new_n770), .C2(new_n761), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n758), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n734), .B1(new_n772), .B2(G1), .ZN(G364));
  OR2_X1    g0573(.A1(new_n701), .A2(new_n703), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(G330), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n219), .A2(G13), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n292), .B1(new_n776), .B2(G45), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n729), .A2(KEYINPUT94), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT94), .ZN(new_n779));
  INV_X1    g0579(.A(new_n777), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n780), .B2(new_n728), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  AND3_X1   g0582(.A1(new_n775), .A2(new_n704), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n727), .A2(new_n278), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT95), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n785), .A2(G355), .B1(new_n612), .B2(new_n727), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n255), .A2(new_n491), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n278), .A2(new_n223), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT96), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(G45), .B2(new_n732), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n786), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G13), .A2(G33), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n218), .B1(G20), .B2(new_n390), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n782), .B1(new_n791), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G179), .A2(G200), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT99), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(G20), .B2(new_n328), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n219), .A2(KEYINPUT99), .A3(G190), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n798), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n265), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT32), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(G20), .A2(G179), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n807), .A2(G190), .A3(G200), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT98), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n805), .B1(new_n812), .B2(new_n208), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n807), .A2(KEYINPUT97), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT97), .ZN(new_n815));
  AOI21_X1  g0615(.A(G200), .B1(new_n806), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n814), .A2(new_n328), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n813), .B1(G77), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n814), .A2(G190), .A3(new_n816), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n803), .A2(new_n804), .B1(new_n201), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n415), .A2(G179), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n800), .B2(new_n801), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n214), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n822), .A2(G20), .A3(G190), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n806), .A2(new_n415), .A3(G190), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n272), .B1(new_n825), .B2(new_n304), .C1(new_n827), .C2(new_n202), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n798), .A2(G190), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G20), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(new_n213), .ZN(new_n832));
  NOR4_X1   g0632(.A1(new_n821), .A2(new_n824), .A3(new_n828), .A4(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G283), .ZN(new_n834));
  INV_X1    g0634(.A(G329), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n834), .A2(new_n823), .B1(new_n802), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(G294), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n278), .B1(new_n825), .B2(new_n628), .C1(new_n831), .C2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(KEYINPUT33), .B(G317), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n836), .B(new_n838), .C1(new_n826), .C2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n812), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(G326), .ZN(new_n842));
  INV_X1    g0642(.A(new_n820), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G311), .A2(new_n818), .B1(new_n843), .B2(G322), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n819), .A2(new_n833), .B1(new_n840), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n795), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n797), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(new_n700), .B2(new_n794), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n783), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G396));
  NOR2_X1   g0651(.A1(new_n418), .A2(new_n709), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n709), .A2(new_n404), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n416), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n852), .B1(new_n854), .B2(new_n418), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n766), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n419), .A2(new_n709), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n685), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n753), .A2(new_n709), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n736), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n709), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n757), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(G330), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n782), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n860), .A2(new_n865), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n866), .B1(KEYINPUT100), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(KEYINPUT100), .B2(new_n867), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n278), .B1(new_n825), .B2(new_n214), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n870), .B(new_n832), .C1(G283), .C2(new_n826), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n841), .A2(G303), .B1(G294), .B2(new_n843), .ZN(new_n872));
  INV_X1    g0672(.A(new_n823), .ZN(new_n873));
  INV_X1    g0673(.A(new_n802), .ZN(new_n874));
  AOI22_X1  g0674(.A1(G87), .A2(new_n873), .B1(new_n874), .B2(G311), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n818), .A2(G116), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n871), .A2(new_n872), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n843), .A2(G143), .B1(G150), .B2(new_n826), .ZN(new_n878));
  INV_X1    g0678(.A(G137), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n878), .B1(new_n265), .B2(new_n817), .C1(new_n812), .C2(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT34), .Z(new_n881));
  OAI21_X1  g0681(.A(new_n272), .B1(new_n825), .B2(new_n208), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(G58), .B2(new_n830), .ZN(new_n883));
  INV_X1    g0683(.A(G132), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n883), .B1(new_n202), .B2(new_n823), .C1(new_n884), .C2(new_n802), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n877), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n795), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n795), .A2(new_n792), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n782), .B1(new_n401), .B2(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n887), .B(new_n889), .C1(new_n855), .C2(new_n793), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n869), .A2(new_n890), .ZN(G384));
  OR2_X1    g0691(.A1(new_n502), .A2(new_n504), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n892), .A2(KEYINPUT35), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(KEYINPUT35), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n893), .A2(G116), .A3(new_n220), .A4(new_n894), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n895), .B(KEYINPUT36), .Z(new_n896));
  OAI211_X1 g0696(.A(new_n217), .B(G77), .C1(new_n201), .C2(new_n226), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n292), .B(G13), .C1(new_n897), .C2(new_n251), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n776), .A2(new_n292), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n852), .B(KEYINPUT101), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n685), .B2(new_n858), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n383), .A2(new_n393), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n384), .A2(new_n709), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n383), .A2(new_n393), .A3(new_n905), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n903), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n300), .A2(new_n692), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT37), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n324), .A2(new_n911), .A3(new_n912), .A4(new_n331), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n290), .A2(new_n330), .A3(new_n299), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n202), .B1(new_n273), .B2(new_n279), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n257), .B1(new_n270), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(new_n287), .A3(new_n289), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n917), .A2(new_n299), .B1(new_n320), .B2(new_n322), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n691), .B1(new_n917), .B2(new_n299), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n914), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n913), .B1(new_n920), .B2(new_n912), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT102), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT102), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n923), .B(new_n913), .C1(new_n920), .C2(new_n912), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n335), .A2(new_n919), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n922), .A2(KEYINPUT38), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n921), .A2(KEYINPUT102), .B1(new_n335), .B2(new_n919), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n928), .B2(new_n924), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n910), .A2(new_n930), .B1(new_n339), .B2(new_n692), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n658), .A2(new_n695), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT39), .B1(new_n927), .B2(new_n929), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n926), .A2(KEYINPUT103), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT103), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n928), .A2(new_n935), .A3(KEYINPUT38), .A4(new_n924), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n335), .A2(new_n300), .A3(new_n692), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n324), .A2(new_n911), .A3(new_n331), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT37), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n913), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT38), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT39), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n934), .A2(new_n936), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n932), .B1(new_n933), .B2(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n931), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n465), .A2(new_n768), .A3(new_n476), .A4(new_n771), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n665), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n946), .B(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n465), .A2(new_n476), .A3(new_n864), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT104), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n864), .A2(new_n855), .A3(new_n909), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n927), .B2(new_n929), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT40), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n941), .A2(new_n942), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n934), .A2(new_n936), .A3(new_n956), .ZN(new_n957));
  AND4_X1   g0757(.A1(KEYINPUT40), .A2(new_n864), .A3(new_n855), .A4(new_n909), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(G330), .B1(new_n951), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n960), .B2(new_n951), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n900), .B1(new_n949), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT105), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n963), .A2(new_n964), .B1(new_n949), .B2(new_n962), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n899), .B1(new_n965), .B2(new_n966), .ZN(G367));
  NOR2_X1   g0767(.A1(new_n675), .A2(new_n676), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n968), .B(new_n566), .C1(new_n564), .C2(new_n695), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n518), .A2(new_n709), .A3(new_n497), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n722), .A2(new_n723), .A3(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT45), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n722), .A2(new_n723), .ZN(new_n976));
  INV_X1    g0776(.A(new_n971), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT44), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n979), .B(new_n971), .C1(new_n722), .C2(new_n723), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n974), .A2(new_n975), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n719), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n718), .B1(new_n680), .B2(new_n709), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n774), .A2(G330), .A3(new_n722), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n722), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n704), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n984), .A2(new_n772), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n979), .B1(new_n724), .B2(new_n971), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n976), .A2(KEYINPUT44), .A3(new_n977), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n972), .B(new_n973), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n990), .A2(new_n720), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n982), .A2(new_n987), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n772), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n728), .B(KEYINPUT41), .Z(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT108), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT108), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n998), .B(new_n995), .C1(new_n993), .C2(new_n772), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n777), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n723), .A2(KEYINPUT42), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n976), .A2(new_n971), .A3(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n716), .A2(new_n717), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1003), .A2(new_n721), .A3(new_n971), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(KEYINPUT42), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1002), .B(new_n1005), .C1(new_n968), .C2(new_n709), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n695), .A2(new_n534), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n563), .B(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT43), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1008), .B(KEYINPUT43), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT106), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n719), .A2(new_n971), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n1016), .A2(KEYINPUT106), .B1(new_n1017), .B2(KEYINPUT107), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1017), .A2(KEYINPUT107), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1000), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n825), .ZN(new_n1023));
  AOI21_X1  g0823(.A(KEYINPUT46), .B1(new_n1023), .B2(G116), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n831), .A2(new_n214), .B1(new_n827), .B2(new_n837), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(G283), .C2(new_n818), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n874), .A2(G317), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n841), .A2(G311), .B1(G303), .B2(new_n843), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT46), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n825), .A2(new_n1029), .A3(new_n612), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n527), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n272), .B(new_n1030), .C1(new_n1031), .C2(new_n873), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n830), .A2(G68), .ZN(new_n1034));
  INV_X1    g0834(.A(G150), .ZN(new_n1035));
  INV_X1    g0835(.A(G143), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1034), .B1(new_n1035), .B2(new_n820), .C1(new_n812), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT109), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n823), .A2(new_n401), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n272), .B1(new_n825), .B2(new_n201), .C1(new_n827), .C2(new_n265), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(G137), .C2(new_n874), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1039), .B(new_n1042), .C1(new_n208), .C2(new_n817), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1033), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT47), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n795), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1008), .A2(new_n794), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n246), .A2(new_n789), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n795), .B(new_n794), .C1(new_n727), .C2(new_n520), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n782), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1047), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1022), .A2(new_n1052), .ZN(G387));
  AOI21_X1  g0853(.A(new_n278), .B1(new_n1023), .B2(G77), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n520), .A2(new_n830), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n213), .C2(new_n823), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G150), .B2(new_n874), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n817), .A2(new_n202), .B1(new_n296), .B2(new_n827), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT110), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n841), .A2(G159), .B1(G50), .B2(new_n843), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G303), .A2(new_n818), .B1(new_n843), .B2(G317), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1062), .A2(KEYINPUT111), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(KEYINPUT111), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n841), .A2(G322), .B1(G311), .B2(new_n826), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT48), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n831), .A2(new_n834), .B1(new_n825), .B2(new_n837), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(KEYINPUT49), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n272), .B1(new_n874), .B2(G326), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n612), .C2(new_n823), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT49), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1061), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT112), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n847), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n1076), .B2(new_n1075), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n718), .A2(new_n794), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n789), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n242), .B2(G45), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n731), .B2(new_n785), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n395), .A2(new_n208), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT50), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n491), .B1(new_n202), .B2(new_n401), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n1084), .A2(new_n731), .A3(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1082), .A2(new_n1086), .B1(G107), .B2(new_n223), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n782), .B1(new_n1087), .B2(new_n796), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1078), .A2(new_n1079), .A3(new_n1088), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT113), .Z(new_n1090));
  NAND3_X1  g0890(.A1(new_n984), .A2(new_n780), .A3(new_n986), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n987), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n728), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n772), .B1(new_n984), .B2(new_n986), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1090), .B(new_n1091), .C1(new_n1093), .C2(new_n1094), .ZN(G393));
  NAND3_X1  g0895(.A1(new_n982), .A2(new_n992), .A3(new_n780), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n841), .A2(G317), .B1(G311), .B2(new_n843), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT114), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1098), .A2(KEYINPUT52), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n278), .B1(new_n825), .B2(new_n834), .C1(new_n831), .C2(new_n612), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G303), .B2(new_n826), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n824), .B1(G322), .B2(new_n874), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(new_n837), .C2(new_n817), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1098), .A2(KEYINPUT52), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n812), .A2(new_n1035), .B1(new_n265), .B2(new_n820), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT51), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n304), .A2(new_n823), .B1(new_n802), .B2(new_n1036), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n831), .A2(new_n401), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n278), .B(new_n1109), .C1(new_n227), .C2(new_n1023), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n208), .B2(new_n827), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1108), .B(new_n1111), .C1(new_n395), .C2(new_n818), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1104), .A2(new_n1105), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT115), .Z(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n795), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n782), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n977), .A2(new_n794), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n796), .B1(new_n223), .B2(new_n527), .C1(new_n1080), .C2(new_n250), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1096), .A2(new_n1119), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n993), .A2(new_n728), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n982), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n992), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1092), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1120), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(G390));
  AOI21_X1  g0926(.A(new_n909), .B1(new_n758), .B2(new_n855), .ZN(new_n1127));
  AND4_X1   g0927(.A1(G330), .A2(new_n864), .A3(new_n855), .A4(new_n909), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n903), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n909), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n865), .B2(new_n856), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n854), .A2(new_n418), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n695), .B(new_n1132), .C1(new_n770), .C2(new_n761), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n852), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n758), .A2(new_n855), .A3(new_n909), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1131), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1129), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n465), .A2(new_n476), .A3(new_n758), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n665), .A2(new_n947), .A3(new_n1140), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1139), .A2(new_n1141), .A3(KEYINPUT117), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT117), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n932), .B1(new_n902), .B2(new_n1130), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n933), .A2(new_n1145), .A3(new_n944), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1135), .A2(new_n909), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n957), .A2(new_n932), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1128), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT116), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1146), .A2(new_n1148), .A3(new_n1137), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1146), .A2(new_n1148), .A3(new_n1137), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1137), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT116), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1144), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1141), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1129), .A2(new_n1138), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n729), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1158), .A2(new_n780), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n933), .A2(new_n944), .A3(new_n792), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n888), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1116), .B1(new_n395), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n278), .B1(new_n825), .B2(new_n304), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1168), .B(new_n1109), .C1(G107), .C2(new_n826), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n841), .A2(G283), .B1(G116), .B2(new_n843), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G68), .A2(new_n873), .B1(new_n874), .B2(G294), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n818), .A2(new_n1031), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n272), .B1(new_n823), .B2(new_n208), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G125), .B2(new_n874), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT119), .Z(new_n1176));
  XOR2_X1   g0976(.A(KEYINPUT54), .B(G143), .Z(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT118), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n841), .A2(G128), .B1(new_n818), .B2(new_n1178), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n831), .A2(new_n265), .B1(new_n827), .B2(new_n879), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT53), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n825), .B2(new_n1035), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1023), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1180), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1179), .B(new_n1184), .C1(new_n884), .C2(new_n820), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1173), .B1(new_n1176), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1167), .B1(new_n1186), .B2(new_n795), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1165), .A2(new_n1187), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1164), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1163), .A2(new_n1189), .ZN(G378));
  AOI22_X1  g0990(.A1(new_n841), .A2(G116), .B1(new_n520), .B2(new_n818), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n214), .B2(new_n820), .ZN(new_n1192));
  AOI211_X1 g0992(.A(G41), .B(new_n272), .C1(new_n1023), .C2(G77), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1193), .B(new_n1034), .C1(new_n213), .C2(new_n827), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n873), .A2(G58), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n834), .B2(new_n802), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1192), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1197), .A2(KEYINPUT58), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(G33), .A2(G41), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1199), .A2(G50), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n272), .B2(G41), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n1197), .B2(KEYINPUT58), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT120), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n841), .A2(G125), .B1(G137), .B2(new_n818), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n843), .A2(G128), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1178), .A2(new_n1023), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n830), .A2(G150), .B1(G132), .B2(new_n826), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  INV_X1    g1009(.A(G124), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1199), .B1(new_n802), .B2(new_n1210), .C1(new_n265), .C2(new_n823), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1208), .B2(KEYINPUT59), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1198), .B(new_n1203), .C1(new_n1209), .C2(new_n1212), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1116), .B1(G50), .B2(new_n1166), .C1(new_n1213), .C2(new_n847), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n457), .A2(new_n458), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n476), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1216), .A2(new_n431), .A3(new_n692), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n476), .B(new_n1215), .C1(new_n432), .C2(new_n691), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  XOR2_X1   g1019(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1217), .A2(new_n1220), .A3(new_n1218), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1214), .B1(new_n792), .B2(new_n1224), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT121), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n955), .A2(new_n959), .A3(G330), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n931), .A2(new_n945), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n735), .B1(new_n953), .B2(new_n954), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(new_n1224), .A3(new_n959), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1229), .A2(new_n1230), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1230), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1226), .B1(new_n1236), .B2(new_n780), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1141), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT57), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1224), .B1(new_n1231), .B2(new_n959), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n946), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(KEYINPUT57), .A3(new_n1233), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1159), .B1(new_n1158), .B2(new_n1139), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n728), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1237), .B1(new_n1240), .B2(new_n1246), .ZN(G375));
  NAND2_X1  g1047(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1144), .A2(new_n996), .A3(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n782), .B1(new_n202), .B2(new_n888), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n272), .B1(new_n1023), .B2(G97), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1251), .B(new_n1055), .C1(new_n612), .C2(new_n827), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1040), .B(new_n1252), .C1(G303), .C2(new_n874), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n812), .A2(new_n837), .B1(new_n834), .B2(new_n820), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(G107), .B2(new_n818), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n812), .A2(new_n884), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT122), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1178), .A2(new_n826), .B1(G128), .B2(new_n874), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n272), .B1(new_n825), .B2(new_n265), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G50), .B2(new_n830), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(G150), .A2(new_n818), .B1(new_n843), .B2(G137), .ZN(new_n1261));
  AND4_X1   g1061(.A1(new_n1195), .A2(new_n1258), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1253), .A2(new_n1255), .B1(new_n1257), .B2(new_n1262), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1250), .B1(new_n847), .B2(new_n1263), .C1(new_n909), .C2(new_n793), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1139), .B2(new_n780), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1249), .A2(new_n1266), .ZN(new_n1267));
  XOR2_X1   g1067(.A(new_n1267), .B(KEYINPUT123), .Z(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(G381));
  NOR2_X1   g1069(.A1(G387), .A2(G375), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1164), .A2(new_n1188), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(new_n1157), .B2(new_n1162), .ZN(new_n1272));
  NOR4_X1   g1072(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1270), .A2(new_n1272), .A3(new_n1268), .A4(new_n1273), .ZN(G407));
  OR2_X1    g1074(.A1(G378), .A2(G343), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G407), .B(G213), .C1(G375), .C2(new_n1275), .ZN(G409));
  INV_X1    g1076(.A(G213), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1277), .A2(G343), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G378), .B(new_n1237), .C1(new_n1240), .C2(new_n1246), .ZN(new_n1279));
  NOR4_X1   g1079(.A1(new_n1245), .A2(new_n1234), .A3(new_n995), .A4(new_n1235), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1226), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1243), .A2(new_n780), .A3(new_n1233), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1272), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1278), .B1(new_n1279), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT60), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1248), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1159), .A2(new_n1160), .A3(KEYINPUT60), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n728), .A3(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(G384), .A3(new_n1266), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G384), .B1(new_n1289), .B2(new_n1266), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1285), .A2(new_n1293), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1294), .A2(KEYINPUT62), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G2897), .B(new_n1278), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1292), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1278), .A2(G2897), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1290), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1296), .B1(new_n1285), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT127), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1304), .B(new_n1296), .C1(new_n1285), .C2(new_n1301), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1294), .A2(KEYINPUT62), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1295), .A2(new_n1303), .A3(new_n1305), .A4(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT124), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(G393), .B(new_n850), .ZN(new_n1309));
  AOI21_X1  g1109(.A(G390), .B1(new_n1022), .B2(new_n1052), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1052), .ZN(new_n1311));
  AOI211_X1 g1111(.A(new_n1311), .B(new_n1125), .C1(new_n1000), .C2(new_n1021), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1308), .B(new_n1309), .C1(new_n1310), .C2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1309), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(KEYINPUT124), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1310), .A2(new_n1309), .ZN(new_n1316));
  OAI21_X1  g1116(.A(KEYINPUT125), .B1(G387), .B2(new_n1125), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT125), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1312), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1316), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1315), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1307), .A2(new_n1313), .A3(new_n1321), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1285), .A2(KEYINPUT63), .A3(new_n1293), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT63), .B1(new_n1285), .B2(new_n1293), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1323), .A2(new_n1302), .A3(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT126), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1315), .A2(new_n1320), .A3(new_n1313), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1325), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1326), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1322), .B1(new_n1328), .B2(new_n1329), .ZN(G405));
  NAND2_X1  g1130(.A1(G375), .A2(new_n1272), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1279), .ZN(new_n1332));
  XOR2_X1   g1132(.A(new_n1332), .B(new_n1293), .Z(new_n1333));
  XNOR2_X1  g1133(.A(new_n1327), .B(new_n1333), .ZN(G402));
endmodule


