//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1274, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n203), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  INV_X1    g0024(.A(G97), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n201), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n246), .A2(G1), .A3(G13), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G223), .A2(G1698), .ZN(new_n249));
  INV_X1    g0049(.A(G222), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n249), .B1(new_n250), .B2(G1698), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n252), .B1(new_n253), .B2(new_n248), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT64), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n247), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(new_n255), .B2(new_n254), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n247), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  AND2_X1   g0060(.A1(G1), .A2(G13), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(new_n246), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n259), .A2(G226), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n257), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G169), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n215), .ZN(new_n271));
  OAI21_X1  g0071(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n272));
  INV_X1    g0072(.A(G150), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n272), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT65), .B1(new_n278), .B2(G20), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT65), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(new_n207), .A3(G33), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n277), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n271), .B1(new_n276), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(G50), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n271), .B1(new_n206), .B2(G20), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(G50), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n269), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT66), .B(G179), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n267), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n284), .A2(G77), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n286), .B2(G77), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT15), .B(G87), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n279), .B2(new_n281), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n277), .A2(new_n275), .B1(new_n207), .B2(new_n253), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n271), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT67), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n207), .A2(new_n253), .ZN(new_n303));
  XOR2_X1   g0103(.A(KEYINPUT8), .B(G58), .Z(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n274), .ZN(new_n305));
  INV_X1    g0105(.A(new_n297), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n279), .A2(new_n281), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(KEYINPUT67), .A3(new_n271), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n296), .B1(new_n302), .B2(new_n310), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n259), .A2(G244), .B1(new_n262), .B2(new_n265), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT3), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G107), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n247), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(G232), .A2(G1698), .ZN(new_n319));
  INV_X1    g0119(.A(G1698), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(G238), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n248), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n312), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n268), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n312), .A2(new_n323), .A3(new_n290), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n311), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n324), .A2(G200), .ZN(new_n329));
  INV_X1    g0129(.A(G190), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n324), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT67), .B1(new_n309), .B2(new_n271), .ZN(new_n332));
  INV_X1    g0132(.A(new_n271), .ZN(new_n333));
  AOI211_X1 g0133(.A(new_n301), .B(new_n333), .C1(new_n305), .C2(new_n308), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n295), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n293), .A2(new_n328), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT68), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n267), .A2(G200), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT9), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n288), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n283), .A2(KEYINPUT9), .A3(new_n287), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n267), .A2(new_n330), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT10), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n345), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT10), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n347), .A2(new_n348), .A3(new_n339), .A4(new_n343), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n337), .A2(new_n338), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G226), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n320), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n224), .A2(G1698), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n313), .A2(new_n353), .A3(new_n315), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G33), .A2(G97), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n247), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT13), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n265), .A2(new_n247), .A3(G274), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n247), .A2(G238), .A3(new_n258), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n358), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT69), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n357), .A2(new_n362), .A3(KEYINPUT13), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT69), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT13), .B1(new_n357), .B2(new_n362), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n365), .A2(new_n368), .A3(G190), .A4(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n369), .ZN(new_n371));
  OAI21_X1  g0171(.A(G200), .B1(new_n371), .B2(new_n366), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n253), .B1(new_n279), .B2(new_n281), .ZN(new_n374));
  INV_X1    g0174(.A(G50), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n275), .A2(new_n375), .B1(new_n207), .B2(G68), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n271), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT70), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI211_X1 g0179(.A(KEYINPUT70), .B(new_n271), .C1(new_n374), .C2(new_n376), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT11), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT11), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n379), .A2(new_n383), .A3(new_n380), .ZN(new_n384));
  INV_X1    g0184(.A(new_n284), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n202), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT12), .B1(new_n386), .B2(KEYINPUT71), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(KEYINPUT71), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(KEYINPUT71), .A3(KEYINPUT12), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n389), .A2(new_n390), .B1(G68), .B2(new_n286), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n382), .A2(new_n384), .A3(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n373), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(G169), .B1(new_n371), .B2(new_n366), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT14), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n365), .A2(new_n368), .A3(G179), .A4(new_n369), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT14), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n397), .B(G169), .C1(new_n371), .C2(new_n366), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n393), .B1(new_n392), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n351), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT73), .ZN(new_n402));
  OR2_X1    g0202(.A1(G223), .A2(G1698), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n352), .A2(G1698), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n313), .A2(new_n403), .A3(new_n315), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n247), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n259), .A2(G232), .B1(new_n262), .B2(new_n265), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(new_n330), .ZN(new_n410));
  INV_X1    g0210(.A(G200), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n247), .A2(new_n258), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n360), .B1(new_n224), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n411), .B1(new_n413), .B2(new_n407), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n304), .A2(new_n284), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n304), .B2(new_n286), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT7), .B1(new_n316), .B2(new_n207), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n207), .A2(KEYINPUT7), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n248), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(G68), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n201), .A2(new_n202), .ZN(new_n422));
  NOR2_X1   g0222(.A1(G58), .A2(G68), .ZN(new_n423));
  OAI21_X1  g0223(.A(G20), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n274), .A2(G159), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n421), .A2(KEYINPUT16), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n271), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT72), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n313), .A2(new_n315), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n278), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT7), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(G20), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(G20), .B1(new_n313), .B2(new_n315), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n431), .A2(new_n435), .B1(new_n436), .B2(KEYINPUT7), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G68), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT16), .B1(new_n438), .B2(new_n427), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n415), .B(new_n417), .C1(new_n429), .C2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT17), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n417), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n436), .A2(KEYINPUT7), .B1(new_n248), .B2(new_n419), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n426), .B1(new_n444), .B2(G68), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n333), .B1(new_n445), .B2(KEYINPUT16), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT16), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n434), .B(new_n432), .C1(new_n316), .C2(KEYINPUT72), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n433), .B1(new_n248), .B2(G20), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n202), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n447), .B1(new_n450), .B2(new_n426), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n443), .B1(new_n446), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT17), .B1(new_n452), .B2(new_n415), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n402), .B1(new_n442), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n268), .B1(new_n408), .B2(new_n409), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n413), .A2(new_n407), .A3(new_n290), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT18), .B1(new_n452), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n417), .B1(new_n429), .B2(new_n439), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT18), .ZN(new_n460));
  INV_X1    g0260(.A(new_n457), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n440), .A2(new_n441), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n452), .A2(KEYINPUT17), .A3(new_n415), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT73), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n454), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n338), .B1(new_n337), .B2(new_n350), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n401), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(new_n207), .C1(G33), .C2(new_n225), .ZN(new_n472));
  INV_X1    g0272(.A(G116), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G20), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n271), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT20), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n472), .A2(KEYINPUT20), .A3(new_n271), .A4(new_n474), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(KEYINPUT77), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n284), .A2(new_n473), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n206), .A2(G33), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n284), .A2(new_n481), .A3(new_n215), .A4(new_n270), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n480), .B1(new_n483), .B2(new_n473), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT77), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n475), .A2(new_n485), .A3(new_n476), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n479), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G303), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n247), .B1(new_n316), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(G257), .A2(G1698), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n320), .A2(G264), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n248), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n206), .B(G45), .C1(new_n263), .C2(KEYINPUT5), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT75), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n264), .A2(G1), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT75), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT5), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G41), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n263), .A2(KEYINPUT5), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n495), .A2(new_n500), .A3(new_n501), .A4(new_n262), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n496), .A2(new_n501), .A3(new_n499), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(G270), .A3(new_n247), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n493), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n487), .A2(KEYINPUT21), .A3(G169), .A4(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G179), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n487), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT21), .ZN(new_n511));
  INV_X1    g0311(.A(new_n487), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n505), .A2(G169), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n505), .A2(G200), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n512), .B(new_n515), .C1(new_n330), .C2(new_n505), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n510), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n503), .A2(G257), .A3(new_n247), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n502), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(G244), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(G1698), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n521), .A2(new_n313), .A3(new_n315), .A4(KEYINPUT4), .ZN(new_n522));
  AND2_X1   g0322(.A1(G250), .A2(G1698), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n313), .A2(new_n315), .A3(new_n523), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n522), .A2(new_n471), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n521), .A2(new_n313), .A3(new_n315), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT74), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT74), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n530), .A3(new_n527), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n525), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n247), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n519), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G190), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n248), .A2(new_n523), .B1(G33), .B2(G283), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT4), .B1(new_n248), .B2(new_n521), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n536), .B(new_n522), .C1(new_n537), .C2(new_n530), .ZN(new_n538));
  INV_X1    g0338(.A(new_n531), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n533), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n519), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n411), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n535), .B1(new_n542), .B2(KEYINPUT76), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n317), .B1(new_n448), .B2(new_n449), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n317), .A2(KEYINPUT6), .A3(G97), .ZN(new_n545));
  XNOR2_X1  g0345(.A(G97), .B(G107), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT6), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n548), .A2(new_n207), .B1(new_n253), .B2(new_n275), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n271), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n284), .A2(G97), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n483), .B2(G97), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  AOI211_X1 g0353(.A(new_n330), .B(new_n519), .C1(new_n532), .C2(new_n533), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT76), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n543), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n522), .A2(new_n471), .A3(new_n524), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n530), .B1(new_n526), .B2(new_n527), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n539), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n541), .B1(new_n560), .B2(new_n247), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n268), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n534), .A2(new_n290), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n563), .A3(new_n553), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n313), .A2(new_n315), .A3(new_n207), .A4(G68), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n207), .B1(new_n356), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n220), .A2(new_n225), .A3(new_n317), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n225), .B1(new_n279), .B2(new_n281), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n566), .B(new_n570), .C1(new_n571), .C2(KEYINPUT19), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n271), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n297), .A2(new_n385), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n483), .A2(new_n306), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n219), .A2(new_n320), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n520), .A2(G1698), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n313), .A2(new_n577), .A3(new_n315), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G116), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n247), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n496), .A2(new_n260), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n221), .B1(new_n264), .B2(G1), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n247), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n268), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n581), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n290), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n576), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n572), .A2(new_n271), .B1(new_n385), .B2(new_n297), .ZN(new_n590));
  OAI21_X1  g0390(.A(G200), .B1(new_n581), .B2(new_n585), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n579), .A2(new_n580), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n533), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(G190), .A3(new_n584), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n483), .A2(G87), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n590), .A2(new_n591), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n589), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n498), .A2(G41), .ZN(new_n598));
  OAI211_X1 g0398(.A(G264), .B(new_n247), .C1(new_n494), .C2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT78), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n503), .A2(KEYINPUT78), .A3(G264), .A4(new_n247), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n226), .A2(G1698), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(G250), .B2(G1698), .ZN(new_n604));
  INV_X1    g0404(.A(G294), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n604), .A2(new_n316), .B1(new_n278), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n601), .A2(new_n602), .B1(new_n606), .B2(new_n533), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(new_n507), .A3(new_n502), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n601), .A2(new_n602), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n533), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n502), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n268), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n313), .A2(new_n315), .A3(new_n207), .A4(G87), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT22), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT22), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n248), .A2(new_n615), .A3(new_n207), .A4(G87), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n580), .A2(G20), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT23), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n207), .B2(G107), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n317), .A2(KEYINPUT23), .A3(G20), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT24), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT24), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n617), .A2(new_n625), .A3(new_n622), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n333), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n385), .A2(KEYINPUT25), .A3(new_n317), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT25), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n284), .B2(G107), .ZN(new_n630));
  AOI22_X1  g0430(.A1(G107), .A2(new_n483), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n608), .B(new_n612), .C1(new_n627), .C2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n617), .A2(new_n625), .A3(new_n622), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n625), .B1(new_n617), .B2(new_n622), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n271), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n611), .A2(G200), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n607), .A2(G190), .A3(new_n502), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n636), .A2(new_n637), .A3(new_n631), .A4(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n597), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  NOR4_X1   g0440(.A1(new_n470), .A2(new_n517), .A3(new_n565), .A4(new_n640), .ZN(G372));
  INV_X1    g0441(.A(KEYINPUT81), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n350), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n346), .A2(new_n349), .A3(KEYINPUT81), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n399), .A2(new_n392), .ZN(new_n646));
  INV_X1    g0446(.A(new_n328), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n393), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n454), .A3(new_n466), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n463), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n293), .B1(new_n645), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n590), .A2(new_n595), .A3(new_n594), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT79), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n584), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n582), .A2(KEYINPUT79), .A3(new_n247), .A4(new_n583), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n411), .B1(new_n657), .B2(new_n593), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n590), .A2(new_n575), .B1(new_n290), .B2(new_n587), .ZN(new_n660));
  AOI21_X1  g0460(.A(G169), .B1(new_n657), .B2(new_n593), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n653), .A2(new_n659), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n557), .A2(new_n564), .A3(new_n639), .A4(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n514), .A2(new_n509), .A3(new_n506), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n624), .A2(new_n626), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n632), .B1(new_n666), .B2(new_n271), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n612), .A2(new_n608), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT80), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n636), .A2(new_n631), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT80), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n670), .A2(new_n671), .A3(new_n608), .A4(new_n612), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n665), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n664), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n660), .A2(new_n662), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n589), .A2(new_n596), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT26), .B1(new_n564), .B2(new_n676), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n562), .A2(new_n563), .A3(new_n553), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n663), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n675), .B(new_n677), .C1(new_n679), .C2(KEYINPUT26), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n651), .B1(new_n470), .B2(new_n681), .ZN(G369));
  AND2_X1   g0482(.A1(new_n633), .A2(new_n639), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT27), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(new_n206), .A3(new_n207), .A4(G13), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT82), .ZN(new_n686));
  INV_X1    g0486(.A(G213), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n687), .B1(new_n688), .B2(KEYINPUT27), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n686), .A2(KEYINPUT83), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT83), .B1(new_n686), .B2(new_n689), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  OR3_X1    g0494(.A1(new_n667), .A2(KEYINPUT85), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT85), .B1(new_n667), .B2(new_n694), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n683), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n633), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n693), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n694), .A2(new_n512), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n665), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n517), .B2(new_n701), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n703), .A2(KEYINPUT84), .A3(G330), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT84), .B1(new_n703), .B2(G330), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n700), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n669), .A2(new_n672), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n693), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n683), .A2(new_n695), .A3(new_n696), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n665), .A2(new_n694), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n708), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n706), .A2(new_n712), .ZN(G399));
  INV_X1    g0513(.A(new_n210), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n569), .A2(G116), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G1), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n213), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  NOR4_X1   g0520(.A1(new_n565), .A2(new_n640), .A3(new_n517), .A4(new_n693), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  INV_X1    g0522(.A(new_n505), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n607), .A3(G179), .A4(new_n587), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n724), .B2(new_n561), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n723), .A2(new_n291), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n657), .A2(new_n593), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n726), .A2(new_n561), .A3(new_n611), .A4(new_n727), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n607), .A2(new_n587), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(KEYINPUT30), .A3(new_n534), .A4(new_n508), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n725), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n693), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(G330), .B1(new_n721), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n681), .A2(new_n693), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n739), .A2(KEYINPUT29), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n576), .A2(new_n588), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n741), .A2(new_n661), .B1(new_n652), .B2(new_n658), .ZN(new_n742));
  OAI21_X1  g0542(.A(KEYINPUT26), .B1(new_n564), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT26), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n561), .A2(new_n268), .B1(new_n550), .B2(new_n552), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n597), .A2(new_n744), .A3(new_n563), .A4(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n743), .A2(new_n746), .A3(new_n675), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n663), .A2(new_n639), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n543), .A2(new_n556), .B1(new_n745), .B2(new_n563), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n633), .A2(new_n510), .A3(new_n514), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT86), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n747), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n748), .A2(new_n749), .A3(KEYINPUT86), .A4(new_n750), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n693), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT29), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n738), .B1(new_n740), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n720), .B1(new_n757), .B2(G1), .ZN(G364));
  NOR2_X1   g0558(.A1(new_n704), .A2(new_n705), .ZN(new_n759));
  INV_X1    g0559(.A(G13), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n206), .B1(new_n761), .B2(G45), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n715), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n759), .B(new_n765), .C1(G330), .C2(new_n703), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n210), .A2(new_n248), .ZN(new_n767));
  INV_X1    g0567(.A(G355), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n767), .A2(new_n768), .B1(G116), .B2(new_n210), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n714), .A2(new_n248), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n264), .B2(new_n214), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n241), .A2(new_n264), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n769), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT87), .Z(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n215), .B1(G20), .B2(new_n268), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n764), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n207), .A2(new_n411), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n291), .A2(G190), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n207), .A2(new_n330), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n291), .A2(new_n411), .A3(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n784), .A2(G50), .B1(new_n787), .B2(G58), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT88), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n411), .A2(G179), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n316), .B1(new_n792), .B2(G87), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n207), .A2(G190), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n291), .A2(new_n411), .A3(new_n794), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n788), .B1(new_n789), .B2(new_n793), .C1(new_n253), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G179), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G159), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n207), .B1(new_n797), .B2(G190), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n801), .A2(KEYINPUT32), .B1(G97), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n291), .A2(new_n330), .A3(new_n782), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G68), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n793), .A2(new_n789), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT32), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n790), .A2(new_n794), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n800), .A2(new_n809), .B1(new_n811), .B2(G107), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n804), .A2(new_n807), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n795), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G311), .A2(new_n814), .B1(new_n787), .B2(G322), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n784), .A2(G326), .ZN(new_n816));
  XOR2_X1   g0616(.A(KEYINPUT33), .B(G317), .Z(new_n817));
  OAI211_X1 g0617(.A(new_n815), .B(new_n816), .C1(new_n805), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n798), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G283), .A2(new_n811), .B1(new_n819), .B2(G329), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n248), .B1(new_n792), .B2(G303), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(new_n605), .C2(new_n802), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n796), .A2(new_n813), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n781), .B1(new_n823), .B2(new_n778), .ZN(new_n824));
  INV_X1    g0624(.A(new_n777), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n703), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n766), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  NOR2_X1   g0628(.A1(new_n336), .A2(new_n328), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n335), .A2(new_n693), .ZN(new_n830));
  AND3_X1   g0630(.A1(new_n312), .A2(new_n290), .A3(new_n323), .ZN(new_n831));
  AOI21_X1  g0631(.A(G169), .B1(new_n312), .B2(new_n323), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n335), .A2(new_n833), .A3(new_n693), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT91), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n335), .A2(new_n693), .A3(new_n833), .A4(KEYINPUT91), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n829), .A2(new_n830), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(new_n693), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n674), .B2(new_n680), .ZN(new_n840));
  INV_X1    g0640(.A(new_n838), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n739), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n764), .B1(new_n842), .B2(new_n737), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n737), .B2(new_n842), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n778), .A2(new_n775), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n764), .B1(G77), .B2(new_n846), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n473), .A2(new_n795), .B1(new_n783), .B2(new_n488), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(G294), .B2(new_n787), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n316), .B1(new_n791), .B2(new_n317), .ZN(new_n850));
  INV_X1    g0650(.A(G311), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n810), .A2(new_n220), .B1(new_n798), .B2(new_n851), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n850), .B(new_n852), .C1(G97), .C2(new_n803), .ZN(new_n853));
  INV_X1    g0653(.A(G283), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n805), .A2(KEYINPUT89), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n805), .A2(KEYINPUT89), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n849), .B(new_n853), .C1(new_n854), .C2(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n784), .A2(G137), .B1(new_n806), .B2(G150), .ZN(new_n859));
  INV_X1    g0659(.A(G143), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n859), .B1(new_n860), .B2(new_n786), .C1(new_n799), .C2(new_n795), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT34), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n248), .B1(new_n791), .B2(new_n375), .ZN(new_n864));
  INV_X1    g0664(.A(G132), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n810), .A2(new_n202), .B1(new_n798), .B2(new_n865), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n864), .B(new_n866), .C1(G58), .C2(new_n803), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n861), .B2(new_n862), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n858), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n869), .A2(KEYINPUT90), .ZN(new_n870));
  INV_X1    g0670(.A(new_n778), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n869), .B2(KEYINPUT90), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n847), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n776), .B2(new_n841), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n844), .A2(new_n874), .ZN(G384));
  NOR2_X1   g0675(.A1(new_n761), .A2(new_n206), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n445), .A2(KEYINPUT16), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n417), .B1(new_n429), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n690), .A2(new_n691), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n467), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n440), .B1(new_n452), .B2(new_n457), .ZN(new_n884));
  INV_X1    g0684(.A(new_n879), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n452), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n883), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n878), .B1(new_n461), .B2(new_n879), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(KEYINPUT37), .A3(new_n440), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n887), .A2(KEYINPUT38), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n882), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(KEYINPUT92), .B(KEYINPUT38), .Z(new_n893));
  INV_X1    g0693(.A(new_n440), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n451), .A2(new_n271), .A3(new_n428), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n457), .B1(new_n895), .B2(new_n417), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n459), .A2(new_n879), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n897), .A2(KEYINPUT93), .A3(KEYINPUT37), .A4(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT37), .B1(new_n886), .B2(KEYINPUT93), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n459), .A2(new_n461), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n898), .A3(new_n440), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n442), .A2(new_n453), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n898), .B1(new_n463), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n893), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n892), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT94), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n887), .A2(new_n889), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n882), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n890), .B1(new_n467), .B2(new_n881), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT39), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT94), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n892), .A2(new_n907), .A3(new_n915), .A4(new_n908), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n910), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n646), .A2(new_n693), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n463), .A2(new_n879), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n882), .A2(new_n911), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT38), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n913), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n392), .B(new_n693), .C1(new_n393), .C2(new_n399), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n382), .A2(new_n391), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n926), .A2(new_n384), .A3(new_n370), .A4(new_n372), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n392), .A2(new_n693), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n646), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n647), .A2(new_n693), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n931), .B1(new_n840), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n920), .B1(new_n924), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n919), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n756), .B(new_n469), .C1(KEYINPUT29), .C2(new_n739), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n651), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n936), .B(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(G330), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n838), .B1(new_n925), .B2(new_n929), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n721), .B2(new_n736), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n941), .B1(new_n923), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n941), .B1(new_n892), .B2(new_n907), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(KEYINPUT95), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT95), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n942), .B(new_n947), .C1(new_n721), .C2(new_n736), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n944), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n721), .A2(new_n736), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n470), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n940), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n950), .B2(new_n952), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n876), .B1(new_n939), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n939), .B2(new_n954), .ZN(new_n956));
  INV_X1    g0756(.A(new_n548), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(KEYINPUT35), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(KEYINPUT35), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n958), .A2(G116), .A3(new_n216), .A4(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT36), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n213), .A2(new_n253), .A3(new_n422), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n202), .A2(G50), .ZN(new_n963));
  OAI211_X1 g0763(.A(G1), .B(new_n760), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n956), .A2(new_n961), .A3(new_n964), .ZN(G367));
  AOI21_X1  g0765(.A(new_n780), .B1(new_n714), .B2(new_n306), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n770), .A2(new_n237), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n765), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n590), .A2(new_n595), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n693), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n663), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n675), .B2(new_n970), .ZN(new_n972));
  INV_X1    g0772(.A(new_n857), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n814), .A2(G283), .B1(G107), .B2(new_n803), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n973), .A2(G294), .B1(KEYINPUT100), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n791), .A2(new_n473), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT46), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n488), .A2(new_n786), .B1(new_n783), .B2(new_n851), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n810), .A2(new_n225), .ZN(new_n979));
  INV_X1    g0779(.A(G317), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n316), .B1(new_n798), .B2(new_n980), .ZN(new_n981));
  NOR4_X1   g0781(.A1(new_n977), .A2(new_n978), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n975), .B(new_n982), .C1(KEYINPUT100), .C2(new_n974), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n857), .A2(new_n799), .B1(new_n375), .B2(new_n795), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT101), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n810), .A2(new_n253), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G137), .B2(new_n819), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n988), .B(new_n248), .C1(new_n201), .C2(new_n791), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G68), .B2(new_n803), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n784), .A2(G143), .B1(new_n787), .B2(G150), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n986), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n984), .A2(new_n985), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n983), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT47), .Z(new_n995));
  OAI221_X1 g0795(.A(new_n968), .B1(new_n825), .B2(new_n972), .C1(new_n995), .C2(new_n871), .ZN(new_n996));
  INV_X1    g0796(.A(new_n712), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n553), .A2(new_n693), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n749), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n678), .A2(new_n693), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT44), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1001), .B1(KEYINPUT98), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n997), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1002), .A2(KEYINPUT98), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1004), .B(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n712), .A2(new_n1001), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT45), .Z(new_n1009));
  AOI21_X1  g0809(.A(new_n706), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1007), .A2(new_n1009), .A3(new_n706), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT99), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n759), .A2(new_n1014), .ZN(new_n1015));
  MUX2_X1   g0815(.A(new_n697), .B(new_n700), .S(new_n710), .Z(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n759), .A2(new_n1014), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n757), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1013), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n757), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n715), .B(KEYINPUT41), .Z(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n763), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n706), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1001), .B(KEYINPUT96), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT97), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(KEYINPUT97), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1031), .B(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1027), .A2(new_n698), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n693), .B1(new_n1034), .B2(new_n564), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1001), .A2(new_n709), .A3(new_n711), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT42), .Z(new_n1038));
  AOI22_X1  g0838(.A1(new_n1036), .A2(new_n1038), .B1(KEYINPUT43), .B2(new_n972), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1033), .B(new_n1039), .Z(new_n1040));
  OAI21_X1  g0840(.A(new_n996), .B1(new_n1025), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT102), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(G387));
  AOI21_X1  g0843(.A(new_n716), .B1(new_n1019), .B2(new_n757), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n757), .B2(new_n1019), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n264), .B1(new_n202), .B2(new_n253), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n717), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1046), .B1(new_n1047), .B2(KEYINPUT103), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT50), .B1(new_n304), .B2(new_n375), .ZN(new_n1049));
  AND3_X1   g0849(.A1(new_n304), .A2(KEYINPUT50), .A3(new_n375), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1048), .B1(KEYINPUT103), .B2(new_n1047), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n770), .B(new_n1051), .C1(new_n234), .C2(new_n264), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(G107), .B2(new_n210), .C1(new_n717), .C2(new_n767), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n765), .B1(new_n1053), .B2(new_n779), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n700), .B2(new_n825), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n814), .A2(G68), .B1(new_n806), .B2(new_n304), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n784), .A2(G159), .B1(new_n787), .B2(G50), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n791), .A2(new_n253), .B1(new_n798), .B2(new_n273), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n802), .A2(new_n297), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1058), .A2(new_n979), .A3(new_n1059), .A4(new_n316), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1056), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n784), .A2(G322), .B1(new_n787), .B2(G317), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n488), .B2(new_n795), .C1(new_n857), .C2(new_n851), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n792), .A2(G294), .B1(new_n803), .B2(G283), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT49), .Z(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(KEYINPUT104), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n810), .A2(new_n473), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n248), .B(new_n1071), .C1(G326), .C2(new_n819), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1069), .A2(KEYINPUT104), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1061), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1055), .B1(new_n1075), .B2(new_n778), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n1019), .B2(new_n763), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1045), .A2(new_n1077), .ZN(G393));
  NAND2_X1  g0878(.A1(new_n1013), .A2(new_n1020), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1021), .A2(new_n715), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1012), .ZN(new_n1081));
  OAI21_X1  g0881(.A(KEYINPUT105), .B1(new_n1081), .B2(new_n1010), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT105), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1011), .A2(new_n1083), .A3(new_n1012), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n1084), .A3(new_n763), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n779), .B1(new_n225), .B2(new_n210), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n771), .A2(new_n244), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n764), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n851), .A2(new_n786), .B1(new_n783), .B2(new_n980), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT52), .Z(new_n1090));
  AOI22_X1  g0890(.A1(G283), .A2(new_n792), .B1(new_n819), .B2(G322), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1091), .B(new_n316), .C1(new_n317), .C2(new_n810), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G116), .B2(new_n803), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n605), .B2(new_n795), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1090), .B(new_n1094), .C1(G303), .C2(new_n973), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1095), .A2(KEYINPUT106), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(KEYINPUT106), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n802), .A2(new_n253), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G68), .A2(new_n792), .B1(new_n819), .B2(G143), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1099), .B(new_n248), .C1(new_n220), .C2(new_n810), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(new_n304), .C2(new_n814), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n273), .A2(new_n783), .B1(new_n786), .B2(new_n799), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT51), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(new_n375), .C2(new_n857), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1096), .A2(new_n1097), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1088), .B1(new_n1105), .B2(new_n778), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n1027), .B2(new_n825), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1085), .A2(KEYINPUT107), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT107), .B1(new_n1085), .B2(new_n1107), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1080), .B1(new_n1108), .B2(new_n1109), .ZN(G390));
  NAND2_X1  g0910(.A1(new_n469), .A2(new_n738), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n937), .A2(new_n651), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT109), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n937), .A2(KEYINPUT109), .A3(new_n651), .A4(new_n1111), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n564), .A2(new_n742), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1116), .A2(new_n744), .B1(new_n660), .B2(new_n662), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1117), .B(new_n677), .C1(new_n673), .C2(new_n664), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n932), .B1(new_n1118), .B2(new_n839), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n930), .B1(new_n738), .B2(new_n841), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n737), .A2(new_n838), .A3(new_n931), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1122), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n932), .B1(new_n755), .B2(new_n841), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT110), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n838), .B1(new_n737), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n930), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1123), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1114), .A2(new_n1115), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT111), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n918), .B1(new_n892), .B2(new_n907), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1125), .B2(new_n931), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT108), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n934), .B2(new_n918), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n918), .ZN(new_n1139));
  OAI211_X1 g0939(.A(KEYINPUT108), .B(new_n1139), .C1(new_n1119), .C2(new_n931), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1136), .B1(new_n1141), .B2(new_n917), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1122), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1136), .B(new_n1124), .C1(new_n1141), .C2(new_n917), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n716), .B1(new_n1134), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n1145), .B2(new_n1134), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n917), .A2(new_n776), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT54), .B(G143), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n795), .A2(new_n1149), .B1(new_n799), .B2(new_n802), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n973), .B2(G137), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT112), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n316), .B1(new_n819), .B2(G125), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n375), .B2(new_n810), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n792), .A2(G150), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT53), .ZN(new_n1156));
  INV_X1    g0956(.A(G128), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1157), .A2(new_n783), .B1(new_n786), .B2(new_n865), .ZN(new_n1158));
  NOR4_X1   g0958(.A1(new_n1152), .A2(new_n1154), .A3(new_n1156), .A4(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n784), .A2(G283), .B1(new_n814), .B2(G97), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n857), .B2(new_n317), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT113), .Z(new_n1162));
  AOI21_X1  g0962(.A(new_n1098), .B1(new_n787), .B2(G116), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT115), .Z(new_n1164));
  OAI21_X1  g0964(.A(new_n316), .B1(new_n791), .B2(new_n220), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT114), .Z(new_n1166));
  OAI22_X1  g0966(.A1(new_n810), .A2(new_n202), .B1(new_n798), .B2(new_n605), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n1162), .A2(new_n1164), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n778), .B1(new_n1159), .B2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1169), .B(new_n764), .C1(new_n304), .C2(new_n846), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT116), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1145), .A2(new_n763), .B1(new_n1148), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1147), .A2(new_n1172), .ZN(G378));
  INV_X1    g0973(.A(new_n936), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n293), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n643), .A2(new_n644), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n879), .A2(new_n288), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT118), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1181));
  NAND4_X1  g0981(.A1(new_n643), .A2(new_n644), .A3(new_n1175), .A4(new_n1178), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1181), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n944), .A2(new_n949), .A3(G330), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT119), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT120), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n944), .A2(new_n949), .A3(KEYINPUT119), .A4(G330), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1185), .A2(G330), .A3(new_n944), .A4(new_n949), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1188), .A2(new_n1190), .B1(new_n1193), .B2(new_n1189), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1174), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1185), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n1190), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1193), .A2(new_n1189), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n936), .A3(new_n1191), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1143), .A2(new_n1144), .A3(new_n1131), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT121), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1203), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1195), .B(new_n1201), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT57), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(KEYINPUT121), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1202), .A2(new_n1204), .A3(new_n1203), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1200), .A2(new_n936), .A3(new_n1191), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n936), .B1(new_n1200), .B2(new_n1191), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1213), .A2(new_n1216), .A3(KEYINPUT57), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1209), .A2(new_n1217), .A3(new_n715), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n764), .B1(G50), .B2(new_n846), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT117), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n791), .A2(new_n1149), .B1(new_n802), .B2(new_n273), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n784), .A2(G125), .B1(new_n787), .B2(G128), .ZN(new_n1222));
  INV_X1    g1022(.A(G137), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1222), .B1(new_n1223), .B2(new_n795), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1221), .B(new_n1224), .C1(G132), .C2(new_n806), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT59), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n278), .B(new_n263), .C1(new_n810), .C2(new_n799), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G124), .B2(new_n819), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n248), .A2(G41), .ZN(new_n1232));
  AOI211_X1 g1032(.A(G50), .B(new_n1232), .C1(new_n278), .C2(new_n263), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n791), .A2(new_n253), .B1(new_n798), .B2(new_n854), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1232), .B1(new_n201), .B2(new_n810), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(G68), .C2(new_n803), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n784), .A2(G116), .B1(new_n814), .B2(new_n306), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n787), .A2(G107), .B1(new_n806), .B2(G97), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT58), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1233), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1231), .B(new_n1241), .C1(new_n1240), .C2(new_n1239), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1220), .B1(new_n1242), .B2(new_n778), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1185), .B2(new_n776), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1195), .A2(new_n1201), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1244), .B1(new_n1245), .B2(new_n762), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1218), .A2(new_n1247), .ZN(G375));
  NAND2_X1  g1048(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1249), .B(new_n1123), .C1(new_n1130), .C2(new_n1126), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(new_n1024), .A3(new_n1132), .ZN(new_n1251));
  XOR2_X1   g1051(.A(new_n762), .B(KEYINPUT122), .Z(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n931), .A2(new_n775), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n316), .B1(new_n811), .B2(G58), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1256), .A2(KEYINPUT123), .B1(new_n787), .B2(G137), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1257), .B1(new_n865), .B2(new_n783), .C1(new_n273), .C2(new_n795), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(G159), .A2(new_n792), .B1(new_n819), .B2(G128), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1259), .B1(new_n375), .B2(new_n802), .C1(new_n1256), .C2(KEYINPUT123), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n857), .B2(new_n1149), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n317), .A2(new_n795), .B1(new_n783), .B2(new_n605), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(G283), .B2(new_n787), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n791), .A2(new_n225), .B1(new_n798), .B2(new_n488), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(new_n1265), .A2(new_n987), .A3(new_n1059), .A4(new_n248), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1264), .B(new_n1266), .C1(new_n857), .C2(new_n473), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n871), .B1(new_n1262), .B2(new_n1267), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n765), .B(new_n1268), .C1(new_n202), .C2(new_n845), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n1131), .A2(new_n1253), .B1(new_n1254), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1251), .A2(new_n1270), .ZN(G381));
  AND3_X1   g1071(.A1(new_n1045), .A2(new_n827), .A3(new_n1077), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  OR4_X1    g1073(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1273), .ZN(new_n1274));
  OR4_X1    g1074(.A1(G387), .A2(new_n1274), .A3(G378), .A4(G375), .ZN(G407));
  AOI21_X1  g1075(.A(new_n716), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1246), .B1(new_n1276), .B2(new_n1217), .ZN(new_n1277));
  INV_X1    g1077(.A(G378), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n687), .A2(G343), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(G407), .A2(G213), .A3(new_n1280), .ZN(G409));
  AOI21_X1  g1081(.A(new_n827), .B1(new_n1045), .B2(new_n1077), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1272), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G390), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1042), .B1(new_n1272), .B2(new_n1282), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1285), .B(new_n1080), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1284), .A2(new_n1041), .A3(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1041), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1218), .A2(G378), .A3(new_n1247), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1024), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1245), .B1(new_n1292), .B2(new_n1252), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1244), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1278), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1279), .B1(new_n1291), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT60), .ZN(new_n1297));
  OR3_X1    g1097(.A1(new_n1204), .A2(new_n1297), .A3(new_n1131), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1132), .A2(KEYINPUT60), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1250), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1300), .A3(new_n715), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(G384), .B(KEYINPUT124), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(new_n1270), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1279), .A2(G2897), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1301), .A2(new_n1270), .ZN(new_n1305));
  AND2_X1   g1105(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1303), .B(new_n1304), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1304), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1301), .A2(new_n1270), .A3(new_n1302), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1306), .B1(new_n1301), .B2(new_n1270), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1308), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1307), .A2(new_n1311), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1289), .B(new_n1290), .C1(new_n1296), .C2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT125), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1303), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1316));
  AOI211_X1 g1116(.A(new_n1279), .B(new_n1316), .C1(new_n1291), .C2(new_n1295), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1315), .B1(new_n1317), .B2(KEYINPUT63), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(KEYINPUT63), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1279), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1316), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1323), .A2(KEYINPUT125), .A3(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1314), .A2(new_n1318), .A3(new_n1319), .A4(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1289), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1307), .A2(new_n1311), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1023), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1216), .B1(new_n1329), .B2(new_n1253), .ZN(new_n1330));
  AOI21_X1  g1130(.A(G378), .B1(new_n1330), .B2(new_n1244), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1331), .B1(G378), .B2(new_n1277), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1328), .B1(new_n1332), .B2(new_n1279), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT62), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1320), .A2(new_n1334), .A3(new_n1321), .A4(new_n1322), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1333), .A2(new_n1335), .A3(new_n1290), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1317), .A2(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1327), .B1(new_n1336), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1326), .A2(new_n1339), .ZN(G405));
  XNOR2_X1  g1140(.A(new_n1277), .B(new_n1278), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1322), .A2(KEYINPUT127), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1327), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1345), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1347), .A2(new_n1289), .A3(new_n1343), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1346), .A2(new_n1348), .ZN(G402));
endmodule


