

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597;

  XOR2_X1 U326 ( .A(n462), .B(KEYINPUT41), .Z(n569) );
  NOR2_X1 U327 ( .A1(n522), .A2(n513), .ZN(n518) );
  XOR2_X1 U328 ( .A(KEYINPUT28), .B(n483), .Z(n538) );
  XOR2_X1 U329 ( .A(KEYINPUT82), .B(G190GAT), .Z(n294) );
  XNOR2_X2 U330 ( .A(n414), .B(n413), .ZN(n564) );
  XNOR2_X1 U331 ( .A(n477), .B(KEYINPUT48), .ZN(n478) );
  XNOR2_X1 U332 ( .A(n447), .B(KEYINPUT31), .ZN(n448) );
  XNOR2_X1 U333 ( .A(n479), .B(n478), .ZN(n533) );
  XNOR2_X1 U334 ( .A(n393), .B(KEYINPUT97), .ZN(n415) );
  XNOR2_X1 U335 ( .A(n449), .B(n448), .ZN(n451) );
  INV_X1 U336 ( .A(KEYINPUT38), .ZN(n454) );
  XNOR2_X1 U337 ( .A(n454), .B(KEYINPUT99), .ZN(n455) );
  INV_X1 U338 ( .A(n574), .ZN(n575) );
  XOR2_X1 U339 ( .A(n344), .B(n343), .Z(n527) );
  XNOR2_X1 U340 ( .A(n456), .B(n455), .ZN(n511) );
  XNOR2_X1 U341 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U342 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U343 ( .A(n490), .B(n489), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n460), .B(n459), .ZN(G1328GAT) );
  XNOR2_X1 U345 ( .A(KEYINPUT84), .B(KEYINPUT3), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n295), .B(KEYINPUT85), .ZN(n296) );
  XOR2_X1 U347 ( .A(n296), .B(KEYINPUT2), .Z(n298) );
  XNOR2_X1 U348 ( .A(G155GAT), .B(G162GAT), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n298), .B(n297), .ZN(n357) );
  XOR2_X1 U350 ( .A(KEYINPUT88), .B(KEYINPUT90), .Z(n300) );
  XNOR2_X1 U351 ( .A(KEYINPUT89), .B(KEYINPUT6), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U353 ( .A(KEYINPUT1), .B(KEYINPUT87), .Z(n302) );
  XNOR2_X1 U354 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U356 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U357 ( .A(KEYINPUT81), .B(KEYINPUT0), .Z(n306) );
  XNOR2_X1 U358 ( .A(G134GAT), .B(KEYINPUT80), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n321) );
  XNOR2_X1 U360 ( .A(G1GAT), .B(G127GAT), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n307), .B(G57GAT), .ZN(n383) );
  XNOR2_X1 U362 ( .A(n321), .B(n383), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U364 ( .A(G120GAT), .B(G148GAT), .Z(n446) );
  XOR2_X1 U365 ( .A(G113GAT), .B(G141GAT), .Z(n422) );
  XOR2_X1 U366 ( .A(n446), .B(n422), .Z(n311) );
  NAND2_X1 U367 ( .A1(G225GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U369 ( .A(n313), .B(n312), .Z(n315) );
  XNOR2_X1 U370 ( .A(G29GAT), .B(G85GAT), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n357), .B(n316), .ZN(n370) );
  XNOR2_X1 U373 ( .A(KEYINPUT91), .B(n370), .ZN(n523) );
  XNOR2_X1 U374 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n294), .B(n317), .ZN(n318) );
  XNOR2_X1 U376 ( .A(KEYINPUT19), .B(n318), .ZN(n337) );
  XOR2_X1 U377 ( .A(G176GAT), .B(G183GAT), .Z(n320) );
  XNOR2_X1 U378 ( .A(G113GAT), .B(KEYINPUT20), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n331) );
  XOR2_X1 U380 ( .A(G99GAT), .B(n321), .Z(n323) );
  XNOR2_X1 U381 ( .A(G43GAT), .B(G71GAT), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U383 ( .A(n324), .B(G120GAT), .Z(n329) );
  XOR2_X1 U384 ( .A(G127GAT), .B(G15GAT), .Z(n326) );
  NAND2_X1 U385 ( .A1(G227GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U386 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U387 ( .A(G169GAT), .B(n327), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(n337), .B(n332), .Z(n363) );
  XOR2_X1 U391 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n334) );
  NAND2_X1 U392 ( .A1(G226GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U394 ( .A(G204GAT), .B(n335), .ZN(n344) );
  XNOR2_X1 U395 ( .A(G176GAT), .B(G92GAT), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n336), .B(G64GAT), .ZN(n442) );
  XOR2_X1 U397 ( .A(G197GAT), .B(KEYINPUT21), .Z(n350) );
  XOR2_X1 U398 ( .A(n442), .B(n350), .Z(n339) );
  XOR2_X1 U399 ( .A(G169GAT), .B(G8GAT), .Z(n419) );
  XOR2_X1 U400 ( .A(n419), .B(n337), .Z(n338) );
  XNOR2_X1 U401 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U402 ( .A(G183GAT), .B(G211GAT), .Z(n390) );
  XOR2_X1 U403 ( .A(n340), .B(n390), .Z(n342) );
  XNOR2_X1 U404 ( .A(G36GAT), .B(G218GAT), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U406 ( .A(n527), .B(KEYINPUT27), .ZN(n367) );
  NAND2_X1 U407 ( .A1(n523), .A2(n367), .ZN(n534) );
  XOR2_X1 U408 ( .A(G78GAT), .B(KEYINPUT83), .Z(n346) );
  XNOR2_X1 U409 ( .A(G141GAT), .B(KEYINPUT23), .ZN(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n361) );
  XOR2_X1 U411 ( .A(G211GAT), .B(G148GAT), .Z(n348) );
  XNOR2_X1 U412 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U414 ( .A(n349), .B(KEYINPUT22), .Z(n352) );
  XNOR2_X1 U415 ( .A(G50GAT), .B(n350), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U417 ( .A(G106GAT), .B(G204GAT), .Z(n450) );
  XOR2_X1 U418 ( .A(KEYINPUT86), .B(n450), .Z(n354) );
  NAND2_X1 U419 ( .A1(G228GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U420 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U421 ( .A(n356), .B(n355), .Z(n359) );
  XOR2_X1 U422 ( .A(G218GAT), .B(KEYINPUT76), .Z(n410) );
  XNOR2_X1 U423 ( .A(n357), .B(n410), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n483) );
  NOR2_X1 U426 ( .A1(n534), .A2(n538), .ZN(n362) );
  NAND2_X1 U427 ( .A1(n363), .A2(n362), .ZN(n373) );
  INV_X1 U428 ( .A(n363), .ZN(n536) );
  NAND2_X1 U429 ( .A1(n536), .A2(n527), .ZN(n364) );
  NAND2_X1 U430 ( .A1(n483), .A2(n364), .ZN(n365) );
  XOR2_X1 U431 ( .A(KEYINPUT25), .B(n365), .Z(n369) );
  NOR2_X1 U432 ( .A1(n483), .A2(n536), .ZN(n366) );
  XNOR2_X1 U433 ( .A(n366), .B(KEYINPUT26), .ZN(n581) );
  NAND2_X1 U434 ( .A1(n367), .A2(n581), .ZN(n368) );
  NAND2_X1 U435 ( .A1(n369), .A2(n368), .ZN(n371) );
  NAND2_X1 U436 ( .A1(n371), .A2(n370), .ZN(n372) );
  NAND2_X1 U437 ( .A1(n373), .A2(n372), .ZN(n493) );
  XOR2_X1 U438 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n375) );
  NAND2_X1 U439 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U440 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U441 ( .A(n376), .B(KEYINPUT15), .Z(n385) );
  INV_X1 U442 ( .A(KEYINPUT13), .ZN(n377) );
  NAND2_X1 U443 ( .A1(KEYINPUT74), .A2(n377), .ZN(n380) );
  INV_X1 U444 ( .A(KEYINPUT74), .ZN(n378) );
  NAND2_X1 U445 ( .A1(n378), .A2(KEYINPUT13), .ZN(n379) );
  NAND2_X1 U446 ( .A1(n380), .A2(n379), .ZN(n382) );
  XNOR2_X1 U447 ( .A(G71GAT), .B(G78GAT), .ZN(n381) );
  XNOR2_X1 U448 ( .A(n382), .B(n381), .ZN(n443) );
  XNOR2_X1 U449 ( .A(n383), .B(n443), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U451 ( .A(KEYINPUT12), .B(G64GAT), .Z(n387) );
  XNOR2_X1 U452 ( .A(G8GAT), .B(G155GAT), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U454 ( .A(n389), .B(n388), .Z(n392) );
  XOR2_X1 U455 ( .A(G15GAT), .B(G22GAT), .Z(n418) );
  XNOR2_X1 U456 ( .A(n418), .B(n390), .ZN(n391) );
  XNOR2_X1 U457 ( .A(n392), .B(n391), .ZN(n560) );
  INV_X1 U458 ( .A(n560), .ZN(n592) );
  NAND2_X1 U459 ( .A1(n493), .A2(n592), .ZN(n393) );
  XOR2_X1 U460 ( .A(KEYINPUT66), .B(KEYINPUT65), .Z(n395) );
  XNOR2_X1 U461 ( .A(G190GAT), .B(G92GAT), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n414) );
  XOR2_X1 U463 ( .A(KEYINPUT10), .B(KEYINPUT68), .Z(n397) );
  XNOR2_X1 U464 ( .A(G162GAT), .B(G106GAT), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n397), .B(n396), .ZN(n399) );
  INV_X1 U466 ( .A(KEYINPUT11), .ZN(n398) );
  XNOR2_X1 U467 ( .A(n399), .B(n398), .ZN(n401) );
  XNOR2_X1 U468 ( .A(G99GAT), .B(G85GAT), .ZN(n452) );
  XOR2_X1 U469 ( .A(G134GAT), .B(n452), .Z(n400) );
  XNOR2_X1 U470 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U471 ( .A(KEYINPUT77), .B(KEYINPUT9), .Z(n403) );
  NAND2_X1 U472 ( .A1(G232GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U473 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U474 ( .A(n405), .B(n404), .Z(n412) );
  XNOR2_X1 U475 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n406) );
  XNOR2_X1 U476 ( .A(n406), .B(G29GAT), .ZN(n407) );
  XOR2_X1 U477 ( .A(n407), .B(KEYINPUT8), .Z(n409) );
  XNOR2_X1 U478 ( .A(G43GAT), .B(G50GAT), .ZN(n408) );
  XNOR2_X1 U479 ( .A(n409), .B(n408), .ZN(n433) );
  XNOR2_X1 U480 ( .A(n433), .B(n410), .ZN(n411) );
  XNOR2_X1 U481 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U482 ( .A(KEYINPUT36), .B(n564), .ZN(n468) );
  NAND2_X1 U483 ( .A1(n415), .A2(n468), .ZN(n417) );
  XOR2_X1 U484 ( .A(KEYINPUT98), .B(KEYINPUT37), .Z(n416) );
  XNOR2_X1 U485 ( .A(n417), .B(n416), .ZN(n521) );
  XOR2_X1 U486 ( .A(n419), .B(n418), .Z(n421) );
  NAND2_X1 U487 ( .A1(G229GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U488 ( .A(n421), .B(n420), .ZN(n423) );
  XOR2_X1 U489 ( .A(n423), .B(n422), .Z(n431) );
  XOR2_X1 U490 ( .A(KEYINPUT30), .B(KEYINPUT71), .Z(n425) );
  XNOR2_X1 U491 ( .A(G197GAT), .B(G1GAT), .ZN(n424) );
  XNOR2_X1 U492 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U493 ( .A(KEYINPUT69), .B(KEYINPUT72), .Z(n427) );
  XNOR2_X1 U494 ( .A(KEYINPUT70), .B(KEYINPUT29), .ZN(n426) );
  XNOR2_X1 U495 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U496 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U498 ( .A(n433), .B(n432), .Z(n554) );
  XOR2_X1 U499 ( .A(KEYINPUT73), .B(n554), .Z(n567) );
  INV_X1 U500 ( .A(KEYINPUT33), .ZN(n434) );
  NAND2_X1 U501 ( .A1(KEYINPUT75), .A2(n434), .ZN(n437) );
  INV_X1 U502 ( .A(KEYINPUT75), .ZN(n435) );
  NAND2_X1 U503 ( .A1(n435), .A2(KEYINPUT33), .ZN(n436) );
  NAND2_X1 U504 ( .A1(n437), .A2(n436), .ZN(n439) );
  NAND2_X1 U505 ( .A1(G230GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U506 ( .A(n439), .B(n438), .ZN(n441) );
  INV_X1 U507 ( .A(KEYINPUT32), .ZN(n440) );
  XNOR2_X1 U508 ( .A(n441), .B(n440), .ZN(n445) );
  XNOR2_X1 U509 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U510 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U511 ( .A(G57GAT), .B(n446), .Z(n447) );
  XNOR2_X1 U512 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n453), .B(n452), .ZN(n461) );
  NAND2_X1 U514 ( .A1(n567), .A2(n461), .ZN(n495) );
  NOR2_X1 U515 ( .A1(n521), .A2(n495), .ZN(n456) );
  NAND2_X1 U516 ( .A1(n523), .A2(n511), .ZN(n460) );
  XOR2_X1 U517 ( .A(G29GAT), .B(KEYINPUT100), .Z(n458) );
  XOR2_X1 U518 ( .A(KEYINPUT39), .B(KEYINPUT101), .Z(n457) );
  INV_X1 U519 ( .A(n461), .ZN(n462) );
  NAND2_X1 U520 ( .A1(n554), .A2(n569), .ZN(n463) );
  XNOR2_X1 U521 ( .A(KEYINPUT46), .B(n463), .ZN(n464) );
  XNOR2_X1 U522 ( .A(KEYINPUT106), .B(n592), .ZN(n576) );
  NAND2_X1 U523 ( .A1(n464), .A2(n576), .ZN(n465) );
  NOR2_X1 U524 ( .A1(n465), .A2(n564), .ZN(n467) );
  INV_X1 U525 ( .A(KEYINPUT47), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n467), .B(n466), .ZN(n476) );
  NAND2_X1 U527 ( .A1(n468), .A2(n560), .ZN(n470) );
  XNOR2_X1 U528 ( .A(KEYINPUT67), .B(KEYINPUT45), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n470), .B(n469), .ZN(n471) );
  AND2_X1 U530 ( .A1(n471), .A2(n461), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n472), .B(KEYINPUT107), .ZN(n473) );
  NOR2_X1 U532 ( .A1(n567), .A2(n473), .ZN(n474) );
  XNOR2_X1 U533 ( .A(KEYINPUT108), .B(n474), .ZN(n475) );
  NOR2_X1 U534 ( .A1(n476), .A2(n475), .ZN(n479) );
  XOR2_X1 U535 ( .A(KEYINPUT64), .B(KEYINPUT109), .Z(n477) );
  INV_X1 U536 ( .A(n527), .ZN(n480) );
  NOR2_X1 U537 ( .A1(n533), .A2(n480), .ZN(n481) );
  XOR2_X1 U538 ( .A(KEYINPUT54), .B(n481), .Z(n482) );
  NOR2_X1 U539 ( .A1(n523), .A2(n482), .ZN(n582) );
  NAND2_X1 U540 ( .A1(n582), .A2(n483), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n484), .B(KEYINPUT55), .ZN(n485) );
  NAND2_X1 U542 ( .A1(n485), .A2(n536), .ZN(n486) );
  XNOR2_X2 U543 ( .A(n486), .B(KEYINPUT119), .ZN(n574) );
  NAND2_X1 U544 ( .A1(n574), .A2(n564), .ZN(n490) );
  XOR2_X1 U545 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n488) );
  INV_X1 U546 ( .A(G190GAT), .ZN(n487) );
  NOR2_X1 U547 ( .A1(n564), .A2(n592), .ZN(n491) );
  XOR2_X1 U548 ( .A(KEYINPUT79), .B(n491), .Z(n492) );
  XNOR2_X1 U549 ( .A(n492), .B(KEYINPUT16), .ZN(n494) );
  NAND2_X1 U550 ( .A1(n494), .A2(n493), .ZN(n513) );
  NOR2_X1 U551 ( .A1(n495), .A2(n513), .ZN(n503) );
  NAND2_X1 U552 ( .A1(n503), .A2(n523), .ZN(n496) );
  XNOR2_X1 U553 ( .A(n496), .B(KEYINPUT34), .ZN(n497) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(n497), .ZN(G1324GAT) );
  NAND2_X1 U555 ( .A1(n527), .A2(n503), .ZN(n498) );
  XNOR2_X1 U556 ( .A(n498), .B(KEYINPUT94), .ZN(n499) );
  XNOR2_X1 U557 ( .A(G8GAT), .B(n499), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT95), .B(KEYINPUT35), .Z(n501) );
  NAND2_X1 U559 ( .A1(n503), .A2(n536), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U561 ( .A(G15GAT), .B(n502), .Z(G1326GAT) );
  NAND2_X1 U562 ( .A1(n538), .A2(n503), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n504), .B(KEYINPUT96), .ZN(n505) );
  XNOR2_X1 U564 ( .A(G22GAT), .B(n505), .ZN(G1327GAT) );
  NAND2_X1 U565 ( .A1(n511), .A2(n527), .ZN(n506) );
  XNOR2_X1 U566 ( .A(n506), .B(KEYINPUT102), .ZN(n507) );
  XNOR2_X1 U567 ( .A(G36GAT), .B(n507), .ZN(G1329GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n509) );
  NAND2_X1 U569 ( .A1(n511), .A2(n536), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U571 ( .A(G43GAT), .B(n510), .ZN(G1330GAT) );
  NAND2_X1 U572 ( .A1(n511), .A2(n538), .ZN(n512) );
  XNOR2_X1 U573 ( .A(n512), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n515) );
  INV_X1 U575 ( .A(n554), .ZN(n583) );
  NAND2_X1 U576 ( .A1(n569), .A2(n583), .ZN(n522) );
  NAND2_X1 U577 ( .A1(n523), .A2(n518), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n515), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U579 ( .A1(n527), .A2(n518), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n516), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n536), .A2(n518), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U584 ( .A1(n518), .A2(n538), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n525) );
  NOR2_X1 U587 ( .A1(n521), .A2(n522), .ZN(n530) );
  NAND2_X1 U588 ( .A1(n530), .A2(n523), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(n526), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n527), .A2(n530), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n536), .A2(n530), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n529), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U595 ( .A1(n538), .A2(n530), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(KEYINPUT110), .ZN(n552) );
  NAND2_X1 U600 ( .A1(n536), .A2(n552), .ZN(n537) );
  NOR2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n548), .A2(n567), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n539), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U605 ( .A1(n548), .A2(n569), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U607 ( .A(G120GAT), .B(n542), .Z(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT112), .Z(n544) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(KEYINPUT113), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n547) );
  INV_X1 U611 ( .A(n548), .ZN(n545) );
  NOR2_X1 U612 ( .A1(n576), .A2(n545), .ZN(n546) );
  XOR2_X1 U613 ( .A(n547), .B(n546), .Z(G1342GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U615 ( .A1(n548), .A2(n564), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G134GAT), .B(n551), .ZN(G1343GAT) );
  NAND2_X1 U618 ( .A1(n552), .A2(n581), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(KEYINPUT115), .ZN(n563) );
  NAND2_X1 U620 ( .A1(n563), .A2(n554), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n559) );
  XOR2_X1 U623 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U624 ( .A1(n563), .A2(n569), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  XOR2_X1 U627 ( .A(G155GAT), .B(KEYINPUT117), .Z(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n560), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1346GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT118), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G162GAT), .B(n566), .ZN(G1347GAT) );
  NAND2_X1 U633 ( .A1(n574), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U635 ( .A1(n574), .A2(n569), .ZN(n571) );
  XOR2_X1 U636 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1349GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U641 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1350GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n580) );
  XNOR2_X1 U644 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n587) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n594) );
  NOR2_X1 U647 ( .A1(n583), .A2(n594), .ZN(n585) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(n587), .B(n586), .Z(G1352GAT) );
  NOR2_X1 U651 ( .A1(n594), .A2(n461), .ZN(n591) );
  XOR2_X1 U652 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n589) );
  XNOR2_X1 U653 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(G1353GAT) );
  NOR2_X1 U656 ( .A1(n592), .A2(n594), .ZN(n593) );
  XOR2_X1 U657 ( .A(G211GAT), .B(n593), .Z(G1354GAT) );
  INV_X1 U658 ( .A(n594), .ZN(n595) );
  NAND2_X1 U659 ( .A1(n595), .A2(n468), .ZN(n596) );
  XNOR2_X1 U660 ( .A(n596), .B(KEYINPUT62), .ZN(n597) );
  XNOR2_X1 U661 ( .A(G218GAT), .B(n597), .ZN(G1355GAT) );
endmodule

