

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583;

  XNOR2_X2 U324 ( .A(n413), .B(KEYINPUT48), .ZN(n545) );
  NOR2_X1 U325 ( .A1(n561), .A2(n405), .ZN(n406) );
  XNOR2_X1 U326 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U327 ( .A(n385), .B(n384), .ZN(n573) );
  XNOR2_X1 U328 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U329 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT83), .B(KEYINPUT0), .Z(n293) );
  XNOR2_X1 U331 ( .A(G113GAT), .B(KEYINPUT82), .ZN(n292) );
  XNOR2_X1 U332 ( .A(n293), .B(n292), .ZN(n325) );
  XOR2_X1 U333 ( .A(n325), .B(G134GAT), .Z(n295) );
  NAND2_X1 U334 ( .A1(G227GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U335 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U336 ( .A(n296), .B(G190GAT), .Z(n304) );
  XOR2_X1 U337 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n298) );
  XNOR2_X1 U338 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n297) );
  XNOR2_X1 U339 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U340 ( .A(G169GAT), .B(n299), .Z(n424) );
  XOR2_X1 U341 ( .A(G127GAT), .B(G183GAT), .Z(n301) );
  XNOR2_X1 U342 ( .A(KEYINPUT87), .B(KEYINPUT86), .ZN(n300) );
  XNOR2_X1 U343 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U344 ( .A(n424), .B(n302), .ZN(n303) );
  XNOR2_X1 U345 ( .A(n304), .B(n303), .ZN(n312) );
  XOR2_X1 U346 ( .A(KEYINPUT84), .B(G71GAT), .Z(n306) );
  XNOR2_X1 U347 ( .A(KEYINPUT20), .B(G176GAT), .ZN(n305) );
  XNOR2_X1 U348 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U349 ( .A(G120GAT), .B(G99GAT), .Z(n308) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(G15GAT), .ZN(n307) );
  XNOR2_X1 U351 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U352 ( .A(n310), .B(n309), .Z(n311) );
  XOR2_X1 U353 ( .A(n312), .B(n311), .Z(n529) );
  INV_X1 U354 ( .A(n529), .ZN(n522) );
  XOR2_X1 U355 ( .A(KEYINPUT97), .B(KEYINPUT1), .Z(n314) );
  XNOR2_X1 U356 ( .A(G155GAT), .B(G85GAT), .ZN(n313) );
  XNOR2_X1 U357 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U358 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n316) );
  XNOR2_X1 U359 ( .A(KEYINPUT4), .B(KEYINPUT96), .ZN(n315) );
  XNOR2_X1 U360 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U361 ( .A(n318), .B(n317), .Z(n323) );
  XOR2_X1 U362 ( .A(G29GAT), .B(G134GAT), .Z(n338) );
  XOR2_X1 U363 ( .A(G120GAT), .B(G148GAT), .Z(n371) );
  XOR2_X1 U364 ( .A(G1GAT), .B(G127GAT), .Z(n351) );
  XOR2_X1 U365 ( .A(n371), .B(n351), .Z(n320) );
  NAND2_X1 U366 ( .A1(G225GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U368 ( .A(n338), .B(n321), .ZN(n322) );
  XNOR2_X1 U369 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U370 ( .A(n324), .B(G57GAT), .Z(n327) );
  XNOR2_X1 U371 ( .A(n325), .B(KEYINPUT98), .ZN(n326) );
  XNOR2_X1 U372 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U373 ( .A(KEYINPUT92), .B(G162GAT), .Z(n329) );
  XNOR2_X1 U374 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n328) );
  XNOR2_X1 U375 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U376 ( .A(G141GAT), .B(n330), .Z(n434) );
  XOR2_X1 U377 ( .A(n331), .B(n434), .Z(n468) );
  XNOR2_X1 U378 ( .A(KEYINPUT99), .B(n468), .ZN(n517) );
  XOR2_X1 U379 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n333) );
  XNOR2_X1 U380 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n332) );
  XNOR2_X1 U381 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U382 ( .A(G99GAT), .B(G85GAT), .Z(n366) );
  XOR2_X1 U383 ( .A(n334), .B(n366), .Z(n336) );
  XNOR2_X1 U384 ( .A(G218GAT), .B(G106GAT), .ZN(n335) );
  XNOR2_X1 U385 ( .A(n336), .B(n335), .ZN(n342) );
  XNOR2_X1 U386 ( .A(G36GAT), .B(G190GAT), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n337), .B(KEYINPUT77), .ZN(n418) );
  XOR2_X1 U388 ( .A(n418), .B(n338), .Z(n340) );
  NAND2_X1 U389 ( .A1(G232GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U391 ( .A(n342), .B(n341), .Z(n350) );
  XOR2_X1 U392 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n344) );
  XNOR2_X1 U393 ( .A(G50GAT), .B(G43GAT), .ZN(n343) );
  XNOR2_X1 U394 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U395 ( .A(KEYINPUT70), .B(n345), .Z(n395) );
  XOR2_X1 U396 ( .A(KEYINPUT78), .B(KEYINPUT65), .Z(n347) );
  XNOR2_X1 U397 ( .A(G162GAT), .B(KEYINPUT67), .ZN(n346) );
  XNOR2_X1 U398 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U399 ( .A(n395), .B(n348), .ZN(n349) );
  XNOR2_X1 U400 ( .A(n350), .B(n349), .ZN(n561) );
  XNOR2_X1 U401 ( .A(G15GAT), .B(n351), .ZN(n352) );
  XNOR2_X1 U402 ( .A(n352), .B(G64GAT), .ZN(n365) );
  XNOR2_X1 U403 ( .A(G22GAT), .B(G155GAT), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n353), .B(G78GAT), .ZN(n436) );
  XOR2_X1 U405 ( .A(KEYINPUT80), .B(n436), .Z(n355) );
  NAND2_X1 U406 ( .A1(G231GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U407 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U408 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n357) );
  XNOR2_X1 U409 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U411 ( .A(n359), .B(n358), .Z(n363) );
  XNOR2_X1 U412 ( .A(G8GAT), .B(G183GAT), .ZN(n360) );
  XNOR2_X1 U413 ( .A(n360), .B(G211GAT), .ZN(n421) );
  XNOR2_X1 U414 ( .A(G71GAT), .B(G57GAT), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n361), .B(KEYINPUT13), .ZN(n367) );
  XNOR2_X1 U416 ( .A(n421), .B(n367), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U418 ( .A(n365), .B(n364), .Z(n552) );
  XOR2_X1 U419 ( .A(KEYINPUT116), .B(n552), .Z(n558) );
  XNOR2_X1 U420 ( .A(n367), .B(n366), .ZN(n369) );
  AND2_X1 U421 ( .A1(G230GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U423 ( .A(n370), .B(G78GAT), .ZN(n376) );
  XOR2_X1 U424 ( .A(KEYINPUT71), .B(KEYINPUT31), .Z(n373) );
  XOR2_X1 U425 ( .A(G106GAT), .B(KEYINPUT73), .Z(n442) );
  XNOR2_X1 U426 ( .A(n442), .B(n371), .ZN(n372) );
  XOR2_X1 U427 ( .A(n373), .B(n372), .Z(n374) );
  XNOR2_X1 U428 ( .A(n374), .B(KEYINPUT76), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n376), .B(n375), .ZN(n385) );
  XOR2_X1 U430 ( .A(G92GAT), .B(G64GAT), .Z(n378) );
  XNOR2_X1 U431 ( .A(G176GAT), .B(KEYINPUT75), .ZN(n377) );
  XNOR2_X1 U432 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U433 ( .A(G204GAT), .B(n379), .ZN(n423) );
  INV_X1 U434 ( .A(n423), .ZN(n383) );
  XOR2_X1 U435 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n381) );
  XNOR2_X1 U436 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U438 ( .A(n573), .B(KEYINPUT41), .Z(n453) );
  XOR2_X1 U439 ( .A(G8GAT), .B(G1GAT), .Z(n387) );
  XNOR2_X1 U440 ( .A(G141GAT), .B(G197GAT), .ZN(n386) );
  XNOR2_X1 U441 ( .A(n387), .B(n386), .ZN(n401) );
  NAND2_X1 U442 ( .A1(G229GAT), .A2(G233GAT), .ZN(n393) );
  XOR2_X1 U443 ( .A(G22GAT), .B(G113GAT), .Z(n389) );
  XNOR2_X1 U444 ( .A(G169GAT), .B(G15GAT), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n391) );
  XOR2_X1 U446 ( .A(G36GAT), .B(G29GAT), .Z(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U448 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U450 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n397) );
  XNOR2_X1 U451 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n396) );
  XNOR2_X1 U452 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U453 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U454 ( .A(n401), .B(n400), .Z(n458) );
  INV_X1 U455 ( .A(n458), .ZN(n570) );
  AND2_X1 U456 ( .A1(n453), .A2(n570), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n402), .B(KEYINPUT46), .ZN(n403) );
  NOR2_X1 U458 ( .A1(n558), .A2(n403), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n404), .B(KEYINPUT117), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n406), .B(KEYINPUT47), .ZN(n412) );
  XNOR2_X1 U461 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n408) );
  XOR2_X1 U462 ( .A(KEYINPUT36), .B(n561), .Z(n580) );
  NOR2_X1 U463 ( .A1(n580), .A2(n552), .ZN(n407) );
  XOR2_X1 U464 ( .A(n408), .B(n407), .Z(n409) );
  NOR2_X1 U465 ( .A1(n573), .A2(n409), .ZN(n410) );
  NAND2_X1 U466 ( .A1(n410), .A2(n458), .ZN(n411) );
  NAND2_X1 U467 ( .A1(n412), .A2(n411), .ZN(n413) );
  XNOR2_X1 U468 ( .A(KEYINPUT89), .B(KEYINPUT21), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n414), .B(KEYINPUT90), .ZN(n415) );
  XOR2_X1 U470 ( .A(n415), .B(KEYINPUT91), .Z(n417) );
  XNOR2_X1 U471 ( .A(G197GAT), .B(G218GAT), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n450) );
  XOR2_X1 U473 ( .A(KEYINPUT100), .B(n418), .Z(n420) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U476 ( .A(n422), .B(n421), .Z(n426) );
  XOR2_X1 U477 ( .A(n424), .B(n423), .Z(n425) );
  XNOR2_X1 U478 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U479 ( .A(n450), .B(n427), .Z(n519) );
  INV_X1 U480 ( .A(n519), .ZN(n459) );
  NAND2_X1 U481 ( .A1(n545), .A2(n459), .ZN(n429) );
  XOR2_X1 U482 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n430) );
  NAND2_X1 U484 ( .A1(n517), .A2(n430), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n431), .B(KEYINPUT64), .ZN(n569) );
  XOR2_X1 U486 ( .A(G211GAT), .B(G148GAT), .Z(n433) );
  XNOR2_X1 U487 ( .A(KEYINPUT94), .B(KEYINPUT88), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U489 ( .A(n435), .B(n434), .Z(n448) );
  XOR2_X1 U490 ( .A(KEYINPUT95), .B(n436), .Z(n438) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n446) );
  XOR2_X1 U493 ( .A(G204GAT), .B(KEYINPUT23), .Z(n440) );
  XNOR2_X1 U494 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U496 ( .A(n441), .B(KEYINPUT93), .Z(n444) );
  XNOR2_X1 U497 ( .A(G50GAT), .B(n442), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n471) );
  NOR2_X1 U502 ( .A1(n569), .A2(n471), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n451), .B(KEYINPUT55), .ZN(n452) );
  NOR2_X2 U504 ( .A1(n522), .A2(n452), .ZN(n562) );
  INV_X1 U505 ( .A(n453), .ZN(n502) );
  INV_X1 U506 ( .A(n502), .ZN(n548) );
  NAND2_X1 U507 ( .A1(n562), .A2(n548), .ZN(n457) );
  XOR2_X1 U508 ( .A(G176GAT), .B(KEYINPUT124), .Z(n455) );
  XNOR2_X1 U509 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n454) );
  NOR2_X1 U510 ( .A1(n573), .A2(n458), .ZN(n490) );
  NAND2_X1 U511 ( .A1(n529), .A2(n459), .ZN(n460) );
  XOR2_X1 U512 ( .A(KEYINPUT102), .B(n460), .Z(n461) );
  NOR2_X1 U513 ( .A1(n471), .A2(n461), .ZN(n463) );
  XNOR2_X1 U514 ( .A(KEYINPUT103), .B(KEYINPUT25), .ZN(n462) );
  XNOR2_X1 U515 ( .A(n463), .B(n462), .ZN(n466) );
  XNOR2_X1 U516 ( .A(KEYINPUT27), .B(n519), .ZN(n469) );
  NAND2_X1 U517 ( .A1(n471), .A2(n522), .ZN(n464) );
  XNOR2_X1 U518 ( .A(n464), .B(KEYINPUT26), .ZN(n568) );
  NOR2_X1 U519 ( .A1(n469), .A2(n568), .ZN(n465) );
  NOR2_X1 U520 ( .A1(n466), .A2(n465), .ZN(n467) );
  NOR2_X1 U521 ( .A1(n468), .A2(n467), .ZN(n473) );
  NOR2_X1 U522 ( .A1(n517), .A2(n469), .ZN(n470) );
  XOR2_X1 U523 ( .A(KEYINPUT101), .B(n470), .Z(n544) );
  XOR2_X1 U524 ( .A(KEYINPUT28), .B(n471), .Z(n526) );
  NAND2_X1 U525 ( .A1(n544), .A2(n526), .ZN(n531) );
  NOR2_X1 U526 ( .A1(n529), .A2(n531), .ZN(n472) );
  NOR2_X1 U527 ( .A1(n473), .A2(n472), .ZN(n486) );
  XNOR2_X1 U528 ( .A(KEYINPUT16), .B(KEYINPUT81), .ZN(n475) );
  NOR2_X1 U529 ( .A1(n561), .A2(n552), .ZN(n474) );
  XNOR2_X1 U530 ( .A(n475), .B(n474), .ZN(n476) );
  NOR2_X1 U531 ( .A1(n486), .A2(n476), .ZN(n503) );
  NAND2_X1 U532 ( .A1(n490), .A2(n503), .ZN(n484) );
  NOR2_X1 U533 ( .A1(n517), .A2(n484), .ZN(n478) );
  XNOR2_X1 U534 ( .A(KEYINPUT34), .B(KEYINPUT104), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U536 ( .A(G1GAT), .B(n479), .Z(G1324GAT) );
  NOR2_X1 U537 ( .A1(n519), .A2(n484), .ZN(n481) );
  XNOR2_X1 U538 ( .A(G8GAT), .B(KEYINPUT105), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(G1325GAT) );
  NOR2_X1 U540 ( .A1(n522), .A2(n484), .ZN(n483) );
  XNOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U543 ( .A1(n526), .A2(n484), .ZN(n485) );
  XOR2_X1 U544 ( .A(G22GAT), .B(n485), .Z(G1327GAT) );
  NOR2_X1 U545 ( .A1(n580), .A2(n486), .ZN(n487) );
  NAND2_X1 U546 ( .A1(n552), .A2(n487), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT37), .B(n488), .ZN(n489) );
  XNOR2_X1 U548 ( .A(KEYINPUT106), .B(n489), .ZN(n515) );
  NAND2_X1 U549 ( .A1(n515), .A2(n490), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n491), .B(KEYINPUT38), .ZN(n499) );
  NOR2_X1 U551 ( .A1(n499), .A2(n517), .ZN(n493) );
  XNOR2_X1 U552 ( .A(KEYINPUT39), .B(KEYINPUT107), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U554 ( .A(G29GAT), .B(n494), .Z(G1328GAT) );
  NOR2_X1 U555 ( .A1(n519), .A2(n499), .ZN(n495) );
  XOR2_X1 U556 ( .A(G36GAT), .B(n495), .Z(G1329GAT) );
  NOR2_X1 U557 ( .A1(n499), .A2(n522), .ZN(n497) );
  XNOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT108), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U560 ( .A(G43GAT), .B(n498), .Z(G1330GAT) );
  NOR2_X1 U561 ( .A1(n499), .A2(n526), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(KEYINPUT109), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(G1331GAT) );
  NOR2_X1 U564 ( .A1(n570), .A2(n502), .ZN(n516) );
  NAND2_X1 U565 ( .A1(n516), .A2(n503), .ZN(n511) );
  NOR2_X1 U566 ( .A1(n517), .A2(n511), .ZN(n504) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n504), .Z(n505) );
  XNOR2_X1 U568 ( .A(KEYINPUT42), .B(n505), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n519), .A2(n511), .ZN(n507) );
  XNOR2_X1 U570 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U573 ( .A1(n522), .A2(n511), .ZN(n509) );
  XOR2_X1 U574 ( .A(KEYINPUT112), .B(n509), .Z(n510) );
  XNOR2_X1 U575 ( .A(G71GAT), .B(n510), .ZN(G1334GAT) );
  NOR2_X1 U576 ( .A1(n526), .A2(n511), .ZN(n513) );
  XNOR2_X1 U577 ( .A(KEYINPUT43), .B(KEYINPUT113), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U579 ( .A(G78GAT), .B(n514), .Z(G1335GAT) );
  NAND2_X1 U580 ( .A1(n516), .A2(n515), .ZN(n525) );
  NOR2_X1 U581 ( .A1(n517), .A2(n525), .ZN(n518) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n518), .Z(G1336GAT) );
  NOR2_X1 U583 ( .A1(n519), .A2(n525), .ZN(n520) );
  XOR2_X1 U584 ( .A(KEYINPUT114), .B(n520), .Z(n521) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n521), .ZN(G1337GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n525), .ZN(n524) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(KEYINPUT115), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(G1338GAT) );
  NOR2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(n527), .Z(n528) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NAND2_X1 U592 ( .A1(n529), .A2(n545), .ZN(n530) );
  NOR2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n540), .A2(n570), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n532), .B(KEYINPUT118), .ZN(n533) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U598 ( .A1(n540), .A2(n548), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U600 ( .A(G120GAT), .B(n536), .Z(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT120), .B(KEYINPUT50), .Z(n538) );
  NAND2_X1 U602 ( .A1(n540), .A2(n558), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U604 ( .A(G127GAT), .B(n539), .Z(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT51), .B(KEYINPUT121), .Z(n542) );
  NAND2_X1 U606 ( .A1(n540), .A2(n561), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U608 ( .A(G134GAT), .B(n543), .Z(G1343GAT) );
  NAND2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U610 ( .A1(n568), .A2(n546), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n554), .A2(n570), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n547), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  NAND2_X1 U614 ( .A1(n554), .A2(n548), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  INV_X1 U617 ( .A(n552), .ZN(n576) );
  NAND2_X1 U618 ( .A1(n576), .A2(n554), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n554), .A2(n561), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U622 ( .A(G169GAT), .B(KEYINPUT123), .Z(n557) );
  NAND2_X1 U623 ( .A1(n562), .A2(n570), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(G183GAT), .B(KEYINPUT125), .Z(n560) );
  NAND2_X1 U626 ( .A1(n562), .A2(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1350GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT58), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n566) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT126), .B(n567), .Z(n572) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n578) );
  NAND2_X1 U636 ( .A1(n578), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U639 ( .A1(n578), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n578), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U643 ( .A(KEYINPUT62), .ZN(n582) );
  INV_X1 U644 ( .A(n578), .ZN(n579) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

