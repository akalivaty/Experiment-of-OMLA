

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U325 ( .A(n458), .B(n457), .ZN(n471) );
  NOR2_X2 U326 ( .A1(n521), .A2(n479), .ZN(n570) );
  XNOR2_X1 U327 ( .A(n411), .B(KEYINPUT99), .ZN(n417) );
  XNOR2_X1 U328 ( .A(n326), .B(n325), .ZN(n330) );
  OR2_X1 U329 ( .A1(n520), .A2(n493), .ZN(n459) );
  XOR2_X1 U330 ( .A(n480), .B(KEYINPUT28), .Z(n533) );
  AND2_X1 U331 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U332 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n294) );
  XOR2_X1 U333 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n295) );
  INV_X1 U334 ( .A(KEYINPUT45), .ZN(n469) );
  XNOR2_X1 U335 ( .A(n470), .B(n469), .ZN(n472) );
  XNOR2_X1 U336 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U337 ( .A(n392), .B(n391), .ZN(n394) );
  INV_X1 U338 ( .A(KEYINPUT102), .ZN(n422) );
  XNOR2_X1 U339 ( .A(n324), .B(n293), .ZN(n325) );
  XNOR2_X1 U340 ( .A(n423), .B(n422), .ZN(n424) );
  NOR2_X1 U341 ( .A1(n480), .A2(n530), .ZN(n409) );
  XOR2_X1 U342 ( .A(KEYINPUT36), .B(n555), .Z(n583) );
  XNOR2_X1 U343 ( .A(n384), .B(n383), .ZN(n497) );
  XNOR2_X1 U344 ( .A(n335), .B(n334), .ZN(n555) );
  XNOR2_X1 U345 ( .A(n460), .B(n459), .ZN(n505) );
  XNOR2_X1 U346 ( .A(n484), .B(G190GAT), .ZN(n485) );
  XNOR2_X1 U347 ( .A(n487), .B(G43GAT), .ZN(n488) );
  XNOR2_X1 U348 ( .A(n486), .B(n485), .ZN(G1351GAT) );
  XNOR2_X1 U349 ( .A(n489), .B(n488), .ZN(G1330GAT) );
  XOR2_X1 U350 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n297) );
  XNOR2_X1 U351 ( .A(G1GAT), .B(G148GAT), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U353 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n299) );
  XNOR2_X1 U354 ( .A(KEYINPUT92), .B(KEYINPUT5), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U356 ( .A(n301), .B(n300), .Z(n313) );
  XOR2_X1 U357 ( .A(G155GAT), .B(KEYINPUT89), .Z(n303) );
  XNOR2_X1 U358 ( .A(G141GAT), .B(KEYINPUT88), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U360 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n305) );
  XNOR2_X1 U361 ( .A(G162GAT), .B(KEYINPUT90), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U363 ( .A(n307), .B(n306), .Z(n369) );
  XNOR2_X1 U364 ( .A(G120GAT), .B(G85GAT), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n308), .B(G57GAT), .ZN(n454) );
  XOR2_X1 U366 ( .A(G29GAT), .B(G134GAT), .Z(n319) );
  XOR2_X1 U367 ( .A(n454), .B(n319), .Z(n310) );
  NAND2_X1 U368 ( .A1(G225GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U370 ( .A(n369), .B(n311), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n313), .B(n312), .ZN(n318) );
  XOR2_X1 U372 ( .A(KEYINPUT0), .B(KEYINPUT80), .Z(n315) );
  XNOR2_X1 U373 ( .A(KEYINPUT79), .B(G127GAT), .ZN(n314) );
  XNOR2_X1 U374 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U375 ( .A(G113GAT), .B(n316), .Z(n405) );
  INV_X1 U376 ( .A(n405), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n318), .B(n317), .ZN(n420) );
  XNOR2_X1 U378 ( .A(KEYINPUT94), .B(n420), .ZN(n521) );
  XNOR2_X1 U379 ( .A(KEYINPUT38), .B(KEYINPUT105), .ZN(n460) );
  XOR2_X1 U380 ( .A(KEYINPUT71), .B(G85GAT), .Z(n321) );
  XOR2_X1 U381 ( .A(G50GAT), .B(KEYINPUT69), .Z(n358) );
  XNOR2_X1 U382 ( .A(n358), .B(n319), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n326) );
  XOR2_X1 U384 ( .A(KEYINPUT70), .B(G92GAT), .Z(n323) );
  XNOR2_X1 U385 ( .A(G99GAT), .B(G106GAT), .ZN(n322) );
  XNOR2_X1 U386 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U387 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n328) );
  XNOR2_X1 U388 ( .A(G162GAT), .B(KEYINPUT9), .ZN(n327) );
  XNOR2_X1 U389 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U390 ( .A(n330), .B(n329), .Z(n335) );
  XNOR2_X1 U391 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n331), .B(KEYINPUT7), .ZN(n433) );
  XOR2_X1 U393 ( .A(KEYINPUT72), .B(G218GAT), .Z(n333) );
  XNOR2_X1 U394 ( .A(G36GAT), .B(G190GAT), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n374) );
  XNOR2_X1 U396 ( .A(n433), .B(n374), .ZN(n334) );
  XOR2_X1 U397 ( .A(KEYINPUT77), .B(G155GAT), .Z(n337) );
  XNOR2_X1 U398 ( .A(G127GAT), .B(G183GAT), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U400 ( .A(KEYINPUT74), .B(KEYINPUT78), .Z(n339) );
  XNOR2_X1 U401 ( .A(G57GAT), .B(KEYINPUT73), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U403 ( .A(n341), .B(n340), .Z(n346) );
  XOR2_X1 U404 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n343) );
  NAND2_X1 U405 ( .A1(G231GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U407 ( .A(KEYINPUT75), .B(n344), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n355) );
  XOR2_X1 U409 ( .A(KEYINPUT76), .B(KEYINPUT15), .Z(n348) );
  XNOR2_X1 U410 ( .A(G8GAT), .B(G64GAT), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n353) );
  XOR2_X1 U412 ( .A(G71GAT), .B(KEYINPUT13), .Z(n444) );
  XOR2_X1 U413 ( .A(n444), .B(G211GAT), .Z(n351) );
  XNOR2_X1 U414 ( .A(G22GAT), .B(G15GAT), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n349), .B(G1GAT), .ZN(n429) );
  XNOR2_X1 U416 ( .A(n429), .B(G78GAT), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U418 ( .A(n353), .B(n352), .Z(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n567) );
  NOR2_X1 U420 ( .A1(n583), .A2(n567), .ZN(n426) );
  XOR2_X1 U421 ( .A(G211GAT), .B(KEYINPUT87), .Z(n357) );
  XNOR2_X1 U422 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n382) );
  XOR2_X1 U424 ( .A(G204GAT), .B(n382), .Z(n360) );
  XNOR2_X1 U425 ( .A(G218GAT), .B(n358), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n360), .B(n359), .ZN(n365) );
  XNOR2_X1 U427 ( .A(G106GAT), .B(G78GAT), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n361), .B(G148GAT), .ZN(n446) );
  XOR2_X1 U429 ( .A(n446), .B(KEYINPUT91), .Z(n363) );
  NAND2_X1 U430 ( .A1(G228GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U431 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U432 ( .A(n365), .B(n364), .Z(n371) );
  XOR2_X1 U433 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n367) );
  XNOR2_X1 U434 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n366) );
  XNOR2_X1 U435 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U437 ( .A(n371), .B(n370), .ZN(n480) );
  XOR2_X1 U438 ( .A(G169GAT), .B(G8GAT), .Z(n428) );
  XOR2_X1 U439 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n376) );
  XNOR2_X1 U440 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n295), .B(n372), .ZN(n373) );
  XOR2_X1 U442 ( .A(KEYINPUT19), .B(n373), .Z(n395) );
  XNOR2_X1 U443 ( .A(n395), .B(n374), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U445 ( .A(n428), .B(n377), .Z(n379) );
  NAND2_X1 U446 ( .A1(G226GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U447 ( .A(n379), .B(n378), .ZN(n384) );
  XOR2_X1 U448 ( .A(G64GAT), .B(G92GAT), .Z(n381) );
  XNOR2_X1 U449 ( .A(G176GAT), .B(G204GAT), .ZN(n380) );
  XNOR2_X1 U450 ( .A(n381), .B(n380), .ZN(n453) );
  XOR2_X1 U451 ( .A(n382), .B(n453), .Z(n383) );
  INV_X1 U452 ( .A(n497), .ZN(n385) );
  XNOR2_X1 U453 ( .A(KEYINPUT27), .B(n385), .ZN(n410) );
  NAND2_X1 U454 ( .A1(n410), .A2(n521), .ZN(n386) );
  XOR2_X1 U455 ( .A(KEYINPUT97), .B(n386), .Z(n528) );
  NOR2_X1 U456 ( .A1(n533), .A2(n528), .ZN(n387) );
  XNOR2_X1 U457 ( .A(KEYINPUT98), .B(n387), .ZN(n408) );
  XNOR2_X1 U458 ( .A(G176GAT), .B(G120GAT), .ZN(n388) );
  XNOR2_X1 U459 ( .A(n294), .B(n388), .ZN(n392) );
  NAND2_X1 U460 ( .A1(G227GAT), .A2(G233GAT), .ZN(n390) );
  INV_X1 U461 ( .A(KEYINPUT83), .ZN(n389) );
  INV_X1 U462 ( .A(G71GAT), .ZN(n393) );
  XNOR2_X1 U463 ( .A(n394), .B(n393), .ZN(n397) );
  XNOR2_X1 U464 ( .A(G15GAT), .B(n395), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U466 ( .A(G99GAT), .B(G190GAT), .Z(n399) );
  XNOR2_X1 U467 ( .A(G43GAT), .B(G134GAT), .ZN(n398) );
  XOR2_X1 U468 ( .A(n399), .B(n398), .Z(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n407) );
  XOR2_X1 U470 ( .A(KEYINPUT81), .B(KEYINPUT20), .Z(n403) );
  XNOR2_X1 U471 ( .A(G169GAT), .B(KEYINPUT82), .ZN(n402) );
  XNOR2_X1 U472 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U473 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U474 ( .A(n407), .B(n406), .ZN(n483) );
  NAND2_X1 U475 ( .A1(n408), .A2(n483), .ZN(n425) );
  INV_X1 U476 ( .A(n483), .ZN(n530) );
  XNOR2_X1 U477 ( .A(KEYINPUT26), .B(n409), .ZN(n569) );
  NAND2_X1 U478 ( .A1(n410), .A2(n569), .ZN(n411) );
  INV_X1 U479 ( .A(n480), .ZN(n413) );
  NOR2_X1 U480 ( .A1(n483), .A2(n497), .ZN(n412) );
  NOR2_X1 U481 ( .A1(n413), .A2(n412), .ZN(n415) );
  XOR2_X1 U482 ( .A(KEYINPUT100), .B(KEYINPUT25), .Z(n414) );
  XNOR2_X1 U483 ( .A(n415), .B(n414), .ZN(n416) );
  NOR2_X1 U484 ( .A1(n417), .A2(n416), .ZN(n419) );
  INV_X1 U485 ( .A(KEYINPUT101), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n421) );
  NOR2_X1 U487 ( .A1(n421), .A2(n420), .ZN(n423) );
  NAND2_X1 U488 ( .A1(n425), .A2(n424), .ZN(n491) );
  NAND2_X1 U489 ( .A1(n426), .A2(n491), .ZN(n427) );
  XOR2_X1 U490 ( .A(KEYINPUT37), .B(n427), .Z(n520) );
  XOR2_X1 U491 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U492 ( .A1(G229GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U494 ( .A(n432), .B(KEYINPUT29), .Z(n435) );
  XNOR2_X1 U495 ( .A(n433), .B(KEYINPUT65), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n443) );
  XOR2_X1 U497 ( .A(G197GAT), .B(G36GAT), .Z(n437) );
  XNOR2_X1 U498 ( .A(G50GAT), .B(G29GAT), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U500 ( .A(KEYINPUT64), .B(KEYINPUT30), .Z(n439) );
  XNOR2_X1 U501 ( .A(G141GAT), .B(G113GAT), .ZN(n438) );
  XNOR2_X1 U502 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U503 ( .A(n441), .B(n440), .Z(n442) );
  XNOR2_X1 U504 ( .A(n443), .B(n442), .ZN(n559) );
  XNOR2_X1 U505 ( .A(G99GAT), .B(n444), .ZN(n445) );
  XNOR2_X1 U506 ( .A(n445), .B(KEYINPUT68), .ZN(n458) );
  XOR2_X1 U507 ( .A(n446), .B(KEYINPUT32), .Z(n448) );
  NAND2_X1 U508 ( .A1(G230GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n452) );
  XOR2_X1 U510 ( .A(KEYINPUT31), .B(KEYINPUT67), .Z(n450) );
  XNOR2_X1 U511 ( .A(KEYINPUT33), .B(KEYINPUT66), .ZN(n449) );
  XNOR2_X1 U512 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U513 ( .A(n452), .B(n451), .Z(n456) );
  XNOR2_X1 U514 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n456), .B(n455), .ZN(n457) );
  INV_X1 U516 ( .A(n471), .ZN(n575) );
  NAND2_X1 U517 ( .A1(n559), .A2(n575), .ZN(n493) );
  NAND2_X1 U518 ( .A1(n521), .A2(n505), .ZN(n463) );
  XOR2_X1 U519 ( .A(KEYINPUT39), .B(KEYINPUT106), .Z(n461) );
  XNOR2_X1 U520 ( .A(n461), .B(G29GAT), .ZN(n462) );
  XNOR2_X1 U521 ( .A(n463), .B(n462), .ZN(G1328GAT) );
  INV_X1 U522 ( .A(n559), .ZN(n571) );
  XNOR2_X1 U523 ( .A(KEYINPUT41), .B(n471), .ZN(n547) );
  NOR2_X1 U524 ( .A1(n571), .A2(n547), .ZN(n464) );
  XNOR2_X1 U525 ( .A(n464), .B(KEYINPUT46), .ZN(n465) );
  NOR2_X1 U526 ( .A1(n567), .A2(n465), .ZN(n466) );
  XNOR2_X1 U527 ( .A(n466), .B(KEYINPUT113), .ZN(n467) );
  NOR2_X1 U528 ( .A1(n555), .A2(n467), .ZN(n468) );
  XNOR2_X1 U529 ( .A(n468), .B(KEYINPUT47), .ZN(n475) );
  INV_X1 U530 ( .A(n567), .ZN(n580) );
  NOR2_X1 U531 ( .A1(n583), .A2(n580), .ZN(n470) );
  NOR2_X1 U532 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U533 ( .A1(n473), .A2(n571), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n477) );
  XOR2_X1 U535 ( .A(KEYINPUT114), .B(KEYINPUT48), .Z(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(n529) );
  NOR2_X1 U537 ( .A1(n529), .A2(n497), .ZN(n478) );
  XOR2_X1 U538 ( .A(KEYINPUT54), .B(n478), .Z(n479) );
  NAND2_X1 U539 ( .A1(n570), .A2(n480), .ZN(n481) );
  XOR2_X1 U540 ( .A(KEYINPUT55), .B(n481), .Z(n482) );
  NOR2_X2 U541 ( .A1(n483), .A2(n482), .ZN(n562) );
  NAND2_X1 U542 ( .A1(n562), .A2(n555), .ZN(n486) );
  XOR2_X1 U543 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n484) );
  NAND2_X1 U544 ( .A1(n505), .A2(n530), .ZN(n489) );
  XOR2_X1 U545 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n487) );
  XOR2_X1 U546 ( .A(KEYINPUT34), .B(KEYINPUT103), .Z(n495) );
  NOR2_X1 U547 ( .A1(n555), .A2(n580), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n490), .B(KEYINPUT16), .ZN(n492) );
  NAND2_X1 U549 ( .A1(n492), .A2(n491), .ZN(n508) );
  NOR2_X1 U550 ( .A1(n493), .A2(n508), .ZN(n502) );
  NAND2_X1 U551 ( .A1(n502), .A2(n521), .ZN(n494) );
  XNOR2_X1 U552 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U553 ( .A(G1GAT), .B(n496), .ZN(G1324GAT) );
  NAND2_X1 U554 ( .A1(n502), .A2(n385), .ZN(n498) );
  XNOR2_X1 U555 ( .A(n498), .B(KEYINPUT104), .ZN(n499) );
  XNOR2_X1 U556 ( .A(G8GAT), .B(n499), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(G15GAT), .B(KEYINPUT35), .Z(n501) );
  NAND2_X1 U558 ( .A1(n502), .A2(n530), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n501), .B(n500), .ZN(G1326GAT) );
  NAND2_X1 U560 ( .A1(n502), .A2(n533), .ZN(n503) );
  XNOR2_X1 U561 ( .A(n503), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U562 ( .A1(n505), .A2(n385), .ZN(n504) );
  XNOR2_X1 U563 ( .A(G36GAT), .B(n504), .ZN(G1329GAT) );
  NAND2_X1 U564 ( .A1(n505), .A2(n533), .ZN(n506) );
  XNOR2_X1 U565 ( .A(n506), .B(KEYINPUT108), .ZN(n507) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n507), .ZN(G1331GAT) );
  XNOR2_X1 U567 ( .A(n547), .B(KEYINPUT109), .ZN(n561) );
  NAND2_X1 U568 ( .A1(n571), .A2(n561), .ZN(n519) );
  NOR2_X1 U569 ( .A1(n508), .A2(n519), .ZN(n509) );
  XNOR2_X1 U570 ( .A(n509), .B(KEYINPUT110), .ZN(n515) );
  NAND2_X1 U571 ( .A1(n521), .A2(n515), .ZN(n510) );
  XNOR2_X1 U572 ( .A(KEYINPUT42), .B(n510), .ZN(n511) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n511), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n515), .A2(n385), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n512), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U576 ( .A(G71GAT), .B(KEYINPUT111), .Z(n514) );
  NAND2_X1 U577 ( .A1(n515), .A2(n530), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U580 ( .A1(n533), .A2(n515), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U583 ( .A1(n520), .A2(n519), .ZN(n525) );
  NAND2_X1 U584 ( .A1(n525), .A2(n521), .ZN(n522) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n525), .A2(n385), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n530), .A2(n525), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U590 ( .A1(n525), .A2(n533), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n526), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n535) );
  NOR2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n545) );
  NAND2_X1 U595 ( .A1(n545), .A2(n530), .ZN(n531) );
  XOR2_X1 U596 ( .A(KEYINPUT115), .B(n531), .Z(n532) );
  NOR2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n542), .A2(n559), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U601 ( .A1(n542), .A2(n561), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n538), .Z(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n540) );
  NAND2_X1 U605 ( .A1(n542), .A2(n567), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U609 ( .A1(n542), .A2(n555), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U611 ( .A1(n545), .A2(n569), .ZN(n556) );
  NOR2_X1 U612 ( .A1(n571), .A2(n556), .ZN(n546) );
  XOR2_X1 U613 ( .A(G141GAT), .B(n546), .Z(G1344GAT) );
  NOR2_X1 U614 ( .A1(n547), .A2(n556), .ZN(n552) );
  XOR2_X1 U615 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n549) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U618 ( .A(KEYINPUT53), .B(n550), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n580), .A2(n556), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(G1346GAT) );
  INV_X1 U623 ( .A(n555), .ZN(n557) );
  NOR2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(G162GAT), .B(n558), .Z(G1347GAT) );
  NAND2_X1 U626 ( .A1(n562), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n566) );
  XOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT56), .Z(n564) );
  NAND2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  NAND2_X1 U633 ( .A1(n567), .A2(n562), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n582) );
  NOR2_X1 U636 ( .A1(n571), .A2(n582), .ZN(n573) );
  XNOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(n574), .ZN(G1352GAT) );
  NOR2_X1 U640 ( .A1(n582), .A2(n575), .ZN(n579) );
  XOR2_X1 U641 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n577) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n582), .ZN(n581) );
  XOR2_X1 U646 ( .A(G211GAT), .B(n581), .Z(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(G218GAT), .B(n586), .Z(G1355GAT) );
endmodule

