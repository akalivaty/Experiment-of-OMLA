//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n207), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n203), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT65), .B(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G107), .A2(G264), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n229));
  AND3_X1   g0029(.A1(new_n218), .A2(new_n228), .A3(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT66), .B(G50), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT77), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n214), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n206), .A2(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n253), .A2(new_n257), .B1(new_n248), .B2(new_n255), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT67), .A2(G41), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT67), .A2(G41), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n259), .A2(new_n260), .A3(G45), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n206), .A2(G274), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G1), .A3(G13), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G232), .ZN(new_n267));
  OAI22_X1  g0067(.A1(new_n261), .A2(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT76), .ZN(new_n269));
  INV_X1    g0069(.A(G226), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G1698), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(G223), .B2(G1698), .ZN(new_n272));
  AND2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G87), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n272), .A2(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n264), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n268), .A2(new_n269), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G190), .ZN(new_n281));
  OAI221_X1 g0081(.A(KEYINPUT76), .B1(new_n266), .B2(new_n267), .C1(new_n261), .C2(new_n262), .ZN(new_n282));
  AND3_X1   g0082(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(G200), .B1(new_n280), .B2(new_n282), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G159), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G58), .A2(G68), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT65), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G68), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n288), .B1(new_n292), .B2(G58), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n287), .B1(new_n293), .B2(new_n207), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT3), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n276), .ZN(new_n296));
  NAND2_X1  g0096(.A1(KEYINPUT3), .A2(G33), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n296), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n297), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n273), .A2(new_n274), .A3(G20), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT7), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT73), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT73), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT7), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n298), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n292), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n294), .B1(KEYINPUT74), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n296), .A2(new_n207), .A3(new_n297), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI211_X1 g0110(.A(KEYINPUT74), .B(new_n219), .C1(new_n310), .C2(new_n298), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT16), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n275), .A2(new_n309), .A3(new_n207), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n308), .A2(KEYINPUT7), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n315), .A3(G68), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n203), .B1(new_n219), .B2(new_n201), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G20), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n316), .A2(new_n318), .A3(KEYINPUT16), .A4(new_n287), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n251), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT75), .B1(new_n313), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT16), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n317), .A2(G20), .B1(G159), .B2(new_n286), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n219), .B1(new_n310), .B2(new_n298), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT74), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n322), .B1(new_n326), .B2(new_n311), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n319), .A2(new_n251), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT75), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AOI211_X1 g0130(.A(new_n258), .B(new_n285), .C1(new_n321), .C2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT17), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n247), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n258), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n283), .A2(new_n284), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n329), .B1(new_n327), .B2(new_n328), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n334), .B(new_n335), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(KEYINPUT77), .A3(KEYINPUT17), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT78), .B1(new_n338), .B2(KEYINPUT17), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n258), .B1(new_n321), .B2(new_n330), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT78), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n341), .A2(new_n342), .A3(new_n332), .A4(new_n335), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n333), .A2(new_n339), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n280), .A2(new_n282), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G179), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(new_n346), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT18), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT18), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n345), .A2(new_n352), .A3(new_n349), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n344), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n356));
  INV_X1    g0156(.A(G150), .ZN(new_n357));
  INV_X1    g0157(.A(new_n286), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n207), .A2(G33), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n254), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n251), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n252), .A2(G50), .A3(new_n256), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n362), .B(new_n363), .C1(G50), .C2(new_n248), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT9), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n261), .A2(new_n262), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n266), .A2(new_n270), .ZN(new_n367));
  AOI21_X1  g0167(.A(G1698), .B1(new_n296), .B2(new_n297), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G222), .ZN(new_n369));
  INV_X1    g0169(.A(G77), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n296), .A2(new_n297), .ZN(new_n371));
  INV_X1    g0171(.A(G1698), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n296), .B2(new_n297), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT68), .B(G223), .ZN(new_n375));
  OAI221_X1 g0175(.A(new_n369), .B1(new_n370), .B2(new_n371), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  AOI211_X1 g0176(.A(new_n366), .B(new_n367), .C1(new_n376), .C2(new_n279), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G190), .ZN(new_n378));
  INV_X1    g0178(.A(G200), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n365), .B(new_n378), .C1(new_n379), .C2(new_n377), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT10), .ZN(new_n381));
  INV_X1    g0181(.A(G179), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n364), .B1(new_n377), .B2(G169), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XOR2_X1   g0185(.A(new_n254), .B(KEYINPUT69), .Z(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n286), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT15), .B(G87), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n387), .B1(new_n207), .B2(new_n370), .C1(new_n360), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n251), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n252), .A2(G77), .A3(new_n256), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(G77), .B2(new_n248), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n368), .A2(G232), .B1(new_n275), .B2(G107), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n220), .B2(new_n374), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n279), .ZN(new_n397));
  INV_X1    g0197(.A(new_n266), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n366), .B1(G244), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n382), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n399), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n348), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n394), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(G200), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n397), .A2(G190), .A3(new_n399), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n390), .A2(new_n393), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n385), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n252), .A2(G68), .A3(new_n256), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT12), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n292), .A2(new_n411), .A3(new_n248), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT12), .B1(new_n249), .B2(new_n202), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n286), .A2(G50), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT70), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n415), .B(new_n416), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n292), .A2(new_n207), .B1(new_n370), .B2(new_n360), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n251), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT11), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n410), .B(new_n414), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n419), .A2(new_n420), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT71), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT71), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n421), .B2(new_n422), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT14), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n373), .A2(G232), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G97), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n371), .A2(new_n372), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n429), .B(new_n430), .C1(new_n270), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n279), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT13), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n366), .B1(G238), .B2(new_n398), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n434), .B1(new_n433), .B2(new_n435), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n428), .B(G169), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n438), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(G179), .A3(new_n436), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n436), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n428), .B1(new_n443), .B2(G169), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n427), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(G200), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n440), .A2(G190), .A3(new_n436), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n423), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT72), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n449), .B(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n355), .A2(new_n409), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT79), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT79), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n355), .A2(new_n409), .A3(new_n454), .A4(new_n451), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G41), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT5), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n264), .A2(G274), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT85), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT67), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n457), .ZN(new_n463));
  NAND2_X1  g0263(.A1(KEYINPUT67), .A2(G41), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT5), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G45), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G1), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n461), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT5), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(new_n259), .B2(new_n260), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(KEYINPUT85), .A3(new_n467), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n469), .A2(KEYINPUT86), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT86), .B1(new_n469), .B2(new_n472), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n460), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G179), .ZN(new_n476));
  INV_X1    g0276(.A(G257), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n296), .B2(new_n297), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(G1698), .B1(G33), .B2(G294), .ZN(new_n479));
  OAI211_X1 g0279(.A(G250), .B(new_n372), .C1(new_n273), .C2(new_n274), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n480), .A2(KEYINPUT95), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(KEYINPUT95), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n279), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n469), .A2(new_n472), .A3(new_n458), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(G264), .A3(new_n264), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT96), .B1(new_n476), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n484), .A2(new_n486), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT96), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(G179), .A4(new_n475), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n475), .A2(new_n486), .A3(new_n484), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G169), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n488), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT97), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT97), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n488), .A2(new_n491), .A3(new_n493), .A4(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(G20), .B1(new_n296), .B2(new_n297), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT22), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT93), .B1(new_n499), .B2(KEYINPUT92), .ZN(new_n500));
  OR2_X1    g0300(.A1(new_n499), .A2(KEYINPUT93), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n498), .A2(G87), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n207), .B(G87), .C1(new_n273), .C2(new_n274), .ZN(new_n503));
  INV_X1    g0303(.A(new_n500), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G116), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(G20), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT23), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n207), .B2(G107), .ZN(new_n509));
  INV_X1    g0309(.A(G107), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(KEYINPUT23), .A3(G20), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n502), .A2(new_n505), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT94), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT24), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT94), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n502), .A2(new_n516), .A3(new_n505), .A4(new_n512), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n515), .B1(new_n514), .B2(new_n517), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n251), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n206), .A2(G33), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n248), .A2(new_n521), .A3(new_n214), .A4(new_n250), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n522), .A2(KEYINPUT82), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(KEYINPUT82), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(new_n510), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT25), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n248), .B2(G107), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n249), .A2(KEYINPUT25), .A3(new_n510), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n520), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n495), .A2(new_n497), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT98), .ZN(new_n533));
  INV_X1    g0333(.A(new_n531), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT86), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n465), .A2(new_n461), .A3(new_n468), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT85), .B1(new_n471), .B2(new_n467), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n469), .A2(KEYINPUT86), .A3(new_n472), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n459), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n379), .B1(new_n487), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n475), .A2(new_n281), .A3(new_n486), .A4(new_n484), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n534), .A2(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n532), .A2(new_n533), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n533), .B1(new_n532), .B2(new_n544), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT87), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n538), .A2(new_n539), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G283), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n550), .B(KEYINPUT84), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(G250), .B2(new_n373), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT4), .ZN(new_n553));
  INV_X1    g0353(.A(G244), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n431), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n368), .A2(KEYINPUT4), .A3(G244), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n549), .A2(new_n460), .B1(new_n279), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n485), .A2(G257), .A3(new_n264), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n548), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(new_n279), .ZN(new_n561));
  AND4_X1   g0361(.A1(new_n548), .A2(new_n475), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n348), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n475), .A2(new_n559), .A3(new_n561), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(G179), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n305), .A2(G107), .B1(G77), .B2(new_n286), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  OR2_X1    g0368(.A1(KEYINPUT80), .A2(KEYINPUT6), .ZN(new_n569));
  NAND2_X1  g0369(.A1(KEYINPUT80), .A2(KEYINPUT6), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(G97), .A3(new_n510), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT81), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n569), .A2(new_n570), .ZN(new_n574));
  XNOR2_X1  g0374(.A(G97), .B(G107), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n572), .A2(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n571), .A2(KEYINPUT81), .A3(G97), .A4(new_n510), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n207), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n251), .B1(new_n568), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n249), .A2(G97), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n525), .B2(G97), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n563), .A2(new_n566), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n564), .A2(G200), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n250), .A2(new_n214), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n574), .A2(new_n575), .ZN(new_n587));
  INV_X1    g0387(.A(G97), .ZN(new_n588));
  AOI211_X1 g0388(.A(new_n588), .B(G107), .C1(new_n569), .C2(new_n570), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n587), .B1(new_n589), .B2(KEYINPUT81), .ZN(new_n590));
  INV_X1    g0390(.A(new_n577), .ZN(new_n591));
  OAI21_X1  g0391(.A(G20), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n586), .B1(new_n592), .B2(new_n567), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT83), .B1(new_n593), .B2(new_n581), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT83), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n579), .A2(new_n595), .A3(new_n582), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n585), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n564), .A2(KEYINPUT87), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n558), .A2(new_n548), .A3(new_n559), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n599), .A3(G190), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n368), .A2(G238), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n371), .A2(G244), .A3(G1698), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n603), .A3(new_n506), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n279), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT88), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n606), .A2(new_n607), .A3(new_n264), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n607), .B1(new_n606), .B2(new_n264), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(G250), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n206), .B2(G45), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT89), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n612), .A2(new_n264), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n612), .B2(new_n264), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n605), .A2(new_n610), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G200), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n605), .A2(G190), .A3(new_n610), .A4(new_n616), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n498), .A2(G68), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT19), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n207), .B1(new_n430), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n277), .A2(new_n588), .A3(new_n510), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n621), .B1(new_n360), .B2(new_n588), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n620), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n251), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n523), .A2(G87), .A3(new_n524), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n388), .A2(new_n249), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n618), .A2(new_n619), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n605), .A2(G179), .A3(new_n610), .A4(new_n616), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n373), .A2(G244), .B1(G33), .B2(G116), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n264), .B1(new_n634), .B2(new_n602), .ZN(new_n635));
  OAI22_X1  g0435(.A1(new_n608), .A2(new_n609), .B1(new_n614), .B2(new_n615), .ZN(new_n636));
  OAI21_X1  g0436(.A(G169), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n633), .A2(new_n637), .A3(KEYINPUT90), .ZN(new_n638));
  INV_X1    g0438(.A(new_n388), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n523), .A2(new_n639), .A3(new_n524), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n627), .A2(new_n640), .A3(new_n629), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n633), .A2(new_n637), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT90), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n632), .B1(new_n638), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n584), .A2(new_n601), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n485), .A2(G270), .A3(new_n264), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n478), .A2(new_n372), .B1(new_n275), .B2(G303), .ZN(new_n649));
  INV_X1    g0449(.A(G264), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n649), .B1(new_n650), .B2(new_n374), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n279), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n475), .A2(new_n648), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT20), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n207), .B1(new_n588), .B2(G33), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n551), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n251), .B1(new_n207), .B2(G116), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n657), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n659), .B(KEYINPUT20), .C1(new_n551), .C2(new_n655), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  MUX2_X1   g0461(.A(new_n248), .B(new_n522), .S(G116), .Z(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n653), .A2(new_n664), .A3(new_n382), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n348), .B1(new_n661), .B2(new_n662), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n653), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT21), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT21), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n653), .A2(new_n669), .A3(new_n666), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n665), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT91), .ZN(new_n672));
  INV_X1    g0472(.A(new_n653), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G190), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n653), .A2(G200), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n664), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n671), .A2(new_n672), .A3(new_n676), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n674), .A2(new_n664), .A3(new_n675), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n673), .A2(G179), .A3(new_n663), .ZN(new_n679));
  INV_X1    g0479(.A(new_n670), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n669), .B1(new_n653), .B2(new_n666), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT91), .B1(new_n678), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n647), .B1(new_n677), .B2(new_n683), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n456), .A2(new_n547), .A3(new_n684), .ZN(G372));
  NAND2_X1  g0485(.A1(new_n594), .A2(new_n596), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n643), .A2(new_n641), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n631), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n563), .A2(new_n566), .A3(new_n686), .A4(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n598), .A2(new_n599), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n565), .B1(new_n692), .B2(new_n348), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(KEYINPUT26), .A3(new_n583), .A4(new_n646), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n494), .A2(new_n531), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n671), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n631), .A2(new_n687), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n534), .B2(new_n543), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n697), .A2(new_n584), .A3(new_n601), .A4(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n695), .A2(new_n700), .A3(new_n687), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n456), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n383), .A2(new_n384), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n342), .B1(new_n331), .B2(new_n332), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n338), .A2(KEYINPUT78), .A3(KEYINPUT17), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n338), .A2(KEYINPUT77), .A3(KEYINPUT17), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT77), .B1(new_n338), .B2(KEYINPUT17), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n704), .A2(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n448), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n445), .B1(new_n709), .B2(new_n403), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n354), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n711), .A2(KEYINPUT99), .ZN(new_n712));
  INV_X1    g0512(.A(new_n381), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n711), .B2(KEYINPUT99), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n703), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n702), .A2(new_n715), .ZN(G369));
  NAND3_X1  g0516(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n717), .A2(KEYINPUT27), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(KEYINPUT27), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G213), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(G343), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n547), .B1(new_n534), .B2(new_n723), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n532), .A2(new_n723), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n683), .A2(new_n677), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n664), .B2(new_n723), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n682), .A2(new_n663), .A3(new_n722), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT100), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT100), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n728), .A2(new_n732), .A3(new_n729), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(G330), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n726), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n671), .A2(new_n722), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n545), .B2(new_n546), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n494), .A2(new_n531), .A3(new_n723), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT101), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n738), .A2(KEYINPUT101), .A3(new_n739), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n736), .A2(new_n744), .ZN(G399));
  INV_X1    g0545(.A(new_n210), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n259), .A2(new_n260), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n623), .A2(G116), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(G1), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(new_n216), .B2(new_n750), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT28), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n693), .A2(new_n690), .A3(new_n583), .A4(new_n646), .ZN(new_n755));
  INV_X1    g0555(.A(new_n687), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n689), .B2(KEYINPUT26), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n532), .A2(new_n671), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n693), .A2(new_n583), .B1(new_n597), .B2(new_n600), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n699), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n755), .B(new_n757), .C1(new_n758), .C2(new_n760), .ZN(new_n761));
  AND3_X1   g0561(.A1(new_n761), .A2(KEYINPUT102), .A3(new_n723), .ZN(new_n762));
  AOI21_X1  g0562(.A(KEYINPUT102), .B1(new_n761), .B2(new_n723), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT29), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n701), .A2(new_n723), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT29), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n684), .B(new_n723), .C1(new_n545), .C2(new_n546), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n617), .A2(new_n382), .ZN(new_n770));
  AND4_X1   g0570(.A1(new_n492), .A2(new_n770), .A3(new_n653), .A4(new_n564), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n653), .A2(new_n487), .A3(new_n633), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n772), .A2(new_n598), .A3(new_n599), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT30), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n772), .A2(KEYINPUT30), .A3(new_n598), .A4(new_n599), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n723), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT31), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n769), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G330), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n768), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n754), .B1(new_n783), .B2(G1), .ZN(G364));
  NAND2_X1  g0584(.A1(new_n207), .A2(G13), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT103), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G45), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G1), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n749), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n734), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n731), .A2(new_n733), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n791), .B1(G330), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G13), .A2(G33), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n207), .A2(G179), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G190), .A2(G200), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT104), .B(G159), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT32), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n207), .A2(new_n382), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n801), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n808), .A2(G190), .A3(new_n379), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n371), .B1(new_n809), .B2(new_n370), .C1(new_n201), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n808), .A2(G200), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n281), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G50), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n281), .A2(G179), .A3(G200), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n207), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n814), .A2(new_n815), .B1(new_n588), .B2(new_n817), .ZN(new_n818));
  OR3_X1    g0618(.A1(new_n807), .A2(new_n811), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n800), .A2(new_n281), .A3(G200), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n510), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n800), .A2(G190), .A3(G200), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n812), .A2(G190), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n822), .B1(new_n277), .B2(new_n823), .C1(new_n825), .C2(new_n202), .ZN(new_n826));
  INV_X1    g0626(.A(new_n823), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n813), .A2(G326), .B1(new_n827), .B2(G303), .ZN(new_n828));
  INV_X1    g0628(.A(G283), .ZN(new_n829));
  INV_X1    g0629(.A(G294), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n828), .B1(new_n829), .B2(new_n820), .C1(new_n830), .C2(new_n817), .ZN(new_n831));
  INV_X1    g0631(.A(new_n810), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n832), .A2(G322), .B1(new_n803), .B2(G329), .ZN(new_n833));
  XNOR2_X1  g0633(.A(KEYINPUT33), .B(G317), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n834), .A2(KEYINPUT105), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(KEYINPUT105), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n835), .A2(new_n824), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n809), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n371), .B1(new_n838), .B2(G311), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n833), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n819), .A2(new_n826), .B1(new_n831), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n214), .B1(G20), .B2(new_n348), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n797), .A2(new_n842), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n746), .A2(new_n371), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(G45), .B2(new_n216), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(new_n242), .B2(G45), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n746), .A2(new_n275), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(G355), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(G116), .B2(new_n210), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n844), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n843), .A2(new_n851), .A3(new_n789), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n794), .B1(new_n799), .B2(new_n852), .ZN(G396));
  NOR2_X1   g0653(.A1(new_n842), .A2(new_n795), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n790), .B1(new_n370), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n842), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n832), .A2(G143), .B1(new_n838), .B2(new_n805), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n857), .B1(new_n814), .B2(new_n858), .C1(new_n357), .C2(new_n825), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT34), .ZN(new_n860));
  INV_X1    g0660(.A(G132), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n371), .B1(new_n802), .B2(new_n861), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n817), .A2(new_n201), .B1(new_n823), .B2(new_n815), .ZN(new_n863));
  INV_X1    g0663(.A(new_n820), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n862), .B(new_n863), .C1(G68), .C2(new_n864), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n824), .A2(G283), .B1(new_n838), .B2(G116), .ZN(new_n866));
  INV_X1    g0666(.A(G303), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n866), .B1(new_n867), .B2(new_n814), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT106), .Z(new_n869));
  OAI22_X1  g0669(.A1(new_n817), .A2(new_n588), .B1(new_n810), .B2(new_n830), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT107), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n823), .A2(new_n510), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n820), .A2(new_n277), .ZN(new_n873));
  INV_X1    g0673(.A(G311), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n275), .B1(new_n802), .B2(new_n874), .ZN(new_n875));
  NOR4_X1   g0675(.A1(new_n871), .A2(new_n872), .A3(new_n873), .A4(new_n875), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n860), .A2(new_n865), .B1(new_n869), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n403), .A2(new_n722), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n394), .A2(new_n722), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n406), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n878), .B1(new_n403), .B2(new_n880), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n855), .B1(new_n856), .B2(new_n877), .C1(new_n881), .C2(new_n796), .ZN(new_n882));
  INV_X1    g0682(.A(new_n881), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n765), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n407), .A2(new_n723), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n701), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n789), .B1(new_n781), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n781), .A2(new_n888), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n882), .B1(new_n890), .B2(new_n891), .ZN(G384));
  NOR2_X1   g0692(.A1(new_n590), .A2(new_n591), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n894), .A2(KEYINPUT35), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(KEYINPUT35), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n895), .A2(G116), .A3(new_n215), .A4(new_n896), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT36), .Z(new_n898));
  OAI211_X1 g0698(.A(new_n217), .B(G77), .C1(new_n201), .C2(new_n219), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n815), .A2(G68), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n206), .B(G13), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n354), .ZN(new_n903));
  INV_X1    g0703(.A(new_n720), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT110), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n445), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n427), .B(KEYINPUT110), .C1(new_n442), .C2(new_n444), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n424), .A2(new_n426), .A3(new_n722), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n448), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n908), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n442), .A2(new_n444), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n427), .B(new_n722), .C1(new_n913), .C2(new_n709), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT109), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n878), .B(KEYINPUT108), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n916), .B1(new_n887), .B2(new_n918), .ZN(new_n919));
  AOI211_X1 g0719(.A(KEYINPUT109), .B(new_n917), .C1(new_n701), .C2(new_n886), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT38), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT16), .B1(new_n323), .B2(new_n316), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n334), .B1(new_n320), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n904), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n708), .B2(new_n903), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n345), .A2(new_n904), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT37), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n350), .A2(new_n927), .A3(new_n928), .A4(new_n338), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n924), .B1(new_n349), .B2(new_n904), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n338), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT37), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n922), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n925), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n344), .B2(new_n354), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(KEYINPUT38), .A3(new_n933), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n906), .B1(new_n921), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT111), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n541), .A2(new_n542), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n688), .B1(new_n943), .B2(new_n531), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n671), .B2(new_n696), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n756), .B1(new_n945), .B2(new_n759), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n885), .B1(new_n946), .B2(new_n695), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT109), .B1(new_n947), .B2(new_n917), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n887), .A2(new_n916), .A3(new_n918), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(new_n939), .A3(new_n915), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT111), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n952), .A3(new_n906), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n942), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n927), .B1(new_n708), .B2(new_n903), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n927), .A2(new_n350), .A3(new_n338), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(new_n928), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n922), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT39), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n958), .A2(new_n959), .A3(new_n938), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n959), .B1(new_n935), .B2(new_n938), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT112), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n926), .A2(new_n922), .A3(new_n934), .ZN(new_n963));
  AOI21_X1  g0763(.A(KEYINPUT38), .B1(new_n937), .B2(new_n933), .ZN(new_n964));
  OAI21_X1  g0764(.A(KEYINPUT39), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n958), .A2(new_n938), .A3(new_n959), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT112), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n962), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n908), .A2(new_n909), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(new_n722), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n954), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n764), .A2(new_n456), .A3(new_n767), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n715), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n973), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n915), .A2(new_n881), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n769), .B2(new_n779), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n963), .B2(new_n964), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT40), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(new_n958), .B2(new_n938), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n979), .A2(new_n980), .B1(new_n981), .B2(new_n978), .ZN(new_n982));
  AND3_X1   g0782(.A1(new_n982), .A2(new_n456), .A3(new_n780), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n982), .B1(new_n456), .B2(new_n780), .ZN(new_n984));
  INV_X1    g0784(.A(G330), .ZN(new_n985));
  OR3_X1    g0785(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n976), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n206), .B2(new_n786), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n976), .A2(new_n986), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n902), .B1(new_n988), .B2(new_n989), .ZN(G367));
  NOR2_X1   g0790(.A1(new_n630), .A2(new_n723), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n756), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n698), .B2(new_n991), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n994));
  AND3_X1   g0794(.A1(new_n693), .A2(new_n686), .A3(new_n722), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n686), .A2(new_n722), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n995), .B1(new_n759), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n547), .A2(new_n737), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n584), .B1(new_n997), .B2(new_n532), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n723), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n994), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT113), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1005), .B(new_n1007), .Z(new_n1008));
  NOR2_X1   g0808(.A1(new_n736), .A2(new_n997), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n749), .B(KEYINPUT41), .Z(new_n1012));
  AOI21_X1  g0812(.A(new_n997), .B1(new_n742), .B2(new_n743), .ZN(new_n1013));
  XOR2_X1   g0813(.A(KEYINPUT114), .B(KEYINPUT45), .Z(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n744), .A2(new_n998), .A3(new_n1014), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n742), .A2(new_n743), .A3(new_n997), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT44), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n735), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n724), .B(new_n725), .C1(new_n671), .C2(new_n722), .ZN(new_n1021));
  AND3_X1   g0821(.A1(new_n1021), .A2(new_n734), .A3(new_n738), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n734), .B1(new_n1021), .B2(new_n738), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1024), .A2(new_n782), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT44), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1018), .B(new_n1026), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1027), .A2(new_n736), .A3(new_n1016), .A4(new_n1015), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1020), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1012), .B1(new_n1029), .B2(new_n783), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1010), .B(new_n1011), .C1(new_n1030), .C2(new_n788), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n845), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n844), .B1(new_n210), .B2(new_n388), .C1(new_n1032), .C2(new_n237), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT115), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n790), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n1034), .B2(new_n1033), .ZN(new_n1036));
  INV_X1    g0836(.A(G317), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n275), .B1(new_n802), .B2(new_n1037), .C1(new_n810), .C2(new_n867), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n825), .A2(new_n830), .B1(new_n814), .B2(new_n874), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(G97), .C2(new_n864), .ZN(new_n1040));
  INV_X1    g0840(.A(G116), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT117), .B1(new_n823), .B2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT46), .Z(new_n1043));
  OAI22_X1  g0843(.A1(new_n817), .A2(new_n510), .B1(new_n809), .B2(new_n829), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT116), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1040), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n810), .A2(new_n357), .B1(new_n802), .B2(new_n858), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n275), .B(new_n1047), .C1(G50), .C2(new_n838), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n824), .A2(new_n805), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n817), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1050), .A2(G68), .B1(new_n827), .B2(G58), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n813), .A2(G143), .B1(new_n864), .B2(G77), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1046), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT47), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1036), .B1(new_n1055), .B2(new_n842), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n993), .B2(new_n798), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1031), .A2(new_n1057), .ZN(G387));
  OAI22_X1  g0858(.A1(new_n810), .A2(new_n815), .B1(new_n809), .B2(new_n202), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n275), .B(new_n1059), .C1(G150), .C2(new_n803), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n824), .A2(new_n255), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n639), .A2(new_n1050), .B1(new_n813), .B2(G159), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n827), .A2(G77), .B1(new_n864), .B2(G97), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n371), .B1(new_n803), .B2(G326), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n817), .A2(new_n829), .B1(new_n823), .B2(new_n830), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n832), .A2(G317), .B1(new_n838), .B2(G303), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n813), .A2(G322), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(new_n874), .C2(new_n825), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n1070), .B2(new_n1069), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT49), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1065), .B1(new_n1041), .B2(new_n820), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1064), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n842), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n751), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n848), .A2(new_n1078), .B1(new_n510), .B2(new_n746), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n386), .A2(new_n815), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT50), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n751), .B(new_n466), .C1(new_n202), .C2(new_n370), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT118), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n845), .B1(new_n234), .B2(new_n466), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1079), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n790), .B1(new_n1086), .B2(new_n844), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1077), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n726), .B2(new_n797), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1024), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n788), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1025), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n749), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1090), .A2(new_n783), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(G393));
  NAND3_X1  g0895(.A1(new_n1020), .A2(new_n1028), .A3(new_n788), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G150), .A2(new_n813), .B1(new_n832), .B2(G159), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT51), .Z(new_n1098));
  NOR2_X1   g0898(.A1(new_n823), .A2(new_n219), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n817), .A2(new_n370), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(G50), .C2(new_n824), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n386), .A2(new_n838), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n275), .B(new_n873), .C1(G143), .C2(new_n803), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1098), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n814), .A2(new_n1037), .B1(new_n874), .B2(new_n810), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT52), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n275), .B1(new_n809), .B2(new_n830), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G322), .B2(new_n803), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n821), .B1(G116), .B2(new_n1050), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n824), .A2(G303), .B1(new_n827), .B2(G283), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n856), .B1(new_n1104), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n845), .A2(new_n245), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n797), .B(new_n842), .C1(new_n746), .C2(G97), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n790), .B(new_n1112), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT119), .Z(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n998), .B2(new_n798), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1096), .A2(new_n1117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1029), .A2(new_n749), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1020), .A2(new_n1028), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n1092), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1118), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(G390));
  INV_X1    g0923(.A(new_n971), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n921), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n962), .A2(new_n968), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n971), .B1(new_n958), .B2(new_n938), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n761), .A2(new_n723), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT102), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n761), .A2(KEYINPUT102), .A3(new_n723), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n878), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n880), .A2(new_n403), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n915), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1127), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1126), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n985), .B1(new_n769), .B2(new_n779), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1139), .A2(new_n881), .A3(new_n915), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1126), .A2(new_n1137), .A3(new_n1140), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n456), .A2(new_n1139), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n974), .A2(new_n715), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n915), .B1(new_n1139), .B2(new_n881), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1135), .A2(new_n1149), .A3(new_n1140), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n950), .B1(new_n1141), .B2(new_n1148), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1147), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n750), .B1(new_n1144), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1146), .B1(new_n1151), .B2(new_n1150), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1142), .A2(new_n1143), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT121), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1142), .A2(new_n788), .A3(new_n1143), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT54), .B(G143), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n810), .A2(new_n861), .B1(new_n809), .B2(new_n1160), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n275), .B(new_n1161), .C1(G125), .C2(new_n803), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n823), .A2(new_n357), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT53), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n813), .A2(G128), .B1(new_n864), .B2(G50), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G159), .A2(new_n1050), .B1(new_n824), .B2(G137), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1162), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n824), .A2(G107), .B1(new_n838), .B2(G97), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n829), .B2(new_n814), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT120), .Z(new_n1170));
  OAI221_X1 g0970(.A(new_n275), .B1(new_n802), .B2(new_n830), .C1(new_n810), .C2(new_n1041), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n202), .A2(new_n820), .B1(new_n823), .B2(new_n277), .ZN(new_n1172));
  OR3_X1    g0972(.A1(new_n1171), .A2(new_n1100), .A3(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1167), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n842), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n790), .B1(new_n254), .B2(new_n854), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n969), .C2(new_n796), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1158), .B1(new_n1159), .B2(new_n1177), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1159), .A2(new_n1158), .A3(new_n1177), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1157), .B1(new_n1178), .B2(new_n1179), .ZN(G378));
  AOI21_X1  g0980(.A(new_n1136), .B1(new_n948), .B2(new_n949), .ZN(new_n1181));
  AOI211_X1 g0981(.A(KEYINPUT111), .B(new_n905), .C1(new_n1181), .C2(new_n939), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n952), .B1(new_n951), .B2(new_n906), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1124), .B1(new_n962), .B2(new_n968), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n979), .A2(new_n980), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n981), .A2(new_n978), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n364), .A2(new_n904), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n385), .B(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  AND4_X1   g0991(.A1(G330), .A2(new_n1186), .A3(new_n1187), .A4(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n982), .B2(G330), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1184), .A2(new_n1185), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1186), .A2(G330), .A3(new_n1187), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1191), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n982), .A2(G330), .A3(new_n1191), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n954), .A2(new_n972), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT123), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1194), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n973), .B(KEYINPUT123), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n788), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n790), .B1(new_n815), .B2(new_n854), .ZN(new_n1204));
  AOI211_X1 g1004(.A(G33), .B(G41), .C1(new_n803), .C2(G124), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n820), .B2(new_n804), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n813), .A2(G125), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n825), .B2(new_n861), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n832), .A2(G128), .B1(new_n838), .B2(G137), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n823), .B2(new_n1160), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1208), .B(new_n1210), .C1(G150), .C2(new_n1050), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1206), .B1(new_n1212), .B2(KEYINPUT59), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(KEYINPUT59), .B2(new_n1212), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n825), .A2(new_n588), .B1(new_n820), .B2(new_n201), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G116), .B2(new_n813), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n371), .B(new_n748), .C1(G283), .C2(new_n803), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n832), .A2(G107), .B1(new_n838), .B2(new_n639), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1050), .A2(G68), .B1(new_n827), .B2(G77), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT58), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n815), .B1(G33), .B2(G41), .C1(new_n748), .C2(new_n371), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1224));
  AND4_X1   g1024(.A1(new_n1214), .A2(new_n1222), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1204), .B1(new_n856), .B2(new_n1225), .C1(new_n1191), .C2(new_n796), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT122), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1203), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT57), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1126), .A2(new_n1137), .A3(new_n1140), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1140), .B1(new_n1126), .B2(new_n1137), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1146), .B1(new_n1233), .B2(new_n1152), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1229), .B1(new_n1230), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1156), .A2(new_n1147), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1229), .B1(new_n1194), .B2(new_n1199), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n750), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1228), .B1(new_n1235), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(G375));
  INV_X1    g1040(.A(new_n1012), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1146), .A2(new_n1151), .A3(new_n1150), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1153), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1136), .A2(new_n795), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n825), .A2(new_n1041), .B1(new_n588), .B2(new_n823), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G294), .B2(new_n813), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n864), .A2(G77), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1050), .A2(new_n639), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n810), .A2(new_n829), .B1(new_n809), .B2(new_n510), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n371), .B(new_n1249), .C1(G303), .C2(new_n803), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n1250), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n810), .A2(new_n858), .B1(new_n809), .B2(new_n357), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n275), .B(new_n1252), .C1(G128), .C2(new_n803), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n827), .A2(G159), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1160), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G132), .A2(new_n813), .B1(new_n824), .B2(new_n1255), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1050), .A2(G50), .B1(new_n864), .B2(G58), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1253), .A2(new_n1254), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n856), .B1(new_n1251), .B2(new_n1258), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n790), .B(new_n1259), .C1(new_n202), .C2(new_n854), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1152), .A2(new_n788), .B1(new_n1244), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1243), .A2(new_n1261), .ZN(G381));
  AND3_X1   g1062(.A1(new_n1031), .A2(new_n1057), .A3(new_n1122), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1159), .A2(new_n1177), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1263), .A2(new_n1239), .A3(new_n1265), .A4(new_n1266), .ZN(G407));
  NAND3_X1  g1067(.A1(new_n1239), .A2(new_n721), .A3(new_n1265), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(G407), .A2(G213), .A3(new_n1268), .ZN(G409));
  XNOR2_X1  g1069(.A(G393), .B(G396), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1122), .B1(new_n1031), .B2(new_n1057), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1271), .B1(new_n1263), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G387), .A2(G390), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1031), .A2(new_n1122), .A3(new_n1057), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1270), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1146), .A2(new_n1150), .A3(KEYINPUT60), .A4(new_n1151), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(KEYINPUT125), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1242), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n749), .B(new_n1153), .C1(new_n1281), .C2(KEYINPUT60), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1261), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(G384), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G384), .B(new_n1261), .C1(new_n1280), .C2(new_n1282), .ZN(new_n1286));
  INV_X1    g1086(.A(G213), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1287), .A2(G343), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(G2897), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1285), .A2(new_n1286), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1289), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1194), .A2(new_n1199), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT124), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1194), .A2(new_n1199), .A3(KEYINPUT124), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1295), .A2(new_n788), .A3(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1236), .A2(new_n1241), .A3(new_n1202), .A4(new_n1201), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n1227), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n1239), .A2(G378), .B1(new_n1265), .B2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1292), .B1(new_n1300), .B2(new_n1288), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1235), .A2(new_n1238), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1228), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(G378), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1299), .A2(new_n1265), .ZN(new_n1306));
  AOI211_X1 g1106(.A(new_n1302), .B(new_n1288), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT62), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1278), .B(new_n1301), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1288), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NOR3_X1   g1112(.A1(new_n1312), .A2(KEYINPUT62), .A3(new_n1302), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1277), .B1(new_n1309), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1312), .B2(new_n1302), .ZN(new_n1316));
  AOI21_X1  g1116(.A(KEYINPUT61), .B1(new_n1312), .B2(new_n1292), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1307), .A2(KEYINPUT63), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1316), .A2(new_n1317), .A3(new_n1318), .A4(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1314), .A2(new_n1320), .ZN(G405));
  INV_X1    g1121(.A(KEYINPUT126), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1265), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1322), .B1(new_n1239), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1305), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1239), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1285), .B(new_n1286), .C1(new_n1325), .C2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT127), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1319), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1326), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1330), .A2(new_n1302), .A3(new_n1305), .A4(new_n1324), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1277), .A2(KEYINPUT127), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1327), .A2(new_n1329), .A3(new_n1331), .A4(new_n1332), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1327), .A2(new_n1331), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1333), .B1(new_n1334), .B2(new_n1332), .ZN(G402));
endmodule


