

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777;

  NAND2_X1 U372 ( .A1(n353), .A2(n365), .ZN(n732) );
  NAND2_X2 U373 ( .A1(n450), .A2(n452), .ZN(n397) );
  AND2_X2 U374 ( .A1(n440), .A2(n542), .ZN(n456) );
  XNOR2_X2 U375 ( .A(n554), .B(n553), .ZN(n630) );
  INV_X1 U376 ( .A(n584), .ZN(n349) );
  NAND2_X1 U377 ( .A1(n412), .A2(n410), .ZN(n773) );
  AND2_X1 U378 ( .A1(n414), .A2(n413), .ZN(n412) );
  NOR2_X1 U379 ( .A1(n582), .A2(n707), .ZN(n369) );
  INV_X1 U380 ( .A(n350), .ZN(n582) );
  NAND2_X1 U381 ( .A1(n703), .A2(n702), .ZN(n592) );
  XNOR2_X2 U382 ( .A(n630), .B(KEYINPUT1), .ZN(n703) );
  OR2_X1 U383 ( .A1(n594), .A2(KEYINPUT44), .ZN(n595) );
  AND2_X1 U384 ( .A1(n396), .A2(n395), .ZN(n394) );
  NAND2_X1 U385 ( .A1(n433), .A2(n431), .ZN(n772) );
  NAND2_X1 U386 ( .A1(n411), .A2(n360), .ZN(n410) );
  AND2_X1 U387 ( .A1(n430), .A2(n429), .ZN(n433) );
  XNOR2_X1 U388 ( .A(n369), .B(KEYINPUT31), .ZN(n682) );
  XNOR2_X1 U389 ( .A(n476), .B(KEYINPUT33), .ZN(n718) );
  XNOR2_X1 U390 ( .A(n583), .B(n477), .ZN(n616) );
  XNOR2_X1 U391 ( .A(n583), .B(KEYINPUT101), .ZN(n628) );
  XNOR2_X1 U392 ( .A(n472), .B(n470), .ZN(n590) );
  XNOR2_X1 U393 ( .A(n729), .B(n728), .ZN(n460) );
  XNOR2_X1 U394 ( .A(n561), .B(n372), .ZN(n729) );
  XNOR2_X1 U395 ( .A(n483), .B(n505), .ZN(n374) );
  XNOR2_X1 U396 ( .A(n536), .B(KEYINPUT4), .ZN(n761) );
  XNOR2_X1 U397 ( .A(n484), .B(n504), .ZN(n483) );
  XNOR2_X1 U398 ( .A(n459), .B(G128), .ZN(n536) );
  XNOR2_X1 U399 ( .A(n527), .B(KEYINPUT67), .ZN(n551) );
  XNOR2_X1 U400 ( .A(G146), .B(G125), .ZN(n523) );
  BUF_X1 U401 ( .A(G104), .Z(n458) );
  XNOR2_X1 U402 ( .A(G137), .B(G140), .ZN(n563) );
  XNOR2_X2 U403 ( .A(n428), .B(n351), .ZN(n350) );
  XNOR2_X1 U404 ( .A(KEYINPUT0), .B(KEYINPUT83), .ZN(n351) );
  AND2_X1 U405 ( .A1(n722), .A2(n403), .ZN(n723) );
  XNOR2_X1 U406 ( .A(n516), .B(KEYINPUT19), .ZN(n492) );
  BUF_X1 U407 ( .A(n740), .Z(n352) );
  XNOR2_X1 U408 ( .A(n374), .B(n480), .ZN(n740) );
  AND2_X2 U409 ( .A1(n464), .A2(n438), .ZN(n353) );
  OR2_X2 U410 ( .A1(n750), .A2(KEYINPUT2), .ZN(n464) );
  XNOR2_X1 U411 ( .A(n562), .B(G472), .ZN(n583) );
  NOR2_X1 U412 ( .A1(n590), .A2(n591), .ZN(n625) );
  XNOR2_X1 U413 ( .A(KEYINPUT10), .B(n523), .ZN(n757) );
  XNOR2_X1 U414 ( .A(n655), .B(n406), .ZN(n689) );
  INV_X1 U415 ( .A(KEYINPUT38), .ZN(n406) );
  AND2_X1 U416 ( .A1(n453), .A2(n455), .ZN(n452) );
  INV_X1 U417 ( .A(n628), .ZN(n455) );
  XNOR2_X1 U418 ( .A(n561), .B(n375), .ZN(n660) );
  XNOR2_X1 U419 ( .A(n556), .B(n479), .ZN(n478) );
  XNOR2_X1 U420 ( .A(n546), .B(G146), .ZN(n561) );
  INV_X1 U421 ( .A(KEYINPUT64), .ZN(n488) );
  NOR2_X1 U422 ( .A1(n592), .A2(n616), .ZN(n476) );
  XNOR2_X1 U423 ( .A(n378), .B(n377), .ZN(n577) );
  INV_X1 U424 ( .A(KEYINPUT74), .ZN(n377) );
  NAND2_X1 U425 ( .A1(n616), .A2(n379), .ZN(n378) );
  AND2_X1 U426 ( .A1(n703), .A2(n349), .ZN(n379) );
  INV_X1 U427 ( .A(KEYINPUT82), .ZN(n496) );
  XNOR2_X1 U428 ( .A(n467), .B(KEYINPUT95), .ZN(n466) );
  INV_X1 U429 ( .A(KEYINPUT11), .ZN(n467) );
  XNOR2_X1 U430 ( .A(G140), .B(KEYINPUT94), .ZN(n465) );
  NOR2_X1 U431 ( .A1(G953), .A2(G237), .ZN(n557) );
  NOR2_X1 U432 ( .A1(n649), .A2(n391), .ZN(n390) );
  NOR2_X1 U433 ( .A1(n382), .A2(n770), .ZN(n399) );
  XNOR2_X1 U434 ( .A(n481), .B(G107), .ZN(n539) );
  INV_X1 U435 ( .A(G116), .ZN(n481) );
  XNOR2_X1 U436 ( .A(n551), .B(n550), .ZN(n556) );
  INV_X1 U437 ( .A(G134), .ZN(n550) );
  XNOR2_X1 U438 ( .A(n761), .B(G101), .ZN(n546) );
  AND2_X1 U439 ( .A1(n475), .A2(KEYINPUT35), .ZN(n423) );
  XNOR2_X1 U440 ( .A(KEYINPUT73), .B(KEYINPUT32), .ZN(n485) );
  XNOR2_X1 U441 ( .A(n552), .B(G469), .ZN(n553) );
  NOR2_X1 U442 ( .A1(n729), .A2(G902), .ZN(n554) );
  XNOR2_X1 U443 ( .A(n398), .B(KEYINPUT22), .ZN(n575) );
  XNOR2_X1 U444 ( .A(n574), .B(n573), .ZN(n584) );
  XNOR2_X1 U445 ( .A(n572), .B(KEYINPUT25), .ZN(n573) );
  XOR2_X1 U446 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n568) );
  XNOR2_X1 U447 ( .A(G128), .B(KEYINPUT77), .ZN(n567) );
  XNOR2_X1 U448 ( .A(n570), .B(KEYINPUT23), .ZN(n490) );
  XNOR2_X1 U449 ( .A(G119), .B(G110), .ZN(n564) );
  XOR2_X1 U450 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n535) );
  XNOR2_X1 U451 ( .A(n487), .B(n534), .ZN(n566) );
  XNOR2_X1 U452 ( .A(n532), .B(n531), .ZN(n731) );
  XNOR2_X1 U453 ( .A(n556), .B(n409), .ZN(n758) );
  INV_X1 U454 ( .A(n563), .ZN(n409) );
  XNOR2_X1 U455 ( .A(n547), .B(n548), .ZN(n408) );
  XOR2_X1 U456 ( .A(n458), .B(G107), .Z(n548) );
  XNOR2_X1 U457 ( .A(n756), .B(n657), .ZN(n463) );
  NOR2_X1 U458 ( .A1(n645), .A2(n612), .ZN(n613) );
  NOR2_X1 U459 ( .A1(n451), .A2(KEYINPUT65), .ZN(n435) );
  INV_X1 U460 ( .A(KEYINPUT6), .ZN(n477) );
  XNOR2_X1 U461 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U462 ( .A(n756), .B(n401), .ZN(n763) );
  XNOR2_X1 U463 ( .A(n765), .B(n402), .ZN(n401) );
  INV_X1 U464 ( .A(KEYINPUT79), .ZN(n402) );
  XNOR2_X1 U465 ( .A(KEYINPUT84), .B(G110), .ZN(n742) );
  AND2_X2 U466 ( .A1(n464), .A2(n438), .ZN(n440) );
  INV_X1 U467 ( .A(KEYINPUT78), .ZN(n439) );
  XNOR2_X1 U468 ( .A(n693), .B(n469), .ZN(n468) );
  INV_X1 U469 ( .A(KEYINPUT76), .ZN(n469) );
  INV_X1 U470 ( .A(n773), .ZN(n473) );
  INV_X1 U471 ( .A(G131), .ZN(n527) );
  AND2_X1 U472 ( .A1(n683), .A2(n678), .ZN(n693) );
  OR2_X1 U473 ( .A1(G237), .A2(G902), .ZN(n513) );
  OR2_X1 U474 ( .A1(n703), .A2(KEYINPUT102), .ZN(n454) );
  NAND2_X1 U475 ( .A1(n703), .A2(KEYINPUT102), .ZN(n453) );
  XOR2_X1 U476 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n559) );
  XNOR2_X1 U477 ( .A(n555), .B(G116), .ZN(n479) );
  XNOR2_X1 U478 ( .A(G137), .B(KEYINPUT92), .ZN(n555) );
  INV_X1 U479 ( .A(G143), .ZN(n459) );
  XNOR2_X1 U480 ( .A(n524), .B(n501), .ZN(n525) );
  XNOR2_X1 U481 ( .A(n466), .B(n465), .ZN(n524) );
  XOR2_X1 U482 ( .A(KEYINPUT17), .B(KEYINPUT86), .Z(n508) );
  XNOR2_X1 U483 ( .A(n549), .B(n506), .ZN(n510) );
  XNOR2_X1 U484 ( .A(n500), .B(n522), .ZN(n506) );
  NAND2_X1 U485 ( .A1(G234), .A2(G237), .ZN(n517) );
  XNOR2_X1 U486 ( .A(n533), .B(n471), .ZN(n470) );
  OR2_X1 U487 ( .A1(n731), .A2(G902), .ZN(n472) );
  INV_X1 U488 ( .A(G475), .ZN(n471) );
  XNOR2_X1 U489 ( .A(n389), .B(n651), .ZN(n388) );
  INV_X1 U490 ( .A(n686), .ZN(n444) );
  INV_X1 U491 ( .A(KEYINPUT45), .ZN(n601) );
  XOR2_X1 U492 ( .A(G902), .B(KEYINPUT15), .Z(n542) );
  XNOR2_X1 U493 ( .A(n629), .B(n495), .ZN(n494) );
  XNOR2_X1 U494 ( .A(KEYINPUT28), .B(KEYINPUT105), .ZN(n495) );
  NOR2_X1 U495 ( .A1(n694), .A2(n691), .ZN(n626) );
  NAND2_X1 U496 ( .A1(n425), .A2(n419), .ZN(n418) );
  AND2_X1 U497 ( .A1(n423), .A2(KEYINPUT34), .ZN(n419) );
  NOR2_X1 U498 ( .A1(n424), .A2(n415), .ZN(n411) );
  OR2_X1 U499 ( .A1(n421), .A2(KEYINPUT35), .ZN(n415) );
  NAND2_X1 U500 ( .A1(n371), .A2(n370), .ZN(n707) );
  NAND2_X1 U501 ( .A1(n386), .A2(n385), .ZN(n645) );
  AND2_X1 U502 ( .A1(n610), .A2(n387), .ZN(n386) );
  XNOR2_X1 U503 ( .A(n609), .B(n362), .ZN(n385) );
  INV_X1 U504 ( .A(n615), .ZN(n387) );
  XNOR2_X1 U505 ( .A(n491), .B(n489), .ZN(n737) );
  XNOR2_X1 U506 ( .A(n503), .B(n490), .ZN(n489) );
  XNOR2_X1 U507 ( .A(n498), .B(n357), .ZN(n734) );
  XNOR2_X1 U508 ( .A(n538), .B(n499), .ZN(n498) );
  XNOR2_X1 U509 ( .A(n540), .B(n535), .ZN(n499) );
  XNOR2_X1 U510 ( .A(n373), .B(n758), .ZN(n372) );
  XNOR2_X1 U511 ( .A(n408), .B(n407), .ZN(n373) );
  XNOR2_X1 U512 ( .A(n634), .B(KEYINPUT40), .ZN(n382) );
  AND2_X1 U513 ( .A1(n577), .A2(n434), .ZN(n432) );
  NAND2_X1 U514 ( .A1(n435), .A2(n393), .ZN(n392) );
  NOR2_X1 U515 ( .A1(n349), .A2(n588), .ZN(n664) );
  NOR2_X1 U516 ( .A1(n576), .A2(n703), .ZN(n587) );
  INV_X1 U517 ( .A(KEYINPUT63), .ZN(n461) );
  AND2_X1 U518 ( .A1(n769), .A2(n768), .ZN(n400) );
  INV_X1 U519 ( .A(KEYINPUT60), .ZN(n441) );
  INV_X1 U520 ( .A(KEYINPUT56), .ZN(n442) );
  AND2_X1 U521 ( .A1(n721), .A2(n749), .ZN(n403) );
  AND2_X1 U522 ( .A1(n438), .A2(n367), .ZN(n354) );
  OR2_X1 U523 ( .A1(n608), .A2(n521), .ZN(n355) );
  INV_X1 U524 ( .A(n583), .ZN(n370) );
  AND2_X1 U525 ( .A1(n368), .A2(n423), .ZN(n356) );
  INV_X1 U526 ( .A(n644), .ZN(n475) );
  AND2_X1 U527 ( .A1(n566), .A2(G217), .ZN(n357) );
  AND2_X1 U528 ( .A1(n774), .A2(n444), .ZN(n358) );
  AND2_X1 U529 ( .A1(n625), .A2(n698), .ZN(n359) );
  NAND2_X1 U530 ( .A1(n718), .A2(n427), .ZN(n360) );
  AND2_X1 U531 ( .A1(n644), .A2(n474), .ZN(n361) );
  XOR2_X1 U532 ( .A(KEYINPUT104), .B(KEYINPUT30), .Z(n362) );
  INV_X1 U533 ( .A(KEYINPUT35), .ZN(n474) );
  INV_X1 U534 ( .A(KEYINPUT34), .ZN(n427) );
  INV_X1 U535 ( .A(n739), .ZN(n446) );
  XOR2_X1 U536 ( .A(n381), .B(n724), .Z(n363) );
  XOR2_X1 U537 ( .A(n731), .B(n502), .Z(n364) );
  AND2_X1 U538 ( .A1(n542), .A2(G475), .ZN(n365) );
  AND2_X1 U539 ( .A1(n542), .A2(G210), .ZN(n366) );
  AND2_X1 U540 ( .A1(n542), .A2(G472), .ZN(n367) );
  NAND2_X1 U541 ( .A1(n416), .A2(n356), .ZN(n413) );
  NAND2_X1 U542 ( .A1(n426), .A2(KEYINPUT34), .ZN(n368) );
  NAND2_X1 U543 ( .A1(n682), .A2(n666), .ZN(n384) );
  INV_X1 U544 ( .A(n592), .ZN(n371) );
  XNOR2_X1 U545 ( .A(n374), .B(n560), .ZN(n376) );
  XNOR2_X1 U546 ( .A(n376), .B(n478), .ZN(n375) );
  NAND2_X1 U547 ( .A1(n582), .A2(n427), .ZN(n426) );
  BUF_X1 U548 ( .A(n597), .Z(n380) );
  BUF_X1 U549 ( .A(n725), .Z(n381) );
  BUF_X1 U550 ( .A(n611), .Z(n655) );
  XNOR2_X1 U551 ( .A(n457), .B(G143), .ZN(n528) );
  BUF_X1 U552 ( .A(G113), .Z(n457) );
  AND2_X1 U553 ( .A1(n575), .A2(KEYINPUT102), .ZN(n451) );
  BUF_X1 U554 ( .A(n575), .Z(n576) );
  XNOR2_X1 U555 ( .A(n382), .B(n777), .ZN(G33) );
  XNOR2_X1 U556 ( .A(n383), .B(KEYINPUT100), .ZN(n448) );
  NAND2_X1 U557 ( .A1(n384), .A2(n468), .ZN(n383) );
  NAND2_X1 U558 ( .A1(n388), .A2(n358), .ZN(n756) );
  NAND2_X1 U559 ( .A1(n390), .A2(n635), .ZN(n389) );
  INV_X1 U560 ( .A(n775), .ZN(n391) );
  NAND2_X1 U561 ( .A1(n394), .A2(n392), .ZN(n437) );
  INV_X1 U562 ( .A(n397), .ZN(n393) );
  NAND2_X1 U563 ( .A1(n451), .A2(KEYINPUT65), .ZN(n395) );
  NAND2_X1 U564 ( .A1(n397), .A2(KEYINPUT65), .ZN(n396) );
  NAND2_X1 U565 ( .A1(n437), .A2(n349), .ZN(n497) );
  NAND2_X1 U566 ( .A1(n497), .A2(n436), .ZN(n443) );
  XNOR2_X1 U567 ( .A(n443), .B(n496), .ZN(n597) );
  NAND2_X1 U568 ( .A1(n350), .A2(n359), .ZN(n398) );
  XNOR2_X1 U569 ( .A(n565), .B(n569), .ZN(n491) );
  NAND2_X1 U570 ( .A1(n494), .A2(n630), .ZN(n636) );
  INV_X1 U571 ( .A(n523), .ZN(n522) );
  NOR2_X1 U572 ( .A1(n737), .A2(G902), .ZN(n574) );
  XNOR2_X1 U573 ( .A(n727), .B(n460), .ZN(n730) );
  XNOR2_X1 U574 ( .A(n726), .B(n363), .ZN(n447) );
  XNOR2_X1 U575 ( .A(n732), .B(n364), .ZN(n445) );
  NAND2_X1 U576 ( .A1(n628), .A2(n688), .ZN(n609) );
  XNOR2_X1 U577 ( .A(n399), .B(KEYINPUT46), .ZN(n635) );
  XNOR2_X1 U578 ( .A(n400), .B(KEYINPUT125), .ZN(G72) );
  OR2_X1 U579 ( .A1(n577), .A2(n434), .ZN(n429) );
  XNOR2_X1 U580 ( .A(n404), .B(n442), .ZN(G51) );
  NAND2_X1 U581 ( .A1(n447), .A2(n446), .ZN(n404) );
  XNOR2_X1 U582 ( .A(n405), .B(n441), .ZN(G60) );
  NAND2_X1 U583 ( .A1(n445), .A2(n446), .ZN(n405) );
  NOR2_X1 U584 ( .A1(n663), .A2(n739), .ZN(n462) );
  INV_X1 U585 ( .A(n549), .ZN(n407) );
  NOR2_X1 U586 ( .A1(n422), .A2(n361), .ZN(n414) );
  NAND2_X1 U587 ( .A1(n420), .A2(n426), .ZN(n416) );
  NOR2_X1 U588 ( .A1(n718), .A2(n417), .ZN(n424) );
  NAND2_X1 U589 ( .A1(n425), .A2(KEYINPUT34), .ZN(n417) );
  NOR2_X1 U590 ( .A1(n718), .A2(n418), .ZN(n422) );
  INV_X1 U591 ( .A(n718), .ZN(n420) );
  INV_X1 U592 ( .A(n426), .ZN(n421) );
  INV_X1 U593 ( .A(n582), .ZN(n425) );
  NAND2_X1 U594 ( .A1(n492), .A2(n355), .ZN(n428) );
  NAND2_X1 U595 ( .A1(n576), .A2(n485), .ZN(n430) );
  INV_X1 U596 ( .A(n772), .ZN(n436) );
  NAND2_X1 U597 ( .A1(n486), .A2(n432), .ZN(n431) );
  INV_X1 U598 ( .A(n485), .ZN(n434) );
  NAND2_X1 U599 ( .A1(n750), .A2(n463), .ZN(n438) );
  XNOR2_X1 U600 ( .A(n353), .B(n439), .ZN(n722) );
  NAND2_X1 U601 ( .A1(n464), .A2(n354), .ZN(n662) );
  NAND2_X1 U602 ( .A1(n440), .A2(n366), .ZN(n726) );
  INV_X1 U603 ( .A(n576), .ZN(n486) );
  NOR2_X1 U604 ( .A1(n473), .A2(n594), .ZN(n593) );
  NAND2_X1 U605 ( .A1(n597), .A2(n593), .ZN(n449) );
  XNOR2_X1 U606 ( .A(n602), .B(n601), .ZN(n750) );
  NAND2_X1 U607 ( .A1(n448), .A2(n589), .ZN(n594) );
  NAND2_X1 U608 ( .A1(n449), .A2(n595), .ZN(n596) );
  NOR2_X1 U609 ( .A1(n600), .A2(n599), .ZN(n602) );
  OR2_X2 U610 ( .A1(n575), .A2(n454), .ZN(n450) );
  NAND2_X1 U611 ( .A1(n456), .A2(G217), .ZN(n736) );
  NAND2_X1 U612 ( .A1(n456), .A2(G478), .ZN(n733) );
  NAND2_X1 U613 ( .A1(n456), .A2(G469), .ZN(n727) );
  NAND2_X1 U614 ( .A1(n611), .A2(n688), .ZN(n516) );
  XNOR2_X1 U615 ( .A(n515), .B(n514), .ZN(n611) );
  XNOR2_X1 U616 ( .A(n462), .B(n461), .ZN(G57) );
  XNOR2_X2 U617 ( .A(n581), .B(KEYINPUT99), .ZN(n683) );
  XNOR2_X1 U618 ( .A(n529), .B(KEYINPUT16), .ZN(n482) );
  XNOR2_X1 U619 ( .A(n482), .B(n539), .ZN(n480) );
  XNOR2_X2 U620 ( .A(G122), .B(G104), .ZN(n529) );
  XNOR2_X2 U621 ( .A(G119), .B(G113), .ZN(n484) );
  NAND2_X1 U622 ( .A1(n762), .A2(G234), .ZN(n487) );
  XNOR2_X2 U623 ( .A(n488), .B(G953), .ZN(n762) );
  NAND2_X1 U624 ( .A1(n493), .A2(n492), .ZN(n637) );
  INV_X1 U625 ( .A(n636), .ZN(n493) );
  INV_X1 U626 ( .A(n497), .ZN(n670) );
  XNOR2_X1 U627 ( .A(n529), .B(n530), .ZN(n531) );
  NOR2_X1 U628 ( .A1(n762), .A2(G952), .ZN(n739) );
  XOR2_X1 U629 ( .A(KEYINPUT72), .B(KEYINPUT18), .Z(n500) );
  AND2_X1 U630 ( .A1(G214), .A2(n557), .ZN(n501) );
  XNOR2_X1 U631 ( .A(KEYINPUT119), .B(KEYINPUT59), .ZN(n502) );
  XOR2_X1 U632 ( .A(n568), .B(n567), .Z(n503) );
  INV_X1 U633 ( .A(KEYINPUT48), .ZN(n650) );
  XNOR2_X1 U634 ( .A(n650), .B(KEYINPUT80), .ZN(n651) );
  INV_X1 U635 ( .A(KEYINPUT85), .ZN(n504) );
  INV_X1 U636 ( .A(KEYINPUT68), .ZN(n552) );
  INV_X1 U637 ( .A(KEYINPUT97), .ZN(n578) );
  NAND2_X1 U638 ( .A1(G214), .A2(n513), .ZN(n688) );
  XOR2_X1 U639 ( .A(KEYINPUT69), .B(KEYINPUT3), .Z(n505) );
  XNOR2_X1 U640 ( .A(n740), .B(n546), .ZN(n512) );
  XNOR2_X1 U641 ( .A(KEYINPUT70), .B(n742), .ZN(n549) );
  NAND2_X1 U642 ( .A1(G224), .A2(n762), .ZN(n507) );
  XNOR2_X1 U643 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U644 ( .A(n510), .B(n509), .Z(n511) );
  XNOR2_X1 U645 ( .A(n512), .B(n511), .ZN(n725) );
  NOR2_X1 U646 ( .A1(n725), .A2(n542), .ZN(n515) );
  NAND2_X1 U647 ( .A1(G210), .A2(n513), .ZN(n514) );
  XOR2_X1 U648 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n518) );
  XNOR2_X1 U649 ( .A(n518), .B(n517), .ZN(n519) );
  NAND2_X1 U650 ( .A1(G952), .A2(n519), .ZN(n716) );
  NOR2_X1 U651 ( .A1(G953), .A2(n716), .ZN(n608) );
  AND2_X1 U652 ( .A1(G902), .A2(n519), .ZN(n604) );
  INV_X1 U653 ( .A(G953), .ZN(n749) );
  NOR2_X1 U654 ( .A1(G898), .A2(n749), .ZN(n744) );
  NAND2_X1 U655 ( .A1(n604), .A2(n744), .ZN(n520) );
  XOR2_X1 U656 ( .A(KEYINPUT88), .B(n520), .Z(n521) );
  XNOR2_X1 U657 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n533) );
  XNOR2_X1 U658 ( .A(n757), .B(n525), .ZN(n526) );
  XNOR2_X1 U659 ( .A(KEYINPUT12), .B(n526), .ZN(n532) );
  XNOR2_X1 U660 ( .A(n551), .B(n528), .ZN(n530) );
  XOR2_X1 U661 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n534) );
  XNOR2_X1 U662 ( .A(n536), .B(G134), .ZN(n537) );
  XNOR2_X1 U663 ( .A(n537), .B(G122), .ZN(n538) );
  XNOR2_X1 U664 ( .A(n539), .B(KEYINPUT98), .ZN(n540) );
  NOR2_X1 U665 ( .A1(G902), .A2(n734), .ZN(n541) );
  XNOR2_X1 U666 ( .A(G478), .B(n541), .ZN(n579) );
  INV_X1 U667 ( .A(n579), .ZN(n591) );
  XOR2_X1 U668 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n544) );
  INV_X1 U669 ( .A(n542), .ZN(n658) );
  NAND2_X1 U670 ( .A1(G234), .A2(n658), .ZN(n543) );
  XNOR2_X1 U671 ( .A(n544), .B(n543), .ZN(n571) );
  NAND2_X1 U672 ( .A1(n571), .A2(G221), .ZN(n545) );
  XOR2_X1 U673 ( .A(KEYINPUT21), .B(n545), .Z(n698) );
  INV_X1 U674 ( .A(n698), .ZN(n585) );
  NAND2_X1 U675 ( .A1(G227), .A2(n762), .ZN(n547) );
  NAND2_X1 U676 ( .A1(n557), .A2(G210), .ZN(n558) );
  XNOR2_X1 U677 ( .A(n559), .B(n558), .ZN(n560) );
  NOR2_X1 U678 ( .A1(n660), .A2(G902), .ZN(n562) );
  XNOR2_X1 U679 ( .A(n564), .B(n563), .ZN(n570) );
  XNOR2_X1 U680 ( .A(n757), .B(KEYINPUT89), .ZN(n565) );
  NAND2_X1 U681 ( .A1(G221), .A2(n566), .ZN(n569) );
  NAND2_X1 U682 ( .A1(n571), .A2(G217), .ZN(n572) );
  XNOR2_X1 U683 ( .A(n590), .B(n578), .ZN(n580) );
  NAND2_X1 U684 ( .A1(n580), .A2(n579), .ZN(n678) );
  NOR2_X1 U685 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U686 ( .A1(n585), .A2(n349), .ZN(n702) );
  NAND2_X1 U687 ( .A1(n630), .A2(n702), .ZN(n603) );
  NOR2_X1 U688 ( .A1(n582), .A2(n603), .ZN(n586) );
  NAND2_X1 U689 ( .A1(n586), .A2(n583), .ZN(n666) );
  NAND2_X1 U690 ( .A1(n587), .A2(n616), .ZN(n588) );
  INV_X1 U691 ( .A(n664), .ZN(n589) );
  NAND2_X1 U692 ( .A1(n591), .A2(n590), .ZN(n644) );
  XNOR2_X1 U693 ( .A(n596), .B(KEYINPUT81), .ZN(n600) );
  NAND2_X1 U694 ( .A1(n380), .A2(n773), .ZN(n598) );
  NOR2_X1 U695 ( .A1(n598), .A2(KEYINPUT44), .ZN(n599) );
  NOR2_X1 U696 ( .A1(KEYINPUT2), .A2(KEYINPUT79), .ZN(n657) );
  INV_X1 U697 ( .A(n603), .ZN(n610) );
  INV_X1 U698 ( .A(n762), .ZN(n605) );
  NAND2_X1 U699 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U700 ( .A1(G900), .A2(n606), .ZN(n607) );
  NOR2_X1 U701 ( .A1(n608), .A2(n607), .ZN(n615) );
  INV_X1 U702 ( .A(n689), .ZN(n612) );
  XNOR2_X1 U703 ( .A(n613), .B(KEYINPUT39), .ZN(n633) );
  NOR2_X1 U704 ( .A1(n633), .A2(n683), .ZN(n686) );
  XNOR2_X1 U705 ( .A(KEYINPUT107), .B(KEYINPUT36), .ZN(n622) );
  NAND2_X1 U706 ( .A1(n349), .A2(n698), .ZN(n614) );
  NOR2_X1 U707 ( .A1(n615), .A2(n614), .ZN(n627) );
  INV_X1 U708 ( .A(n616), .ZN(n617) );
  NAND2_X1 U709 ( .A1(n627), .A2(n617), .ZN(n618) );
  NOR2_X1 U710 ( .A1(n678), .A2(n618), .ZN(n619) );
  NAND2_X1 U711 ( .A1(n619), .A2(n688), .ZN(n652) );
  INV_X1 U712 ( .A(n655), .ZN(n620) );
  NOR2_X1 U713 ( .A1(n652), .A2(n620), .ZN(n621) );
  XOR2_X1 U714 ( .A(n622), .B(n621), .Z(n623) );
  NAND2_X1 U715 ( .A1(n703), .A2(n623), .ZN(n624) );
  XNOR2_X1 U716 ( .A(KEYINPUT108), .B(n624), .ZN(n775) );
  NAND2_X1 U717 ( .A1(n689), .A2(n688), .ZN(n694) );
  INV_X1 U718 ( .A(n625), .ZN(n691) );
  XNOR2_X1 U719 ( .A(n626), .B(KEYINPUT41), .ZN(n717) );
  NAND2_X1 U720 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U721 ( .A1(n717), .A2(n636), .ZN(n631) );
  XNOR2_X1 U722 ( .A(n631), .B(KEYINPUT42), .ZN(n632) );
  XNOR2_X1 U723 ( .A(KEYINPUT106), .B(n632), .ZN(n770) );
  NOR2_X1 U724 ( .A1(n633), .A2(n678), .ZN(n634) );
  INV_X1 U725 ( .A(KEYINPUT47), .ZN(n638) );
  XNOR2_X1 U726 ( .A(n637), .B(KEYINPUT75), .ZN(n640) );
  INV_X1 U727 ( .A(n640), .ZN(n675) );
  NAND2_X1 U728 ( .A1(n638), .A2(n675), .ZN(n643) );
  NAND2_X1 U729 ( .A1(n638), .A2(KEYINPUT76), .ZN(n639) );
  XOR2_X1 U730 ( .A(n639), .B(n693), .Z(n641) );
  NAND2_X1 U731 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U732 ( .A1(n643), .A2(n642), .ZN(n647) );
  NOR2_X1 U733 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U734 ( .A1(n655), .A2(n646), .ZN(n674) );
  NAND2_X1 U735 ( .A1(n647), .A2(n674), .ZN(n648) );
  XOR2_X1 U736 ( .A(n648), .B(KEYINPUT71), .Z(n649) );
  NOR2_X1 U737 ( .A1(n703), .A2(n652), .ZN(n653) );
  XNOR2_X1 U738 ( .A(n653), .B(KEYINPUT43), .ZN(n654) );
  NOR2_X1 U739 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U740 ( .A(KEYINPUT103), .B(n656), .ZN(n774) );
  XOR2_X1 U741 ( .A(KEYINPUT62), .B(KEYINPUT109), .Z(n659) );
  XNOR2_X1 U742 ( .A(n662), .B(n661), .ZN(n663) );
  XOR2_X1 U743 ( .A(G101), .B(n664), .Z(G3) );
  NOR2_X1 U744 ( .A1(n678), .A2(n666), .ZN(n665) );
  XOR2_X1 U745 ( .A(n458), .B(n665), .Z(G6) );
  NOR2_X1 U746 ( .A1(n683), .A2(n666), .ZN(n668) );
  XNOR2_X1 U747 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n667) );
  XNOR2_X1 U748 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U749 ( .A(G107), .B(n669), .ZN(G9) );
  XOR2_X1 U750 ( .A(G110), .B(n670), .Z(G12) );
  NOR2_X1 U751 ( .A1(n675), .A2(n683), .ZN(n672) );
  XNOR2_X1 U752 ( .A(KEYINPUT29), .B(KEYINPUT110), .ZN(n671) );
  XNOR2_X1 U753 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U754 ( .A(G128), .B(n673), .ZN(G30) );
  XNOR2_X1 U755 ( .A(G143), .B(n674), .ZN(G45) );
  NOR2_X1 U756 ( .A1(n678), .A2(n675), .ZN(n677) );
  XNOR2_X1 U757 ( .A(G146), .B(KEYINPUT111), .ZN(n676) );
  XNOR2_X1 U758 ( .A(n677), .B(n676), .ZN(G48) );
  NOR2_X1 U759 ( .A1(n678), .A2(n682), .ZN(n680) );
  XNOR2_X1 U760 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n679) );
  XNOR2_X1 U761 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U762 ( .A(n457), .B(n681), .ZN(G15) );
  NOR2_X1 U763 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U764 ( .A(KEYINPUT114), .B(n684), .Z(n685) );
  XNOR2_X1 U765 ( .A(G116), .B(n685), .ZN(G18) );
  XNOR2_X1 U766 ( .A(G134), .B(n686), .ZN(n687) );
  XNOR2_X1 U767 ( .A(n687), .B(KEYINPUT115), .ZN(G36) );
  NOR2_X1 U768 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U769 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U770 ( .A(n692), .B(KEYINPUT118), .ZN(n696) );
  NOR2_X1 U771 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U772 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U773 ( .A1(n697), .A2(n718), .ZN(n713) );
  NOR2_X1 U774 ( .A1(n698), .A2(n584), .ZN(n699) );
  XOR2_X1 U775 ( .A(KEYINPUT49), .B(n699), .Z(n700) );
  NOR2_X1 U776 ( .A1(n370), .A2(n700), .ZN(n701) );
  XNOR2_X1 U777 ( .A(n701), .B(KEYINPUT116), .ZN(n706) );
  OR2_X1 U778 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U779 ( .A(KEYINPUT50), .B(n704), .ZN(n705) );
  NAND2_X1 U780 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U781 ( .A1(n708), .A2(n707), .ZN(n710) );
  XOR2_X1 U782 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n709) );
  XNOR2_X1 U783 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U784 ( .A1(n711), .A2(n717), .ZN(n712) );
  NOR2_X1 U785 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U786 ( .A(n714), .B(KEYINPUT52), .ZN(n715) );
  NOR2_X1 U787 ( .A1(n716), .A2(n715), .ZN(n720) );
  NOR2_X1 U788 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U790 ( .A(n723), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U791 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n724) );
  XOR2_X1 U792 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n728) );
  NOR2_X1 U793 ( .A1(n739), .A2(n730), .ZN(G54) );
  XNOR2_X1 U794 ( .A(n733), .B(n734), .ZN(n735) );
  NOR2_X1 U795 ( .A1(n735), .A2(n739), .ZN(G63) );
  XNOR2_X1 U796 ( .A(n736), .B(n737), .ZN(n738) );
  NOR2_X1 U797 ( .A1(n738), .A2(n739), .ZN(G66) );
  XOR2_X1 U798 ( .A(n352), .B(G101), .Z(n741) );
  XNOR2_X1 U799 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U800 ( .A1(n744), .A2(n743), .ZN(n755) );
  NAND2_X1 U801 ( .A1(G224), .A2(G953), .ZN(n745) );
  XNOR2_X1 U802 ( .A(n745), .B(KEYINPUT61), .ZN(n746) );
  XNOR2_X1 U803 ( .A(KEYINPUT120), .B(n746), .ZN(n747) );
  NAND2_X1 U804 ( .A1(n747), .A2(G898), .ZN(n748) );
  XNOR2_X1 U805 ( .A(n748), .B(KEYINPUT121), .ZN(n752) );
  AND2_X1 U806 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U807 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U808 ( .A(n753), .B(KEYINPUT122), .Z(n754) );
  XNOR2_X1 U809 ( .A(n755), .B(n754), .ZN(G69) );
  XNOR2_X1 U810 ( .A(n757), .B(KEYINPUT123), .ZN(n759) );
  XNOR2_X1 U811 ( .A(n758), .B(n759), .ZN(n760) );
  XOR2_X1 U812 ( .A(n761), .B(n760), .Z(n765) );
  NAND2_X1 U813 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U814 ( .A(n764), .B(KEYINPUT124), .ZN(n769) );
  XNOR2_X1 U815 ( .A(G227), .B(n765), .ZN(n766) );
  NAND2_X1 U816 ( .A1(n766), .A2(G900), .ZN(n767) );
  NAND2_X1 U817 ( .A1(n767), .A2(G953), .ZN(n768) );
  XOR2_X1 U818 ( .A(n770), .B(G137), .Z(G39) );
  XOR2_X1 U819 ( .A(G119), .B(KEYINPUT126), .Z(n771) );
  XNOR2_X1 U820 ( .A(n772), .B(n771), .ZN(G21) );
  XNOR2_X1 U821 ( .A(G122), .B(n773), .ZN(G24) );
  XNOR2_X1 U822 ( .A(G140), .B(n774), .ZN(G42) );
  XOR2_X1 U823 ( .A(G125), .B(n775), .Z(n776) );
  XNOR2_X1 U824 ( .A(KEYINPUT37), .B(n776), .ZN(G27) );
  XNOR2_X1 U825 ( .A(G131), .B(KEYINPUT127), .ZN(n777) );
endmodule

