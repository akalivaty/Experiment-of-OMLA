//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT65), .Z(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT67), .Z(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n209), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT68), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT1), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n221), .A2(new_n222), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT66), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G20), .ZN(new_n227));
  AND2_X1   g0027(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR4_X1   g0031(.A1(new_n213), .A2(new_n223), .A3(new_n224), .A4(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G68), .Z(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND2_X1  g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G222), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n249), .ZN(new_n258));
  INV_X1    g0058(.A(G223), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(G1698), .ZN(new_n260));
  OAI221_X1 g0060(.A(new_n254), .B1(new_n202), .B2(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n262), .A2(new_n268), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(G226), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n263), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G190), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(G200), .B2(new_n273), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G150), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n228), .A2(G33), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  OAI221_X1 g0080(.A(new_n278), .B1(new_n207), .B2(new_n201), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n229), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(new_n283), .ZN(new_n287));
  INV_X1    g0087(.A(G50), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n206), .B2(G20), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n287), .A2(new_n289), .B1(new_n288), .B2(new_n286), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT69), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n291), .B(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n276), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n273), .A2(new_n298), .B1(new_n284), .B2(new_n290), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(G179), .B2(new_n273), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G87), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n256), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT72), .B(G33), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n257), .B1(new_n304), .B2(new_n255), .ZN(new_n305));
  INV_X1    g0105(.A(G226), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G1698), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(G223), .B2(G1698), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n303), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n262), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT74), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT74), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n256), .A2(KEYINPUT72), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT72), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n308), .B1(new_n318), .B2(new_n257), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n313), .B(new_n262), .C1(new_n319), .C2(new_n303), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n271), .A2(G232), .ZN(new_n321));
  INV_X1    g0121(.A(G179), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n269), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n312), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n305), .A2(new_n309), .ZN(new_n325));
  INV_X1    g0125(.A(new_n303), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n311), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n269), .A2(new_n321), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n298), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT75), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n287), .ZN(new_n333));
  INV_X1    g0133(.A(new_n280), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n206), .A2(G20), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n333), .A2(new_n336), .B1(new_n285), .B2(new_n334), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n250), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n228), .B(new_n340), .C1(KEYINPUT3), .C2(new_n317), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n257), .A2(new_n207), .A3(new_n249), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n342), .A2(KEYINPUT73), .A3(new_n339), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT73), .B1(new_n342), .B2(new_n339), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n341), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G68), .ZN(new_n346));
  INV_X1    g0146(.A(G58), .ZN(new_n347));
  INV_X1    g0147(.A(G68), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(G58), .A2(G68), .ZN(new_n350));
  OAI21_X1  g0150(.A(G20), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n277), .A2(G159), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT16), .B1(new_n346), .B2(new_n354), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n351), .A2(KEYINPUT16), .A3(new_n352), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n251), .B1(new_n317), .B2(KEYINPUT3), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n339), .B1(new_n357), .B2(new_n207), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n225), .A2(new_n227), .A3(new_n339), .ZN(new_n359));
  OAI21_X1  g0159(.A(G68), .B1(new_n305), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n356), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n283), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n338), .B1(new_n355), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n324), .A2(KEYINPUT75), .A3(new_n329), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n332), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT18), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n363), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT77), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n269), .A2(new_n321), .A3(new_n274), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n312), .A2(new_n320), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G200), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n327), .B2(new_n328), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n368), .A2(KEYINPUT76), .A3(new_n369), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT17), .ZN(new_n376));
  INV_X1    g0176(.A(new_n283), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT7), .B1(new_n305), .B2(G20), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n357), .A2(new_n339), .A3(new_n228), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(G68), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n377), .B1(new_n380), .B2(new_n356), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n353), .B1(new_n345), .B2(G68), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n381), .B1(KEYINPUT16), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(new_n374), .A3(new_n338), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT76), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n376), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n375), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n384), .A2(KEYINPUT77), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n376), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n367), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G1698), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n258), .A2(G226), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G97), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n393), .B(new_n394), .C1(new_n260), .C2(new_n234), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n262), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT70), .ZN(new_n397));
  INV_X1    g0197(.A(new_n268), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n311), .A2(G238), .A3(new_n398), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n269), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n397), .B1(new_n269), .B2(new_n399), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n396), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT13), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT13), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n404), .B(new_n396), .C1(new_n400), .C2(new_n401), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G169), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT14), .ZN(new_n408));
  INV_X1    g0208(.A(new_n401), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n269), .A2(new_n399), .A3(new_n397), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT71), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(new_n404), .A4(new_n396), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n405), .A2(KEYINPUT71), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(G179), .A4(new_n403), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT14), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n406), .A2(new_n416), .A3(G169), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n408), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n277), .A2(G50), .B1(G20), .B2(new_n348), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n279), .B2(new_n202), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n420), .A2(new_n283), .ZN(new_n421));
  OR2_X1    g0221(.A1(new_n421), .A2(KEYINPUT11), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(KEYINPUT11), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n286), .A2(new_n348), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT12), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n287), .A2(G68), .A3(new_n335), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n422), .A2(new_n423), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n427), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n406), .A2(G200), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n413), .A2(new_n414), .A3(G190), .A4(new_n403), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n271), .A2(G244), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n253), .A2(G232), .ZN(new_n435));
  INV_X1    g0235(.A(G107), .ZN(new_n436));
  INV_X1    g0236(.A(G238), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n435), .B1(new_n436), .B2(new_n258), .C1(new_n437), .C2(new_n260), .ZN(new_n438));
  AOI211_X1 g0238(.A(new_n270), .B(new_n434), .C1(new_n438), .C2(new_n262), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n439), .A2(new_n322), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n225), .A2(new_n227), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n334), .A2(new_n277), .B1(new_n441), .B2(G77), .ZN(new_n442));
  XNOR2_X1  g0242(.A(KEYINPUT15), .B(G87), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n279), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n283), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n335), .A2(G77), .ZN(new_n446));
  OAI221_X1 g0246(.A(new_n445), .B1(G77), .B2(new_n285), .C1(new_n333), .C2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n439), .B2(G169), .ZN(new_n448));
  OR2_X1    g0248(.A1(new_n440), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n447), .B1(new_n439), .B2(G190), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n372), .B2(new_n439), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NOR4_X1   g0252(.A1(new_n301), .A2(new_n391), .A3(new_n433), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n283), .B1(new_n207), .B2(G116), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G283), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(G33), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT83), .ZN(new_n459));
  OR3_X1    g0259(.A1(new_n441), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n441), .B2(new_n458), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n455), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n462), .A2(KEYINPUT84), .A3(KEYINPUT20), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n286), .A2(G116), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n287), .B1(G1), .B2(new_n256), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(G116), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n267), .A2(G1), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT5), .B(G41), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n311), .A2(G274), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n262), .B1(new_n468), .B2(new_n469), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G270), .ZN(new_n472));
  MUX2_X1   g0272(.A(G257), .B(G264), .S(G1698), .Z(new_n473));
  AOI22_X1  g0273(.A1(new_n305), .A2(new_n473), .B1(G303), .B2(new_n252), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n470), .B(new_n472), .C1(new_n474), .C2(new_n311), .ZN(new_n475));
  OR2_X1    g0275(.A1(new_n475), .A2(new_n274), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT84), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n462), .B2(KEYINPUT20), .ZN(new_n478));
  INV_X1    g0278(.A(new_n455), .ZN(new_n479));
  INV_X1    g0279(.A(new_n461), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n441), .A2(new_n458), .A3(new_n459), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT20), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n475), .A2(G200), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n467), .A2(new_n476), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT85), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n475), .A2(G169), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(new_n467), .B2(new_n485), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n467), .A2(new_n485), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n475), .A2(new_n322), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n491), .A2(KEYINPUT21), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n490), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n478), .A2(new_n484), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n482), .A2(new_n477), .A3(new_n483), .ZN(new_n497));
  INV_X1    g0297(.A(new_n465), .ZN(new_n498));
  INV_X1    g0298(.A(G116), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n497), .B1(new_n464), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n495), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT21), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n494), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(G250), .A2(G1698), .ZN(new_n506));
  INV_X1    g0306(.A(G257), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(G1698), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n305), .A2(new_n508), .B1(G294), .B2(new_n317), .ZN(new_n509));
  OR2_X1    g0309(.A1(new_n509), .A2(new_n311), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n469), .A2(new_n468), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(new_n311), .A3(G264), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT88), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n471), .A2(KEYINPUT88), .A3(G264), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n510), .A2(new_n470), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n509), .A2(new_n311), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n470), .A2(new_n512), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n517), .A2(new_n372), .B1(new_n520), .B2(new_n274), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n305), .A2(KEYINPUT22), .A3(G87), .A4(new_n228), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT22), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n252), .B2(new_n302), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n317), .A2(new_n207), .A3(G116), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n441), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n436), .A2(G20), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(KEYINPUT23), .B1(KEYINPUT86), .B2(KEYINPUT24), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n526), .A2(new_n527), .A3(new_n529), .A4(new_n531), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n524), .A2(new_n532), .B1(KEYINPUT86), .B2(KEYINPUT24), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n526), .A2(new_n529), .A3(new_n531), .ZN(new_n534));
  NOR2_X1   g0334(.A1(KEYINPUT86), .A2(KEYINPUT24), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n534), .A2(new_n535), .A3(new_n523), .A4(new_n527), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n377), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n206), .A2(G13), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT25), .ZN(new_n539));
  AOI211_X1 g0339(.A(new_n538), .B(new_n530), .C1(KEYINPUT87), .C2(new_n539), .ZN(new_n540));
  OR3_X1    g0340(.A1(new_n540), .A2(KEYINPUT87), .A3(new_n539), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(KEYINPUT87), .B2(new_n539), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n541), .B(new_n542), .C1(new_n436), .C2(new_n465), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n522), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n510), .A2(G179), .A3(new_n470), .A4(new_n516), .ZN(new_n546));
  OAI21_X1  g0346(.A(G169), .B1(new_n518), .B2(new_n519), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n537), .B2(new_n543), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n489), .A2(new_n505), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n511), .A2(new_n311), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n470), .B1(new_n552), .B2(new_n507), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT79), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n471), .A2(G257), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT79), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(new_n470), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n258), .A2(KEYINPUT4), .A3(G244), .A4(new_n392), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n258), .A2(G250), .A3(G1698), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n456), .A3(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT4), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n305), .A2(G244), .A3(new_n392), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n554), .B(new_n557), .C1(new_n563), .C2(new_n311), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G200), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n274), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n285), .A2(G97), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n498), .B2(G97), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n277), .A2(G77), .ZN(new_n569));
  XNOR2_X1  g0369(.A(G97), .B(G107), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(KEYINPUT78), .B2(KEYINPUT6), .ZN(new_n571));
  NOR2_X1   g0371(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(KEYINPUT6), .B2(new_n457), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n571), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n569), .B1(new_n574), .B2(new_n228), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(G107), .B2(new_n345), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n568), .B1(new_n576), .B2(new_n377), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n566), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT80), .B1(new_n564), .B2(G179), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n554), .A2(new_n557), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n562), .A2(new_n561), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n262), .B1(new_n581), .B2(new_n560), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT80), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n580), .A2(new_n582), .A3(new_n583), .A4(new_n322), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n345), .A2(G107), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n283), .B1(new_n586), .B2(new_n575), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(new_n568), .B1(new_n564), .B2(new_n298), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n565), .A2(new_n578), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n305), .A2(G68), .A3(new_n228), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n225), .B(new_n227), .C1(new_n591), .C2(new_n394), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n302), .A2(new_n457), .A3(new_n436), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n279), .A2(new_n457), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n590), .B(new_n594), .C1(new_n595), .C2(KEYINPUT19), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n283), .ZN(new_n597));
  INV_X1    g0397(.A(new_n443), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(new_n285), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n498), .A2(new_n598), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n597), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT81), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n468), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n605), .A2(G250), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n311), .A2(new_n606), .B1(new_n265), .B2(new_n468), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n437), .A2(G1698), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n305), .A2(new_n608), .B1(G116), .B2(new_n317), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n305), .A2(G244), .A3(G1698), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(G179), .B(new_n607), .C1(new_n611), .C2(new_n311), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n311), .B1(new_n609), .B2(new_n610), .ZN(new_n613));
  INV_X1    g0413(.A(new_n607), .ZN(new_n614));
  OAI21_X1  g0414(.A(G169), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n602), .A2(new_n603), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n613), .A2(new_n274), .A3(new_n614), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n613), .A2(new_n614), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n619), .B2(G200), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n465), .A2(new_n302), .ZN(new_n621));
  AOI211_X1 g0421(.A(new_n599), .B(new_n621), .C1(new_n596), .C2(new_n283), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n604), .A2(new_n616), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n589), .A2(KEYINPUT82), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT82), .B1(new_n589), .B2(new_n623), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n551), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n454), .A2(new_n626), .ZN(G372));
  INV_X1    g0427(.A(new_n300), .ZN(new_n628));
  INV_X1    g0428(.A(new_n449), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n629), .A2(new_n432), .B1(new_n418), .B2(new_n427), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n375), .A2(new_n386), .B1(new_n388), .B2(new_n376), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n367), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n628), .B1(new_n632), .B2(new_n297), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n585), .A2(new_n588), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n612), .A2(new_n615), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n602), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n618), .A2(G190), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n372), .B2(new_n618), .ZN(new_n639));
  INV_X1    g0439(.A(new_n622), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n634), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT90), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g0444(.A(KEYINPUT90), .B(new_n634), .C1(new_n635), .C2(new_n641), .ZN(new_n645));
  INV_X1    g0445(.A(new_n635), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(new_n623), .A3(KEYINPUT26), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n637), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n578), .A2(new_n565), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n620), .A2(new_n622), .B1(new_n636), .B2(new_n602), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n635), .A2(new_n650), .A3(new_n545), .A4(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT89), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n549), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n548), .B(KEYINPUT89), .C1(new_n537), .C2(new_n543), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n504), .B(new_n494), .C1(new_n654), .C2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n649), .B1(new_n652), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n648), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n633), .B1(new_n454), .B2(new_n659), .ZN(G369));
  OR3_X1    g0460(.A1(new_n441), .A2(KEYINPUT27), .A3(new_n538), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT27), .B1(new_n441), .B2(new_n538), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G343), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT91), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n492), .A2(new_n665), .ZN(new_n666));
  OR3_X1    g0466(.A1(new_n489), .A2(new_n505), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n505), .A2(new_n666), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g0469(.A(KEYINPUT92), .B(G330), .Z(new_n670));
  AND2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n550), .ZN(new_n672));
  INV_X1    g0472(.A(new_n665), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n672), .B1(new_n544), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n549), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  OR3_X1    g0476(.A1(new_n654), .A2(new_n656), .A3(new_n665), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n665), .B1(new_n494), .B2(new_n504), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n672), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n210), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n206), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n593), .A2(G116), .ZN(new_n684));
  INV_X1    g0484(.A(new_n230), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n683), .A2(new_n684), .B1(new_n685), .B2(new_n682), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT28), .Z(new_n687));
  AOI21_X1  g0487(.A(new_n665), .B1(new_n648), .B2(new_n658), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(KEYINPUT29), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT93), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT93), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n688), .B2(KEYINPUT29), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n646), .A2(new_n623), .A3(new_n634), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT26), .B1(new_n635), .B2(new_n641), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(new_n694), .A3(new_n637), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n521), .A2(new_n537), .A3(new_n543), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n641), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n491), .A2(KEYINPUT21), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n492), .A2(new_n493), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n504), .A2(new_n698), .A3(new_n699), .A4(new_n549), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n697), .A2(new_n589), .A3(new_n700), .ZN(new_n701));
  OAI211_X1 g0501(.A(KEYINPUT29), .B(new_n673), .C1(new_n695), .C2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n690), .A2(new_n692), .A3(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n551), .B(new_n673), .C1(new_n624), .C2(new_n625), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n474), .A2(new_n311), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n618), .A2(new_n705), .A3(new_n472), .ZN(new_n706));
  INV_X1    g0506(.A(new_n564), .ZN(new_n707));
  INV_X1    g0507(.A(new_n546), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n706), .A2(KEYINPUT30), .A3(new_n708), .A4(new_n707), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n475), .A2(new_n322), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n619), .A2(new_n713), .A3(new_n564), .A4(new_n517), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n715), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT31), .B1(new_n715), .B2(new_n665), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n704), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n670), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n703), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n687), .B1(new_n721), .B2(G1), .ZN(G364));
  INV_X1    g0522(.A(G13), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n441), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G45), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n683), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n671), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n670), .B2(new_n669), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n681), .A2(new_n252), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n730), .A2(G355), .B1(new_n499), .B2(new_n681), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n681), .A2(new_n305), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(G45), .B2(new_n230), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n247), .A2(new_n267), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n229), .B1(G20), .B2(new_n298), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n228), .A2(new_n322), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n274), .A2(G200), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n372), .A2(G190), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  XNOR2_X1  g0549(.A(KEYINPUT33), .B(G317), .ZN(new_n750));
  AOI22_X1  g0550(.A1(G322), .A2(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G283), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n441), .A2(new_n322), .A3(new_n747), .ZN(new_n753));
  INV_X1    g0553(.A(G311), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G190), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n742), .A2(new_n755), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n751), .B1(new_n752), .B2(new_n753), .C1(new_n754), .C2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n441), .A2(new_n322), .A3(new_n755), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n441), .B1(new_n745), .B2(G179), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n759), .A2(G329), .B1(G294), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n274), .A2(new_n372), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(G20), .A3(new_n322), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n258), .B1(new_n764), .B2(G303), .ZN(new_n765));
  INV_X1    g0565(.A(G326), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n742), .A2(new_n762), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n761), .B(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n757), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT95), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(KEYINPUT95), .ZN(new_n771));
  INV_X1    g0571(.A(new_n767), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G50), .ZN(new_n773));
  INV_X1    g0573(.A(G159), .ZN(new_n774));
  OR3_X1    g0574(.A1(new_n758), .A2(KEYINPUT32), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(KEYINPUT32), .B1(new_n758), .B2(new_n774), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n252), .B1(new_n764), .B2(G87), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n773), .A2(new_n775), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n756), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G58), .A2(new_n746), .B1(new_n779), .B2(G77), .ZN(new_n780));
  INV_X1    g0580(.A(new_n753), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n749), .A2(G68), .B1(G107), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n760), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n783), .A2(KEYINPUT94), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(KEYINPUT94), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n780), .B(new_n782), .C1(new_n457), .C2(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n770), .B(new_n771), .C1(new_n778), .C2(new_n787), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n726), .B(new_n741), .C1(new_n788), .C2(new_n739), .ZN(new_n789));
  INV_X1    g0589(.A(new_n738), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n789), .B1(new_n669), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n729), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  NOR2_X1   g0593(.A1(new_n449), .A2(new_n665), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n665), .A2(new_n447), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT96), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(KEYINPUT96), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n796), .A2(new_n451), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n794), .B1(new_n798), .B2(new_n449), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n688), .B(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n727), .B1(new_n800), .B2(new_n720), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n720), .B2(new_n800), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G143), .A2(new_n746), .B1(new_n772), .B2(G137), .ZN(new_n803));
  INV_X1    g0603(.A(G150), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n804), .B2(new_n748), .C1(new_n774), .C2(new_n756), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT34), .Z(new_n806));
  OAI221_X1 g0606(.A(new_n305), .B1(new_n288), .B2(new_n763), .C1(new_n783), .C2(new_n347), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n753), .A2(new_n348), .ZN(new_n808));
  INV_X1    g0608(.A(G132), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n758), .A2(new_n809), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n806), .A2(new_n807), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n781), .A2(G87), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n812), .B1(new_n754), .B2(new_n758), .C1(new_n748), .C2(new_n752), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n252), .B1(new_n763), .B2(new_n436), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n772), .B2(G303), .ZN(new_n815));
  INV_X1    g0615(.A(G294), .ZN(new_n816));
  INV_X1    g0616(.A(new_n746), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n499), .B2(new_n756), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n786), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n813), .B(new_n818), .C1(G97), .C2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n739), .B1(new_n811), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n739), .A2(new_n736), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n726), .B1(new_n202), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n821), .B(new_n823), .C1(new_n799), .C2(new_n737), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n802), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G384));
  NOR2_X1   g0626(.A1(new_n724), .A2(new_n206), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n427), .A2(new_n665), .ZN(new_n828));
  INV_X1    g0628(.A(new_n415), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n416), .B1(new_n406), .B2(G169), .ZN(new_n830));
  AOI211_X1 g0630(.A(KEYINPUT14), .B(new_n298), .C1(new_n403), .C2(new_n405), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n432), .B(new_n828), .C1(new_n832), .C2(new_n429), .ZN(new_n833));
  INV_X1    g0633(.A(new_n432), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n427), .B(new_n665), .C1(new_n418), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n799), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n704), .B2(new_n718), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT38), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n363), .A2(new_n663), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n367), .B2(new_n390), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n371), .A2(new_n373), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n385), .B1(new_n363), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(KEYINPUT37), .B1(new_n363), .B2(new_n663), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n383), .A2(new_n374), .A3(KEYINPUT76), .A4(new_n338), .ZN(new_n845));
  AND4_X1   g0645(.A1(new_n365), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n365), .A2(new_n384), .A3(new_n840), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(KEYINPUT37), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n839), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT16), .B1(new_n380), .B2(new_n354), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n338), .B1(new_n850), .B2(new_n362), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n663), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n366), .B2(new_n631), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n332), .A2(new_n364), .A3(new_n851), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n843), .A2(new_n856), .A3(new_n845), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n853), .B1(new_n857), .B2(KEYINPUT100), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT100), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n843), .A2(new_n856), .A3(new_n859), .A4(new_n845), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n855), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(KEYINPUT38), .B(new_n854), .C1(new_n861), .C2(new_n846), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n849), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n838), .A2(new_n863), .A3(KEYINPUT40), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n857), .A2(KEYINPUT100), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(new_n860), .A3(new_n852), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n846), .B1(new_n867), .B2(KEYINPUT37), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n852), .B1(new_n367), .B2(new_n390), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n839), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT101), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(new_n871), .A3(new_n862), .ZN(new_n872));
  OAI211_X1 g0672(.A(KEYINPUT101), .B(new_n839), .C1(new_n868), .C2(new_n869), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(new_n838), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT40), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT103), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n874), .A2(KEYINPUT103), .A3(new_n875), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n865), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n453), .A2(new_n719), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n670), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT104), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n884), .B(new_n885), .C1(new_n881), .C2(new_n880), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n794), .B1(new_n688), .B2(new_n799), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n889), .A2(new_n872), .A3(new_n873), .A4(new_n836), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n367), .B2(new_n663), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n428), .A2(new_n665), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n872), .A2(KEYINPUT39), .A3(new_n873), .ZN(new_n894));
  XNOR2_X1  g0694(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n849), .A2(new_n862), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n893), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n690), .A2(new_n453), .A3(new_n692), .A4(new_n702), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n899), .A2(new_n633), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n898), .B(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n827), .B1(new_n887), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n901), .B2(new_n887), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n574), .B(KEYINPUT97), .Z(new_n904));
  OR2_X1    g0704(.A1(new_n904), .A2(KEYINPUT35), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(KEYINPUT35), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n228), .A2(new_n499), .A3(new_n229), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT98), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT36), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  OAI21_X1  g0712(.A(G77), .B1(new_n347), .B2(new_n348), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n913), .A2(new_n230), .B1(G50), .B2(new_n348), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(G1), .A3(new_n723), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT99), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n903), .A2(new_n911), .A3(new_n912), .A4(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT105), .ZN(G367));
  INV_X1    g0718(.A(new_n732), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n740), .B1(new_n210), .B2(new_n443), .C1(new_n919), .C2(new_n240), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n756), .A2(new_n752), .B1(new_n783), .B2(new_n436), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT110), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n746), .A2(G303), .B1(G317), .B2(new_n759), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n816), .B2(new_n748), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n305), .B1(new_n772), .B2(G311), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n764), .A2(G116), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT46), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n781), .A2(G97), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n922), .A2(new_n924), .A3(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT111), .ZN(new_n931));
  INV_X1    g0731(.A(G137), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n258), .B1(new_n763), .B2(new_n347), .C1(new_n758), .C2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(G143), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n767), .A2(new_n934), .B1(new_n202), .B2(new_n753), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n933), .B(new_n935), .C1(G150), .C2(new_n746), .ZN(new_n936));
  AOI22_X1  g0736(.A1(G50), .A2(new_n779), .B1(new_n749), .B2(G159), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n937), .A2(KEYINPUT112), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n819), .A2(G68), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(KEYINPUT112), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n936), .A2(new_n938), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n931), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT47), .Z(new_n943));
  INV_X1    g0743(.A(new_n739), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n727), .B(new_n920), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT113), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n640), .A2(new_n665), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n651), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n637), .B2(new_n949), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n947), .B(new_n948), .C1(new_n790), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n646), .A2(new_n665), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n665), .A2(new_n577), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n650), .A2(new_n635), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(new_n672), .A3(new_n678), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT106), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(KEYINPUT42), .ZN(new_n959));
  INV_X1    g0759(.A(new_n549), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n650), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n665), .B1(new_n961), .B2(new_n635), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n958), .B2(KEYINPUT42), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT107), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n964), .B2(new_n963), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n676), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n956), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT108), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n968), .A2(new_n971), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  OR3_X1    g0775(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n975), .B1(new_n972), .B2(new_n973), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n725), .A2(G1), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n679), .A2(KEYINPUT109), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT109), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n675), .B2(new_n678), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n980), .B1(new_n982), .B2(new_n679), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(new_n671), .Z(new_n984));
  NAND2_X1  g0784(.A1(new_n721), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n677), .A2(new_n679), .ZN(new_n986));
  INV_X1    g0786(.A(new_n956), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT44), .Z(new_n989));
  NOR2_X1   g0789(.A1(new_n986), .A2(new_n987), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(new_n969), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n985), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n721), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n682), .B(KEYINPUT41), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n979), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n952), .B1(new_n978), .B2(new_n998), .ZN(G387));
  OR2_X1    g0799(.A1(new_n675), .A2(new_n790), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n684), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n730), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(G107), .B2(new_n210), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n919), .B1(new_n237), .B2(G45), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n267), .B1(new_n348), .B2(new_n202), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT114), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1005), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  AND3_X1   g0807(.A1(new_n334), .A2(KEYINPUT50), .A3(new_n288), .ZN(new_n1008));
  AOI21_X1  g0808(.A(KEYINPUT50), .B1(new_n334), .B2(new_n288), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1007), .B1(new_n1006), .B2(new_n1001), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1003), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n740), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n727), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n763), .A2(new_n202), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1014), .A2(new_n357), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1015), .B(new_n928), .C1(new_n804), .C2(new_n758), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT115), .Z(new_n1017));
  NOR2_X1   g0817(.A1(new_n786), .A2(new_n443), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G50), .A2(new_n746), .B1(new_n749), .B2(new_n334), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G68), .A2(new_n779), .B1(new_n772), .B2(G159), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT116), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n305), .B1(new_n759), .B2(G326), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n783), .A2(new_n752), .B1(new_n816), .B2(new_n763), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G317), .A2(new_n746), .B1(new_n772), .B2(G322), .ZN(new_n1026));
  INV_X1    g0826(.A(G303), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1026), .B1(new_n1027), .B2(new_n756), .C1(new_n754), .C2(new_n748), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT48), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1025), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n1029), .B2(new_n1028), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT49), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1024), .B1(new_n499), .B2(new_n753), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1023), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1013), .B1(new_n1035), .B2(new_n739), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n984), .A2(new_n979), .B1(new_n1000), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n985), .A2(new_n682), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n721), .A2(new_n984), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(G393));
  OAI221_X1 g0840(.A(new_n740), .B1(new_n457), .B2(new_n210), .C1(new_n919), .C2(new_n244), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1041), .A2(new_n727), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n817), .A2(new_n774), .B1(new_n804), .B2(new_n767), .ZN(new_n1043));
  XOR2_X1   g0843(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n819), .A2(G77), .ZN(new_n1047));
  AND3_X1   g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n748), .A2(new_n288), .B1(new_n934), .B2(new_n758), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n812), .B(new_n305), .C1(new_n348), .C2(new_n763), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n334), .C2(new_n779), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G311), .A2(new_n746), .B1(new_n772), .B2(G317), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT52), .Z(new_n1053));
  OAI21_X1  g0853(.A(new_n252), .B1(new_n763), .B2(new_n752), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n759), .A2(G322), .B1(G116), .B2(new_n760), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n816), .B2(new_n756), .C1(new_n1027), .C2(new_n748), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1054), .B(new_n1056), .C1(G107), .C2(new_n781), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1048), .A2(new_n1051), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1042), .B1(new_n944), .B2(new_n1058), .C1(new_n956), .C2(new_n790), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n979), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1059), .B1(new_n993), .B2(new_n1060), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n994), .A2(new_n682), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n985), .A2(new_n993), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(G390));
  INV_X1    g0865(.A(new_n836), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n893), .B1(new_n888), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(new_n894), .A3(new_n896), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n892), .B1(new_n849), .B2(new_n862), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n798), .A2(new_n449), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n673), .B(new_n1070), .C1(new_n695), .C2(new_n701), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n794), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT118), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1071), .A2(KEYINPUT118), .A3(new_n1072), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1069), .B1(new_n1077), .B2(new_n1066), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1068), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n719), .A2(G330), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1080), .A2(new_n837), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT119), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n719), .A2(new_n670), .A3(new_n799), .A4(new_n836), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1068), .A2(new_n1078), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT119), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1079), .A2(new_n1086), .A3(new_n1081), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1083), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n894), .A2(new_n736), .A3(new_n896), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n822), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n727), .B1(new_n334), .B2(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n457), .A2(new_n756), .B1(new_n767), .B2(new_n752), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G294), .B2(new_n759), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n258), .B(new_n808), .C1(G87), .C2(new_n764), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G116), .A2(new_n746), .B1(new_n749), .B2(G107), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1047), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n817), .A2(new_n809), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G128), .B2(new_n772), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G50), .A2(new_n781), .B1(new_n759), .B2(G125), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n252), .B1(new_n749), .B2(G137), .ZN(new_n1101));
  XOR2_X1   g0901(.A(KEYINPUT54), .B(G143), .Z(new_n1102));
  NAND3_X1  g0902(.A1(new_n764), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT53), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n763), .B2(new_n804), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n779), .A2(new_n1102), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n786), .A2(new_n774), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1097), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1092), .B1(new_n1109), .B2(new_n739), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1089), .A2(new_n979), .B1(new_n1090), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(G330), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n704), .B2(new_n718), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n453), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n899), .A2(new_n633), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT120), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1071), .A2(KEYINPUT118), .A3(new_n1072), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT118), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1084), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n836), .B1(new_n1113), .B2(new_n799), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1116), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n799), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1066), .B1(new_n1080), .B2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1123), .A2(new_n1077), .A3(KEYINPUT120), .A4(new_n1084), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1066), .B1(new_n720), .B2(new_n1122), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n837), .B2(new_n1080), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n889), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1115), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1088), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1083), .A2(new_n1129), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n682), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1111), .A2(new_n1133), .ZN(G378));
  INV_X1    g0934(.A(new_n898), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n293), .A2(new_n663), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n301), .B(new_n1136), .Z(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1137), .B(new_n1138), .Z(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n880), .B2(G330), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n874), .A2(KEYINPUT103), .A3(new_n875), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT103), .B1(new_n874), .B2(new_n875), .ZN(new_n1142));
  OAI211_X1 g0942(.A(G330), .B(new_n864), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1137), .B(new_n1138), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1135), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n880), .A2(new_n1139), .A3(G330), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1147), .A2(new_n1148), .A3(new_n898), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1115), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1146), .A2(new_n1149), .B1(new_n1150), .B2(new_n1132), .ZN(new_n1151));
  OAI21_X1  g0951(.A(KEYINPUT122), .B1(new_n1151), .B2(KEYINPUT57), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n682), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n1151), .B2(KEYINPUT57), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1132), .A2(new_n1150), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1149), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n898), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT122), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1152), .A2(new_n1154), .A3(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n979), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1144), .A2(new_n736), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n727), .B1(G50), .B2(new_n1091), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n256), .A2(new_n266), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT121), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n288), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n266), .B2(new_n357), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n767), .A2(new_n499), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n756), .A2(new_n443), .B1(new_n752), .B2(new_n758), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(G107), .C2(new_n746), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1014), .A2(new_n305), .A3(G41), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n753), .A2(new_n347), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n749), .B2(G97), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1172), .A2(new_n939), .A3(new_n1173), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT58), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1169), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(G125), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n1179), .A2(new_n767), .B1(new_n756), .B2(new_n932), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G128), .B2(new_n746), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n749), .A2(G132), .B1(new_n764), .B2(new_n1102), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n804), .C2(new_n786), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1167), .B1(new_n759), .B2(G124), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(new_n774), .C2(new_n753), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1178), .B1(new_n1177), .B2(new_n1176), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1165), .B1(new_n1188), .B2(new_n739), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1164), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1163), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1162), .A2(new_n1192), .ZN(G375));
  AOI22_X1  g0993(.A1(new_n1121), .A2(new_n1124), .B1(new_n1127), .B2(new_n889), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(new_n1060), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n727), .B1(G68), .B2(new_n1091), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n817), .A2(new_n932), .B1(new_n804), .B2(new_n756), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G132), .B2(new_n772), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n819), .A2(G50), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n357), .B(new_n1174), .C1(G159), .C2(new_n764), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n749), .A2(new_n1102), .B1(new_n759), .B2(G128), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n758), .A2(new_n1027), .B1(new_n457), .B2(new_n763), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT123), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n258), .B1(new_n781), .B2(G77), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G107), .A2(new_n779), .B1(new_n749), .B2(G116), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G283), .A2(new_n746), .B1(new_n772), .B2(G294), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1019), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1202), .B1(new_n1204), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1196), .B1(new_n1209), .B2(new_n739), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n836), .B2(new_n737), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1195), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1194), .A2(new_n1115), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1130), .A2(new_n997), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1215), .ZN(G381));
  AOI21_X1  g1016(.A(new_n1159), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1155), .B(KEYINPUT57), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n682), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1191), .B1(new_n1220), .B2(new_n1161), .ZN(new_n1221));
  INV_X1    g1021(.A(G378), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1064), .A2(new_n825), .ZN(new_n1224));
  OR4_X1    g1024(.A1(G396), .A2(G387), .A3(G393), .A4(new_n1224), .ZN(new_n1225));
  OR3_X1    g1025(.A1(new_n1223), .A2(new_n1225), .A3(G381), .ZN(G407));
  OAI211_X1 g1026(.A(G407), .B(G213), .C1(G343), .C2(new_n1223), .ZN(G409));
  NAND4_X1  g1027(.A1(new_n1163), .A2(new_n1111), .A3(new_n1133), .A4(new_n1190), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1158), .A2(new_n996), .ZN(new_n1229));
  INV_X1    g1029(.A(G213), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n1228), .A2(new_n1229), .B1(new_n1230), .B2(G343), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1230), .A2(G343), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(G2897), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1194), .A2(KEYINPUT60), .A3(new_n1115), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n682), .ZN(new_n1237));
  OAI21_X1  g1037(.A(KEYINPUT60), .B1(new_n1194), .B2(new_n1115), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1237), .B1(new_n1214), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n825), .B1(new_n1239), .B2(new_n1212), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1214), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(new_n682), .A3(new_n1236), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(G384), .A3(new_n1213), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1240), .A2(KEYINPUT124), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT124), .B1(new_n1240), .B2(new_n1243), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1235), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1240), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1243), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G2897), .B(new_n1234), .C1(new_n1247), .C2(new_n1248), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1246), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT61), .B1(new_n1233), .B2(new_n1250), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1232), .B(new_n1252), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT63), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G387), .A2(new_n1064), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G390), .B(new_n952), .C1(new_n978), .C2(new_n998), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(KEYINPUT125), .A3(new_n1257), .ZN(new_n1258));
  OR3_X1    g1058(.A1(G387), .A2(KEYINPUT125), .A3(new_n1064), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(G393), .B(new_n792), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT126), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1256), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(G387), .A2(KEYINPUT126), .A3(new_n1064), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1260), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .A4(new_n1257), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1261), .A2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1231), .B1(G375), .B2(G378), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1268), .A2(KEYINPUT63), .A3(new_n1252), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1251), .A2(new_n1255), .A3(new_n1267), .A4(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1246), .A2(new_n1249), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1271), .B1(new_n1268), .B2(new_n1272), .ZN(new_n1273));
  XOR2_X1   g1073(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1274));
  NAND2_X1  g1074(.A1(new_n1253), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1268), .A2(KEYINPUT62), .A3(new_n1252), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1273), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1270), .B1(new_n1277), .B2(new_n1267), .ZN(G405));
  NAND2_X1  g1078(.A1(G375), .A2(G378), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1223), .A2(new_n1279), .A3(new_n1252), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(new_n1223), .B2(new_n1279), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1266), .B(new_n1261), .C1(new_n1281), .C2(new_n1283), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1223), .A2(new_n1279), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1267), .B(new_n1280), .C1(new_n1285), .C2(new_n1282), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(G402));
endmodule


