

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775;

  OR2_X1 U376 ( .A1(n617), .A2(n616), .ZN(n626) );
  XNOR2_X1 U377 ( .A(n497), .B(n496), .ZN(n386) );
  XNOR2_X1 U378 ( .A(n421), .B(KEYINPUT10), .ZN(n422) );
  NOR2_X2 U379 ( .A1(G953), .A2(G237), .ZN(n469) );
  NOR2_X1 U380 ( .A1(n660), .A2(n775), .ZN(n366) );
  INV_X2 U381 ( .A(G953), .ZN(n763) );
  XNOR2_X1 U382 ( .A(n577), .B(n576), .ZN(n660) );
  XNOR2_X2 U383 ( .A(n622), .B(n621), .ZN(n774) );
  NOR2_X2 U384 ( .A1(n614), .A2(n613), .ZN(n615) );
  AND2_X2 U385 ( .A1(n529), .A2(n528), .ZN(n623) );
  NOR2_X1 U386 ( .A1(n560), .A2(n600), .ZN(n541) );
  INV_X1 U387 ( .A(KEYINPUT69), .ZN(n421) );
  AND2_X1 U388 ( .A1(n369), .A2(n357), .ZN(n736) );
  NAND2_X1 U389 ( .A1(n377), .A2(n398), .ZN(n516) );
  INV_X2 U390 ( .A(n699), .ZN(n437) );
  AND2_X1 U391 ( .A1(n380), .A2(n378), .ZN(n377) );
  XNOR2_X1 U392 ( .A(n376), .B(n375), .ZN(n374) );
  XNOR2_X1 U393 ( .A(n373), .B(KEYINPUT72), .ZN(n372) );
  XNOR2_X1 U394 ( .A(KEYINPUT16), .B(G122), .ZN(n496) );
  NAND2_X1 U395 ( .A1(n404), .A2(n355), .ZN(n622) );
  NOR2_X1 U396 ( .A1(n619), .A2(n696), .ZN(n355) );
  INV_X2 U397 ( .A(n620), .ZN(n404) );
  BUF_X1 U398 ( .A(n637), .Z(n762) );
  XNOR2_X2 U399 ( .A(n439), .B(n438), .ZN(n601) );
  NOR2_X2 U400 ( .A1(n542), .A2(n589), .ZN(n439) );
  XNOR2_X2 U401 ( .A(n455), .B(n411), .ZN(n760) );
  XNOR2_X1 U402 ( .A(n367), .B(KEYINPUT20), .ZN(n434) );
  XNOR2_X1 U403 ( .A(n370), .B(KEYINPUT70), .ZN(n539) );
  NOR2_X1 U404 ( .A1(n698), .A2(n538), .ZN(n370) );
  NOR2_X1 U405 ( .A1(n736), .A2(KEYINPUT83), .ZN(n552) );
  OR2_X2 U406 ( .A1(n623), .A2(n774), .ZN(n628) );
  XNOR2_X1 U407 ( .A(n362), .B(n385), .ZN(n395) );
  INV_X1 U408 ( .A(KEYINPUT48), .ZN(n385) );
  INV_X1 U409 ( .A(n746), .ZN(n392) );
  INV_X1 U410 ( .A(n359), .ZN(n379) );
  NAND2_X1 U411 ( .A1(n511), .A2(n400), .ZN(n399) );
  INV_X1 U412 ( .A(n513), .ZN(n400) );
  OR2_X1 U413 ( .A1(n680), .A2(KEYINPUT2), .ZN(n683) );
  BUF_X1 U414 ( .A(n540), .Z(n702) );
  OR2_X1 U415 ( .A1(n407), .A2(KEYINPUT104), .ZN(n405) );
  NAND2_X1 U416 ( .A1(n620), .A2(n527), .ZN(n406) );
  INV_X1 U417 ( .A(n565), .ZN(n407) );
  XNOR2_X1 U418 ( .A(n384), .B(n383), .ZN(n433) );
  XNOR2_X1 U419 ( .A(n418), .B(KEYINPUT95), .ZN(n383) );
  OR2_X1 U420 ( .A1(n691), .A2(n534), .ZN(n536) );
  INV_X1 U421 ( .A(KEYINPUT15), .ZN(n417) );
  XNOR2_X1 U422 ( .A(G902), .B(KEYINPUT91), .ZN(n368) );
  AND2_X1 U423 ( .A1(n586), .A2(n739), .ZN(n691) );
  INV_X1 U424 ( .A(G237), .ZN(n458) );
  XNOR2_X1 U425 ( .A(n628), .B(n382), .ZN(n629) );
  INV_X1 U426 ( .A(KEYINPUT88), .ZN(n382) );
  NAND2_X1 U427 ( .A1(n763), .A2(G234), .ZN(n420) );
  NOR2_X1 U428 ( .A1(n395), .A2(n585), .ZN(n394) );
  NOR2_X1 U429 ( .A1(n393), .A2(n392), .ZN(n391) );
  XNOR2_X1 U430 ( .A(n435), .B(n371), .ZN(n698) );
  XNOR2_X1 U431 ( .A(KEYINPUT96), .B(KEYINPUT21), .ZN(n371) );
  INV_X1 U432 ( .A(G902), .ZN(n491) );
  NAND2_X1 U433 ( .A1(n434), .A2(G217), .ZN(n384) );
  XNOR2_X1 U434 ( .A(G128), .B(G119), .ZN(n424) );
  XNOR2_X1 U435 ( .A(G140), .B(KEYINPUT94), .ZN(n426) );
  XOR2_X1 U436 ( .A(KEYINPUT7), .B(G107), .Z(n486) );
  XNOR2_X1 U437 ( .A(G122), .B(G116), .ZN(n485) );
  XOR2_X1 U438 ( .A(G104), .B(G122), .Z(n475) );
  XNOR2_X1 U439 ( .A(G143), .B(G113), .ZN(n474) );
  XOR2_X1 U440 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n471) );
  XNOR2_X1 U441 ( .A(KEYINPUT92), .B(KEYINPUT17), .ZN(n502) );
  XNOR2_X1 U442 ( .A(KEYINPUT18), .B(KEYINPUT80), .ZN(n499) );
  AND2_X1 U443 ( .A1(n572), .A2(n573), .ZN(n397) );
  NOR2_X1 U444 ( .A1(n381), .A2(n379), .ZN(n378) );
  NOR2_X1 U445 ( .A1(n592), .A2(n714), .ZN(n594) );
  INV_X1 U446 ( .A(KEYINPUT34), .ZN(n593) );
  NOR2_X1 U447 ( .A1(n763), .A2(G952), .ZN(n678) );
  NOR2_X1 U448 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U449 ( .A1(n537), .A2(n542), .ZN(n369) );
  NAND2_X1 U450 ( .A1(n404), .A2(n356), .ZN(n403) );
  AND2_X1 U451 ( .A1(n407), .A2(KEYINPUT104), .ZN(n356) );
  XOR2_X1 U452 ( .A(n541), .B(n409), .Z(n357) );
  AND2_X1 U453 ( .A1(n406), .A2(n405), .ZN(n358) );
  NAND2_X1 U454 ( .A1(n512), .A2(G214), .ZN(n359) );
  AND2_X1 U455 ( .A1(n748), .A2(n585), .ZN(n360) );
  INV_X1 U456 ( .A(n402), .ZN(n381) );
  NAND2_X1 U457 ( .A1(n640), .A2(n513), .ZN(n402) );
  AND2_X1 U458 ( .A1(n361), .A2(n468), .ZN(n515) );
  NAND2_X1 U459 ( .A1(n361), .A2(n397), .ZN(n396) );
  XNOR2_X1 U460 ( .A(n601), .B(KEYINPUT106), .ZN(n361) );
  XNOR2_X2 U461 ( .A(n505), .B(G134), .ZN(n487) );
  XNOR2_X2 U462 ( .A(G143), .B(G128), .ZN(n505) );
  NAND2_X1 U463 ( .A1(n365), .A2(n363), .ZN(n362) );
  AND2_X1 U464 ( .A1(n567), .A2(n364), .ZN(n363) );
  XNOR2_X1 U465 ( .A(n744), .B(KEYINPUT87), .ZN(n364) );
  XNOR2_X1 U466 ( .A(n366), .B(KEYINPUT46), .ZN(n365) );
  NAND2_X1 U467 ( .A1(n511), .A2(G234), .ZN(n367) );
  XNOR2_X1 U468 ( .A(n368), .B(n417), .ZN(n511) );
  NAND2_X1 U469 ( .A1(n357), .A2(n543), .ZN(n569) );
  XNOR2_X2 U470 ( .A(n374), .B(n372), .ZN(n498) );
  XNOR2_X2 U471 ( .A(G113), .B(KEYINPUT3), .ZN(n373) );
  XNOR2_X2 U472 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n375) );
  XNOR2_X2 U473 ( .A(G119), .B(G116), .ZN(n376) );
  AND2_X1 U474 ( .A1(n380), .A2(n402), .ZN(n401) );
  OR2_X1 U475 ( .A1(n649), .A2(n399), .ZN(n398) );
  NAND2_X1 U476 ( .A1(n649), .A2(n513), .ZN(n380) );
  NAND2_X1 U477 ( .A1(n670), .A2(G217), .ZN(n673) );
  NAND2_X1 U478 ( .A1(n670), .A2(G478), .ZN(n677) );
  XNOR2_X2 U479 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n500) );
  AND2_X2 U480 ( .A1(n671), .A2(n491), .ZN(n432) );
  XNOR2_X2 U481 ( .A(G146), .B(G125), .ZN(n507) );
  XNOR2_X2 U482 ( .A(n507), .B(n422), .ZN(n761) );
  OR2_X2 U483 ( .A1(n532), .A2(n531), .ZN(n742) );
  XNOR2_X2 U484 ( .A(n498), .B(n386), .ZN(n754) );
  XNOR2_X2 U485 ( .A(n388), .B(n387), .ZN(n497) );
  XNOR2_X2 U486 ( .A(G110), .B(G107), .ZN(n387) );
  XNOR2_X2 U487 ( .A(G104), .B(G101), .ZN(n388) );
  NAND2_X1 U488 ( .A1(n395), .A2(n360), .ZN(n390) );
  NOR2_X2 U489 ( .A1(n394), .A2(n389), .ZN(n637) );
  NAND2_X1 U490 ( .A1(n390), .A2(n391), .ZN(n389) );
  NOR2_X1 U491 ( .A1(n748), .A2(n585), .ZN(n393) );
  INV_X1 U492 ( .A(n575), .ZN(n587) );
  XNOR2_X2 U493 ( .A(n396), .B(KEYINPUT39), .ZN(n575) );
  NAND2_X1 U494 ( .A1(n401), .A2(n398), .ZN(n583) );
  XNOR2_X1 U495 ( .A(n510), .B(n754), .ZN(n649) );
  NAND2_X1 U496 ( .A1(n404), .A2(n407), .ZN(n614) );
  NAND2_X1 U497 ( .A1(n358), .A2(n403), .ZN(n529) );
  XNOR2_X2 U498 ( .A(n408), .B(KEYINPUT22), .ZN(n620) );
  NAND2_X1 U499 ( .A1(n599), .A2(n526), .ZN(n408) );
  XOR2_X1 U500 ( .A(KEYINPUT28), .B(KEYINPUT108), .Z(n409) );
  INV_X1 U501 ( .A(KEYINPUT5), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  INV_X1 U503 ( .A(KEYINPUT8), .ZN(n419) );
  INV_X1 U504 ( .A(n476), .ZN(n411) );
  XNOR2_X1 U505 ( .A(KEYINPUT81), .B(KEYINPUT35), .ZN(n597) );
  XNOR2_X1 U506 ( .A(n457), .B(G472), .ZN(n540) );
  XNOR2_X1 U507 ( .A(n500), .B(G137), .ZN(n410) );
  XNOR2_X2 U508 ( .A(n487), .B(n410), .ZN(n455) );
  XNOR2_X1 U509 ( .A(G140), .B(G131), .ZN(n476) );
  NAND2_X1 U510 ( .A1(n763), .A2(G227), .ZN(n412) );
  XNOR2_X1 U511 ( .A(n412), .B(G146), .ZN(n413) );
  XNOR2_X1 U512 ( .A(n497), .B(n413), .ZN(n414) );
  XNOR2_X1 U513 ( .A(n760), .B(n414), .ZN(n643) );
  OR2_X2 U514 ( .A1(n643), .A2(G902), .ZN(n416) );
  XNOR2_X1 U515 ( .A(KEYINPUT71), .B(G469), .ZN(n415) );
  XNOR2_X2 U516 ( .A(n416), .B(n415), .ZN(n542) );
  XOR2_X1 U517 ( .A(KEYINPUT25), .B(KEYINPUT79), .Z(n418) );
  XNOR2_X2 U518 ( .A(n420), .B(n419), .ZN(n482) );
  NAND2_X1 U519 ( .A1(G221), .A2(n482), .ZN(n423) );
  XNOR2_X1 U520 ( .A(n423), .B(n761), .ZN(n431) );
  XOR2_X1 U521 ( .A(G137), .B(G110), .Z(n425) );
  XNOR2_X1 U522 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U523 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n427) );
  XNOR2_X1 U524 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U525 ( .A(n429), .B(n428), .Z(n430) );
  XNOR2_X1 U526 ( .A(n431), .B(n430), .ZN(n671) );
  XNOR2_X2 U527 ( .A(n433), .B(n432), .ZN(n699) );
  NAND2_X1 U528 ( .A1(n434), .A2(G221), .ZN(n435) );
  INV_X1 U529 ( .A(n698), .ZN(n436) );
  NAND2_X1 U530 ( .A1(n437), .A2(n436), .ZN(n589) );
  INV_X1 U531 ( .A(KEYINPUT97), .ZN(n438) );
  INV_X1 U532 ( .A(G101), .ZN(n440) );
  NAND2_X1 U533 ( .A1(n440), .A2(KEYINPUT76), .ZN(n443) );
  INV_X1 U534 ( .A(KEYINPUT76), .ZN(n441) );
  NAND2_X1 U535 ( .A1(G101), .A2(n441), .ZN(n442) );
  NAND2_X1 U536 ( .A1(n443), .A2(n442), .ZN(n445) );
  NAND2_X1 U537 ( .A1(n469), .A2(G210), .ZN(n444) );
  XNOR2_X1 U538 ( .A(n445), .B(n444), .ZN(n449) );
  XNOR2_X1 U539 ( .A(G146), .B(G131), .ZN(n447) );
  XNOR2_X1 U540 ( .A(n449), .B(n448), .ZN(n450) );
  NAND2_X1 U541 ( .A1(n450), .A2(n498), .ZN(n454) );
  INV_X1 U542 ( .A(n450), .ZN(n452) );
  INV_X1 U543 ( .A(n498), .ZN(n451) );
  NAND2_X1 U544 ( .A1(n452), .A2(n451), .ZN(n453) );
  NAND2_X1 U545 ( .A1(n454), .A2(n453), .ZN(n456) );
  XNOR2_X1 U546 ( .A(n456), .B(n455), .ZN(n663) );
  NAND2_X1 U547 ( .A1(n663), .A2(n491), .ZN(n457) );
  NAND2_X1 U548 ( .A1(n491), .A2(n458), .ZN(n512) );
  NAND2_X1 U549 ( .A1(n540), .A2(n359), .ZN(n460) );
  XNOR2_X1 U550 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n459) );
  XNOR2_X1 U551 ( .A(n460), .B(n459), .ZN(n573) );
  NAND2_X1 U552 ( .A1(G237), .A2(G234), .ZN(n461) );
  XNOR2_X1 U553 ( .A(n461), .B(KEYINPUT14), .ZN(n463) );
  NAND2_X1 U554 ( .A1(n463), .A2(G952), .ZN(n462) );
  XNOR2_X1 U555 ( .A(KEYINPUT93), .B(n462), .ZN(n712) );
  NAND2_X1 U556 ( .A1(n712), .A2(n763), .ZN(n522) );
  NAND2_X1 U557 ( .A1(G902), .A2(n463), .ZN(n519) );
  NOR2_X1 U558 ( .A1(G900), .A2(n519), .ZN(n464) );
  NAND2_X1 U559 ( .A1(n464), .A2(G953), .ZN(n465) );
  NAND2_X1 U560 ( .A1(n522), .A2(n465), .ZN(n467) );
  INV_X1 U561 ( .A(KEYINPUT82), .ZN(n466) );
  XNOR2_X1 U562 ( .A(n467), .B(n466), .ZN(n538) );
  INV_X1 U563 ( .A(n538), .ZN(n571) );
  AND2_X1 U564 ( .A1(n573), .A2(n571), .ZN(n468) );
  NAND2_X1 U565 ( .A1(n469), .A2(G214), .ZN(n470) );
  XNOR2_X1 U566 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U567 ( .A(KEYINPUT99), .B(n472), .ZN(n473) );
  XNOR2_X1 U568 ( .A(n473), .B(n761), .ZN(n479) );
  XNOR2_X1 U569 ( .A(n475), .B(n474), .ZN(n477) );
  XNOR2_X1 U570 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U571 ( .A(n479), .B(n478), .ZN(n655) );
  NOR2_X1 U572 ( .A1(G902), .A2(n655), .ZN(n481) );
  XNOR2_X1 U573 ( .A(KEYINPUT13), .B(G475), .ZN(n480) );
  XNOR2_X1 U574 ( .A(n481), .B(n480), .ZN(n530) );
  INV_X1 U575 ( .A(n530), .ZN(n525) );
  INV_X1 U576 ( .A(n525), .ZN(n495) );
  XOR2_X1 U577 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n484) );
  NAND2_X1 U578 ( .A1(G217), .A2(n482), .ZN(n483) );
  XNOR2_X1 U579 ( .A(n484), .B(n483), .ZN(n490) );
  XNOR2_X1 U580 ( .A(n486), .B(n485), .ZN(n488) );
  XNOR2_X1 U581 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U582 ( .A(n490), .B(n489), .ZN(n675) );
  NAND2_X1 U583 ( .A1(n675), .A2(n491), .ZN(n493) );
  INV_X1 U584 ( .A(G478), .ZN(n492) );
  XNOR2_X1 U585 ( .A(n493), .B(n492), .ZN(n531) );
  INV_X1 U586 ( .A(n531), .ZN(n494) );
  NAND2_X1 U587 ( .A1(n495), .A2(n494), .ZN(n596) );
  XNOR2_X1 U588 ( .A(n500), .B(n499), .ZN(n504) );
  NAND2_X1 U589 ( .A1(n763), .A2(G224), .ZN(n501) );
  XNOR2_X1 U590 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U591 ( .A(n504), .B(n503), .ZN(n509) );
  INV_X1 U592 ( .A(n505), .ZN(n506) );
  XNOR2_X1 U593 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U594 ( .A(n509), .B(n508), .ZN(n510) );
  INV_X1 U595 ( .A(n511), .ZN(n640) );
  NAND2_X1 U596 ( .A1(n512), .A2(G210), .ZN(n513) );
  NOR2_X1 U597 ( .A1(n596), .A2(n583), .ZN(n514) );
  AND2_X1 U598 ( .A1(n515), .A2(n514), .ZN(n554) );
  XOR2_X1 U599 ( .A(G143), .B(n554), .Z(G45) );
  XNOR2_X2 U600 ( .A(n516), .B(KEYINPUT89), .ZN(n562) );
  XNOR2_X1 U601 ( .A(KEYINPUT78), .B(KEYINPUT19), .ZN(n517) );
  XNOR2_X1 U602 ( .A(n517), .B(KEYINPUT66), .ZN(n518) );
  XNOR2_X2 U603 ( .A(n562), .B(n518), .ZN(n537) );
  INV_X1 U604 ( .A(n519), .ZN(n520) );
  NOR2_X1 U605 ( .A1(G898), .A2(n763), .ZN(n755) );
  NAND2_X1 U606 ( .A1(n520), .A2(n755), .ZN(n521) );
  AND2_X1 U607 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X2 U608 ( .A1(n537), .A2(n523), .ZN(n524) );
  XNOR2_X2 U609 ( .A(n524), .B(KEYINPUT0), .ZN(n599) );
  NAND2_X1 U610 ( .A1(n525), .A2(n531), .ZN(n688) );
  NOR2_X1 U611 ( .A1(n688), .A2(n698), .ZN(n526) );
  XNOR2_X1 U612 ( .A(n542), .B(KEYINPUT1), .ZN(n696) );
  INV_X1 U613 ( .A(n696), .ZN(n565) );
  INV_X1 U614 ( .A(KEYINPUT104), .ZN(n527) );
  NOR2_X1 U615 ( .A1(n702), .A2(n437), .ZN(n528) );
  XOR2_X1 U616 ( .A(G110), .B(n623), .Z(G12) );
  XNOR2_X1 U617 ( .A(n530), .B(KEYINPUT100), .ZN(n532) );
  XNOR2_X1 U618 ( .A(n742), .B(KEYINPUT102), .ZN(n586) );
  NAND2_X1 U619 ( .A1(n532), .A2(n531), .ZN(n739) );
  INV_X1 U620 ( .A(KEYINPUT75), .ZN(n533) );
  NAND2_X1 U621 ( .A1(n533), .A2(n545), .ZN(n534) );
  INV_X1 U622 ( .A(KEYINPUT83), .ZN(n535) );
  NAND2_X1 U623 ( .A1(n536), .A2(n535), .ZN(n544) );
  NAND2_X1 U624 ( .A1(n539), .A2(n699), .ZN(n560) );
  INV_X1 U625 ( .A(n540), .ZN(n600) );
  INV_X1 U626 ( .A(n542), .ZN(n543) );
  NAND2_X1 U627 ( .A1(n544), .A2(n736), .ZN(n547) );
  INV_X1 U628 ( .A(KEYINPUT47), .ZN(n545) );
  NAND2_X1 U629 ( .A1(n545), .A2(KEYINPUT83), .ZN(n546) );
  AND2_X1 U630 ( .A1(n547), .A2(n546), .ZN(n551) );
  NOR2_X1 U631 ( .A1(n691), .A2(KEYINPUT47), .ZN(n548) );
  NAND2_X1 U632 ( .A1(n736), .A2(n548), .ZN(n549) );
  NAND2_X1 U633 ( .A1(n549), .A2(KEYINPUT75), .ZN(n550) );
  NAND2_X1 U634 ( .A1(n551), .A2(n550), .ZN(n558) );
  NOR2_X1 U635 ( .A1(n691), .A2(n552), .ZN(n553) );
  OR2_X1 U636 ( .A1(n545), .A2(n553), .ZN(n556) );
  INV_X1 U637 ( .A(n554), .ZN(n555) );
  NAND2_X1 U638 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U639 ( .A1(n558), .A2(n557), .ZN(n567) );
  INV_X1 U640 ( .A(KEYINPUT6), .ZN(n559) );
  XNOR2_X1 U641 ( .A(n702), .B(n559), .ZN(n618) );
  NOR2_X1 U642 ( .A1(n739), .A2(n560), .ZN(n561) );
  NAND2_X1 U643 ( .A1(n618), .A2(n561), .ZN(n579) );
  INV_X1 U644 ( .A(n562), .ZN(n563) );
  NOR2_X1 U645 ( .A1(n579), .A2(n563), .ZN(n564) );
  XNOR2_X1 U646 ( .A(n564), .B(KEYINPUT36), .ZN(n566) );
  AND2_X1 U647 ( .A1(n566), .A2(n565), .ZN(n744) );
  XNOR2_X1 U648 ( .A(n583), .B(KEYINPUT38), .ZN(n686) );
  NAND2_X1 U649 ( .A1(n686), .A2(n359), .ZN(n690) );
  NOR2_X1 U650 ( .A1(n690), .A2(n688), .ZN(n568) );
  XNOR2_X1 U651 ( .A(n568), .B(KEYINPUT41), .ZN(n715) );
  NOR2_X1 U652 ( .A1(n715), .A2(n569), .ZN(n570) );
  XNOR2_X1 U653 ( .A(n570), .B(KEYINPUT42), .ZN(n775) );
  AND2_X1 U654 ( .A1(n686), .A2(n571), .ZN(n572) );
  INV_X1 U655 ( .A(n739), .ZN(n574) );
  NAND2_X1 U656 ( .A1(n575), .A2(n574), .ZN(n577) );
  INV_X1 U657 ( .A(KEYINPUT40), .ZN(n576) );
  NAND2_X1 U658 ( .A1(n696), .A2(n359), .ZN(n578) );
  NOR2_X1 U659 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U660 ( .A(KEYINPUT105), .B(n580), .Z(n582) );
  INV_X1 U661 ( .A(KEYINPUT43), .ZN(n581) );
  XNOR2_X1 U662 ( .A(n582), .B(n581), .ZN(n584) );
  NAND2_X1 U663 ( .A1(n584), .A2(n583), .ZN(n748) );
  INV_X1 U664 ( .A(KEYINPUT86), .ZN(n585) );
  OR2_X1 U665 ( .A1(n587), .A2(n586), .ZN(n746) );
  NAND2_X1 U666 ( .A1(n637), .A2(KEYINPUT2), .ZN(n588) );
  XNOR2_X1 U667 ( .A(n588), .B(KEYINPUT85), .ZN(n635) );
  INV_X1 U668 ( .A(n599), .ZN(n592) );
  BUF_X1 U669 ( .A(n589), .Z(n695) );
  NOR2_X1 U670 ( .A1(n696), .A2(n695), .ZN(n604) );
  NAND2_X1 U671 ( .A1(n604), .A2(n618), .ZN(n591) );
  INV_X1 U672 ( .A(KEYINPUT33), .ZN(n590) );
  XNOR2_X1 U673 ( .A(n591), .B(n590), .ZN(n714) );
  XNOR2_X1 U674 ( .A(n594), .B(n593), .ZN(n595) );
  NOR2_X1 U675 ( .A1(n596), .A2(n595), .ZN(n598) );
  XNOR2_X1 U676 ( .A(n598), .B(n597), .ZN(n772) );
  NAND2_X1 U677 ( .A1(n772), .A2(KEYINPUT44), .ZN(n612) );
  BUF_X1 U678 ( .A(n599), .Z(n606) );
  AND2_X1 U679 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n606), .A2(n602), .ZN(n603) );
  XNOR2_X1 U681 ( .A(n603), .B(KEYINPUT98), .ZN(n729) );
  NAND2_X1 U682 ( .A1(n604), .A2(n702), .ZN(n705) );
  INV_X1 U683 ( .A(n705), .ZN(n605) );
  NAND2_X1 U684 ( .A1(n606), .A2(n605), .ZN(n608) );
  INV_X1 U685 ( .A(KEYINPUT31), .ZN(n607) );
  XNOR2_X1 U686 ( .A(n608), .B(n607), .ZN(n741) );
  NAND2_X1 U687 ( .A1(n729), .A2(n741), .ZN(n610) );
  INV_X1 U688 ( .A(n691), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n617) );
  OR2_X1 U691 ( .A1(n618), .A2(n699), .ZN(n613) );
  XNOR2_X1 U692 ( .A(n615), .B(KEYINPUT103), .ZN(n771) );
  INV_X1 U693 ( .A(n771), .ZN(n616) );
  OR2_X1 U694 ( .A1(n618), .A2(n437), .ZN(n619) );
  INV_X1 U695 ( .A(KEYINPUT32), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n628), .A2(KEYINPUT44), .ZN(n624) );
  XNOR2_X1 U697 ( .A(n624), .B(KEYINPUT65), .ZN(n625) );
  NOR2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n632) );
  OR2_X1 U699 ( .A1(n772), .A2(KEYINPUT44), .ZN(n627) );
  XNOR2_X1 U700 ( .A(n627), .B(KEYINPUT67), .ZN(n630) );
  NAND2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n632), .A2(n631), .ZN(n634) );
  XNOR2_X1 U703 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n633) );
  XNOR2_X2 U704 ( .A(n634), .B(n633), .ZN(n680) );
  NAND2_X1 U705 ( .A1(n635), .A2(n680), .ZN(n636) );
  XNOR2_X2 U706 ( .A(n636), .B(KEYINPUT77), .ZN(n685) );
  NAND2_X1 U707 ( .A1(n680), .A2(n762), .ZN(n639) );
  INV_X1 U708 ( .A(KEYINPUT2), .ZN(n638) );
  NAND2_X1 U709 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U710 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X4 U711 ( .A1(n685), .A2(n642), .ZN(n669) );
  NAND2_X1 U712 ( .A1(n669), .A2(G469), .ZN(n646) );
  XOR2_X1 U713 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n644) );
  XNOR2_X1 U714 ( .A(n643), .B(n644), .ZN(n645) );
  XNOR2_X1 U715 ( .A(n646), .B(n645), .ZN(n647) );
  NOR2_X2 U716 ( .A1(n647), .A2(n678), .ZN(n648) );
  XNOR2_X1 U717 ( .A(n648), .B(KEYINPUT120), .ZN(G54) );
  NAND2_X1 U718 ( .A1(n669), .A2(G210), .ZN(n652) );
  XOR2_X1 U719 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n650) );
  XNOR2_X1 U720 ( .A(n649), .B(n650), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n652), .B(n651), .ZN(n653) );
  NOR2_X2 U722 ( .A1(n653), .A2(n678), .ZN(n654) );
  XNOR2_X1 U723 ( .A(n654), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U724 ( .A1(n669), .A2(G475), .ZN(n657) );
  XOR2_X1 U725 ( .A(KEYINPUT59), .B(n655), .Z(n656) );
  XNOR2_X1 U726 ( .A(n657), .B(n656), .ZN(n658) );
  NOR2_X2 U727 ( .A1(n658), .A2(n678), .ZN(n659) );
  XNOR2_X1 U728 ( .A(n659), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U729 ( .A(G131), .B(KEYINPUT127), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n660), .B(n661), .ZN(G33) );
  NAND2_X1 U731 ( .A1(n669), .A2(G472), .ZN(n665) );
  XOR2_X1 U732 ( .A(KEYINPUT90), .B(KEYINPUT62), .Z(n662) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X2 U735 ( .A1(n666), .A2(n678), .ZN(n668) );
  XNOR2_X1 U736 ( .A(KEYINPUT109), .B(KEYINPUT63), .ZN(n667) );
  XNOR2_X1 U737 ( .A(n668), .B(n667), .ZN(G57) );
  BUF_X1 U738 ( .A(n669), .Z(n670) );
  XOR2_X1 U739 ( .A(n671), .B(KEYINPUT122), .Z(n672) );
  XNOR2_X1 U740 ( .A(n673), .B(n672), .ZN(n674) );
  NOR2_X1 U741 ( .A1(n674), .A2(n678), .ZN(G66) );
  XNOR2_X1 U742 ( .A(n675), .B(KEYINPUT121), .ZN(n676) );
  XNOR2_X1 U743 ( .A(n677), .B(n676), .ZN(n679) );
  NOR2_X1 U744 ( .A1(n679), .A2(n678), .ZN(G63) );
  OR2_X1 U745 ( .A1(n762), .A2(KEYINPUT2), .ZN(n681) );
  XNOR2_X1 U746 ( .A(n681), .B(KEYINPUT84), .ZN(n682) );
  NAND2_X1 U747 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n719) );
  NOR2_X1 U749 ( .A1(n686), .A2(n359), .ZN(n687) );
  NOR2_X1 U750 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U751 ( .A(KEYINPUT117), .B(n689), .Z(n693) );
  NOR2_X1 U752 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U753 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U754 ( .A1(n714), .A2(n694), .ZN(n710) );
  NAND2_X1 U755 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U756 ( .A(n697), .B(KEYINPUT50), .ZN(n704) );
  AND2_X1 U757 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U758 ( .A(KEYINPUT49), .B(n700), .Z(n701) );
  NOR2_X1 U759 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U760 ( .A1(n704), .A2(n703), .ZN(n706) );
  NAND2_X1 U761 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U762 ( .A(KEYINPUT51), .B(n707), .ZN(n708) );
  NOR2_X1 U763 ( .A1(n708), .A2(n715), .ZN(n709) );
  NOR2_X1 U764 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U765 ( .A(KEYINPUT52), .B(n711), .Z(n713) );
  NAND2_X1 U766 ( .A1(n713), .A2(n712), .ZN(n717) );
  OR2_X1 U767 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U768 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U769 ( .A(n720), .B(KEYINPUT118), .ZN(n721) );
  NAND2_X1 U770 ( .A1(n721), .A2(n763), .ZN(n723) );
  XNOR2_X1 U771 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n722) );
  XNOR2_X1 U772 ( .A(n723), .B(n722), .ZN(G75) );
  NOR2_X1 U773 ( .A1(n729), .A2(n739), .ZN(n725) );
  XNOR2_X1 U774 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n724) );
  XNOR2_X1 U775 ( .A(n725), .B(n724), .ZN(n726) );
  XNOR2_X1 U776 ( .A(G104), .B(n726), .ZN(G6) );
  XOR2_X1 U777 ( .A(KEYINPUT112), .B(KEYINPUT26), .Z(n728) );
  XNOR2_X1 U778 ( .A(G107), .B(KEYINPUT27), .ZN(n727) );
  XNOR2_X1 U779 ( .A(n728), .B(n727), .ZN(n731) );
  NOR2_X1 U780 ( .A1(n729), .A2(n742), .ZN(n730) );
  XOR2_X1 U781 ( .A(n731), .B(n730), .Z(G9) );
  INV_X1 U782 ( .A(n736), .ZN(n732) );
  NOR2_X1 U783 ( .A1(n732), .A2(n742), .ZN(n734) );
  XNOR2_X1 U784 ( .A(KEYINPUT113), .B(KEYINPUT29), .ZN(n733) );
  XNOR2_X1 U785 ( .A(n734), .B(n733), .ZN(n735) );
  XOR2_X1 U786 ( .A(G128), .B(n735), .Z(G30) );
  NAND2_X1 U787 ( .A1(n736), .A2(n574), .ZN(n737) );
  XNOR2_X1 U788 ( .A(n737), .B(KEYINPUT114), .ZN(n738) );
  XNOR2_X1 U789 ( .A(G146), .B(n738), .ZN(G48) );
  NOR2_X1 U790 ( .A1(n739), .A2(n741), .ZN(n740) );
  XOR2_X1 U791 ( .A(G113), .B(n740), .Z(G15) );
  NOR2_X1 U792 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U793 ( .A(G116), .B(n743), .Z(G18) );
  XNOR2_X1 U794 ( .A(G125), .B(n744), .ZN(n745) );
  XNOR2_X1 U795 ( .A(n745), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U796 ( .A(G134), .B(n746), .Z(n747) );
  XNOR2_X1 U797 ( .A(n747), .B(KEYINPUT115), .ZN(G36) );
  XNOR2_X1 U798 ( .A(n748), .B(G140), .ZN(n749) );
  XNOR2_X1 U799 ( .A(KEYINPUT116), .B(n749), .ZN(G42) );
  NAND2_X1 U800 ( .A1(n680), .A2(n763), .ZN(n753) );
  NAND2_X1 U801 ( .A1(G953), .A2(G224), .ZN(n750) );
  XNOR2_X1 U802 ( .A(KEYINPUT61), .B(n750), .ZN(n751) );
  NAND2_X1 U803 ( .A1(n751), .A2(G898), .ZN(n752) );
  NAND2_X1 U804 ( .A1(n753), .A2(n752), .ZN(n758) );
  XNOR2_X1 U805 ( .A(n754), .B(KEYINPUT123), .ZN(n756) );
  NOR2_X1 U806 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U807 ( .A(n758), .B(n757), .ZN(n759) );
  XNOR2_X1 U808 ( .A(KEYINPUT124), .B(n759), .ZN(G69) );
  XOR2_X1 U809 ( .A(n761), .B(n760), .Z(n765) );
  XNOR2_X1 U810 ( .A(n762), .B(n765), .ZN(n764) );
  NAND2_X1 U811 ( .A1(n764), .A2(n763), .ZN(n770) );
  XOR2_X1 U812 ( .A(G227), .B(n765), .Z(n766) );
  NAND2_X1 U813 ( .A1(n766), .A2(G900), .ZN(n767) );
  XOR2_X1 U814 ( .A(KEYINPUT125), .B(n767), .Z(n768) );
  NAND2_X1 U815 ( .A1(G953), .A2(n768), .ZN(n769) );
  NAND2_X1 U816 ( .A1(n770), .A2(n769), .ZN(G72) );
  XNOR2_X1 U817 ( .A(n771), .B(G101), .ZN(G3) );
  XOR2_X1 U818 ( .A(G122), .B(n772), .Z(n773) );
  XNOR2_X1 U819 ( .A(KEYINPUT126), .B(n773), .ZN(G24) );
  XOR2_X1 U820 ( .A(G119), .B(n774), .Z(G21) );
  XOR2_X1 U821 ( .A(G137), .B(n775), .Z(G39) );
endmodule

