//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G137), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(G137), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT11), .A3(G134), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n193), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G131), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT67), .B(G131), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n198), .A2(new_n192), .A3(new_n193), .A4(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n204), .A3(G146), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n201), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n205), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT65), .B(G143), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n206), .B1(new_n211), .B2(G146), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(G146), .B1(new_n202), .B2(new_n204), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n215));
  OAI21_X1  g029(.A(G128), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n210), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT76), .B1(new_n218), .B2(G107), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(G107), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n218), .A2(KEYINPUT76), .A3(G107), .ZN(new_n222));
  OAI21_X1  g036(.A(G101), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT3), .B1(new_n218), .B2(G107), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n225));
  INV_X1    g039(.A(G107), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G104), .ZN(new_n227));
  INV_X1    g041(.A(G101), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n224), .A2(new_n227), .A3(new_n228), .A4(new_n220), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n217), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n230), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n205), .A2(new_n207), .A3(new_n209), .ZN(new_n233));
  INV_X1    g047(.A(G146), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n202), .A2(new_n204), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(new_n234), .ZN(new_n237));
  OAI21_X1  g051(.A(G128), .B1(new_n206), .B2(new_n215), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n233), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n232), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n200), .B1(new_n231), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT12), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(G110), .B(G140), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(KEYINPUT75), .ZN(new_n246));
  INV_X1    g060(.A(G953), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n247), .A2(G227), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n246), .B(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n235), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n211), .B2(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT0), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(new_n208), .A3(KEYINPUT64), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT64), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n256), .B1(KEYINPUT0), .B2(G128), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n253), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n259), .A2(KEYINPUT66), .B1(new_n253), .B2(new_n212), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n251), .A2(new_n261), .A3(new_n258), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n224), .A2(new_n227), .A3(new_n220), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(G101), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(G101), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT4), .A3(new_n229), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n260), .A2(new_n262), .A3(new_n265), .A4(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT10), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n269), .B1(new_n217), .B2(new_n230), .ZN(new_n270));
  INV_X1    g084(.A(new_n200), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n251), .A2(new_n238), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n269), .B1(new_n272), .B2(new_n233), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n232), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n268), .A2(new_n270), .A3(new_n271), .A4(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT77), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n255), .A2(new_n257), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n252), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT66), .B1(new_n237), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n212), .A2(new_n253), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n280), .A2(new_n262), .A3(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n267), .A2(new_n265), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n282), .A2(new_n283), .B1(new_n232), .B2(new_n273), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n284), .A2(KEYINPUT77), .A3(new_n271), .A4(new_n270), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n249), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT78), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n244), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI211_X1 g102(.A(KEYINPUT78), .B(new_n249), .C1(new_n277), .C2(new_n285), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n277), .A2(new_n285), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n284), .A2(new_n270), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n200), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n249), .ZN(new_n294));
  OAI22_X1  g108(.A1(new_n288), .A2(new_n289), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G469), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n244), .A2(new_n290), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n299), .A2(new_n249), .B1(new_n292), .B2(new_n286), .ZN(new_n300));
  OAI21_X1  g114(.A(G469), .B1(new_n300), .B2(G902), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n189), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT79), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G234), .ZN(new_n305));
  OAI21_X1  g119(.A(G217), .B1(new_n305), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n307));
  INV_X1    g121(.A(G140), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G125), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n307), .B1(new_n309), .B2(KEYINPUT16), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT16), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n311), .A2(new_n308), .A3(KEYINPUT74), .A4(G125), .ZN(new_n312));
  INV_X1    g126(.A(G125), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n310), .B(new_n312), .C1(new_n315), .C2(new_n311), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(new_n234), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n208), .A2(G119), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n208), .A2(G119), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G110), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n318), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT24), .B(G110), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n317), .B(new_n325), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n327), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n324), .B2(G110), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n316), .A2(new_n234), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n330), .B(new_n331), .C1(G146), .C2(new_n315), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n247), .A2(G221), .A3(G234), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(KEYINPUT22), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(G137), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n328), .A2(new_n332), .A3(new_n336), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n297), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n306), .B1(new_n340), .B2(KEYINPUT25), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(KEYINPUT25), .B2(new_n340), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n338), .A2(new_n339), .ZN(new_n343));
  AOI21_X1  g157(.A(G902), .B1(new_n305), .B2(G217), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n280), .A2(new_n262), .A3(new_n281), .A4(new_n200), .ZN(new_n347));
  INV_X1    g161(.A(new_n193), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n191), .A2(G137), .ZN(new_n349));
  OAI21_X1  g163(.A(G131), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n199), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n240), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT2), .B(G113), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(G116), .B(G119), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XOR2_X1   g171(.A(G116), .B(G119), .Z(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n354), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n353), .A2(KEYINPUT71), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n360), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT68), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n240), .A2(new_n351), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n363), .B1(new_n240), .B2(new_n351), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n362), .B(new_n347), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT71), .B1(new_n353), .B2(new_n360), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT28), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n347), .A2(new_n362), .A3(new_n352), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT28), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(KEYINPUT69), .A2(G237), .ZN(new_n374));
  NOR2_X1   g188(.A1(KEYINPUT69), .A2(G237), .ZN(new_n375));
  OAI211_X1 g189(.A(G210), .B(new_n247), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT27), .ZN(new_n377));
  OR2_X1    g191(.A1(KEYINPUT69), .A2(G237), .ZN(new_n378));
  NAND2_X1  g192(.A1(KEYINPUT69), .A2(G237), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT27), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G210), .A4(new_n247), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT26), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n377), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n383), .B1(new_n377), .B2(new_n382), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n228), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n377), .A2(new_n382), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT26), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n377), .A2(new_n382), .A3(new_n383), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(G101), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n373), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT30), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n251), .A2(new_n238), .B1(new_n212), .B2(new_n209), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n199), .A2(new_n350), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT68), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n240), .A2(new_n351), .A3(new_n363), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n394), .B1(new_n399), .B2(new_n347), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n347), .A2(new_n394), .A3(new_n352), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n360), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT70), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n366), .A2(new_n391), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n366), .A2(new_n391), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT70), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT31), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT31), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n403), .A2(new_n407), .A3(new_n410), .A4(new_n405), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n393), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(G472), .A2(G902), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n412), .A2(KEYINPUT32), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT32), .B1(new_n412), .B2(new_n413), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n347), .B1(new_n364), .B2(new_n365), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT30), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n362), .B1(new_n418), .B2(new_n401), .ZN(new_n419));
  INV_X1    g233(.A(new_n366), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n392), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT72), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT72), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n424), .B(new_n392), .C1(new_n419), .C2(new_n420), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n369), .A2(new_n372), .A3(new_n391), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n422), .A2(new_n423), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n417), .A2(new_n360), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n371), .B1(new_n428), .B2(new_n366), .ZN(new_n429));
  INV_X1    g243(.A(new_n372), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n392), .A2(new_n423), .ZN(new_n432));
  AOI21_X1  g246(.A(G902), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G472), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n346), .B1(new_n416), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G113), .B(G122), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(new_n218), .ZN(new_n438));
  AOI21_X1  g252(.A(G953), .B1(new_n378), .B2(new_n379), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G214), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(KEYINPUT84), .B2(new_n236), .ZN(new_n441));
  AOI21_X1  g255(.A(G143), .B1(new_n203), .B2(KEYINPUT84), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(G214), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(KEYINPUT18), .A2(G131), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n315), .B(G146), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n441), .A2(KEYINPUT18), .A3(G131), .A4(new_n443), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n317), .A2(KEYINPUT86), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n316), .A2(new_n234), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n331), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n198), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n441), .A2(KEYINPUT17), .A3(new_n454), .A4(new_n443), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n450), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n441), .A2(new_n454), .A3(new_n443), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n454), .B1(new_n441), .B2(new_n443), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT17), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n438), .B(new_n449), .C1(new_n456), .C2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n438), .ZN(new_n462));
  INV_X1    g276(.A(new_n449), .ZN(new_n463));
  INV_X1    g277(.A(new_n315), .ZN(new_n464));
  AND2_X1   g278(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n465));
  NOR2_X1   g279(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n467), .B(new_n234), .C1(new_n464), .C2(new_n466), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n331), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n459), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(new_n457), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n462), .B1(new_n463), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n461), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(G475), .A2(G902), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT20), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT20), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n477), .A3(new_n474), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n449), .B1(new_n456), .B2(new_n460), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n462), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n461), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n297), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n476), .A2(new_n478), .B1(new_n482), .B2(G475), .ZN(new_n483));
  INV_X1    g297(.A(new_n187), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(G217), .A3(new_n247), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT87), .ZN(new_n487));
  INV_X1    g301(.A(G122), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n487), .B1(new_n488), .B2(G116), .ZN(new_n489));
  INV_X1    g303(.A(G116), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(KEYINPUT87), .A3(G122), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n490), .A2(G122), .ZN(new_n493));
  OAI21_X1  g307(.A(G107), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n489), .A2(new_n491), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n495), .B(new_n226), .C1(new_n490), .C2(G122), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n211), .A2(G128), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n208), .A2(G143), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n191), .A3(new_n499), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n498), .A2(KEYINPUT13), .A3(new_n499), .ZN(new_n501));
  OAI21_X1  g315(.A(G134), .B1(new_n498), .B2(KEYINPUT13), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n497), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT14), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n493), .B1(new_n492), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n495), .A2(KEYINPUT14), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n226), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n500), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n191), .B1(new_n498), .B2(new_n499), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n496), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n503), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(KEYINPUT88), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT88), .ZN(new_n513));
  INV_X1    g327(.A(new_n507), .ZN(new_n514));
  INV_X1    g328(.A(new_n509), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n500), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n496), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n513), .B1(new_n517), .B2(new_n503), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n486), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n503), .A3(new_n513), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n485), .ZN(new_n521));
  AOI21_X1  g335(.A(G902), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G478), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(KEYINPUT15), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n511), .A2(KEYINPUT88), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n485), .B1(new_n527), .B2(new_n520), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n512), .A2(new_n486), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n297), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n524), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n483), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n247), .A2(G952), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n534), .B1(G234), .B2(G237), .ZN(new_n535));
  AOI211_X1 g349(.A(new_n297), .B(new_n247), .C1(G234), .C2(G237), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT21), .B(G898), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n533), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G214), .B1(G237), .B2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G210), .B1(G237), .B2(G902), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n490), .A2(KEYINPUT5), .A3(G119), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT81), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT5), .ZN(new_n545));
  OAI21_X1  g359(.A(G113), .B1(new_n358), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n357), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n547), .A2(new_n230), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT82), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n547), .A2(new_n549), .A3(new_n230), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n547), .B2(new_n230), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G110), .B(G122), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n283), .A2(KEYINPUT80), .A3(new_n360), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n267), .A2(new_n360), .A3(new_n265), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT80), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n556), .A2(new_n553), .A3(new_n548), .A4(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n240), .A2(G125), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n280), .A2(new_n262), .A3(new_n281), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n562), .B1(new_n563), .B2(G125), .ZN(new_n564));
  INV_X1    g378(.A(G224), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(G953), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT7), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n566), .A2(KEYINPUT83), .ZN(new_n569));
  OR3_X1    g383(.A1(new_n564), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n568), .B1(new_n564), .B2(new_n569), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(G902), .B1(new_n561), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n556), .A2(new_n548), .A3(new_n559), .ZN(new_n574));
  INV_X1    g388(.A(new_n553), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n560), .A3(KEYINPUT6), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n564), .B(new_n567), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT6), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n574), .A2(new_n579), .A3(new_n575), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n542), .B1(new_n573), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n573), .A2(new_n581), .A3(new_n542), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n541), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n304), .A2(new_n436), .A3(new_n539), .A4(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT89), .B(G101), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(G3));
  NAND2_X1  g402(.A1(new_n412), .A2(new_n297), .ZN(new_n589));
  INV_X1    g403(.A(G472), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(KEYINPUT90), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n591), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n412), .B2(new_n297), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n592), .A2(new_n346), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n304), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT92), .B1(new_n522), .B2(G478), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT92), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n530), .A2(new_n599), .A3(new_n523), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n519), .A2(new_n602), .A3(new_n521), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n486), .A2(KEYINPUT91), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n511), .B(new_n604), .Z(new_n605));
  OAI21_X1  g419(.A(new_n603), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n523), .A2(G902), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n477), .B1(new_n473), .B2(new_n474), .ZN(new_n610));
  INV_X1    g424(.A(new_n474), .ZN(new_n611));
  AOI211_X1 g425(.A(KEYINPUT20), .B(new_n611), .C1(new_n461), .C2(new_n472), .ZN(new_n612));
  AOI21_X1  g426(.A(G902), .B1(new_n480), .B2(new_n461), .ZN(new_n613));
  INV_X1    g427(.A(G475), .ZN(new_n614));
  OAI22_X1  g428(.A1(new_n610), .A2(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n538), .ZN(new_n617));
  INV_X1    g431(.A(new_n584), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n617), .B(new_n540), .C1(new_n618), .C2(new_n582), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n597), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NAND2_X1  g437(.A1(new_n526), .A2(new_n531), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n483), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n597), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT93), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT35), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G107), .ZN(G9));
  NOR2_X1   g444(.A1(new_n592), .A2(new_n594), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n333), .B(KEYINPUT94), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n337), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n344), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n342), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n304), .A2(new_n638), .A3(new_n539), .A4(new_n585), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  INV_X1    g455(.A(G900), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n536), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n535), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n625), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n636), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n416), .B2(new_n435), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n304), .A2(new_n585), .A3(new_n647), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT95), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  XNOR2_X1  g466(.A(new_n645), .B(KEYINPUT39), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n304), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT97), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n658));
  OR3_X1    g472(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT98), .ZN(new_n659));
  OAI21_X1  g473(.A(KEYINPUT98), .B1(new_n657), .B2(new_n658), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n618), .A2(new_n582), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT96), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n662), .B(KEYINPUT38), .Z(new_n663));
  NAND2_X1  g477(.A1(new_n428), .A2(new_n366), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n392), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n408), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n666), .B2(G902), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n416), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n648), .A2(new_n624), .A3(new_n615), .A4(new_n540), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n663), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n659), .A2(new_n660), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n236), .ZN(G45));
  AOI22_X1  g486(.A1(new_n598), .A2(new_n600), .B1(new_n606), .B2(new_n607), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n483), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n645), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n304), .A2(new_n585), .A3(new_n649), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  AOI21_X1  g492(.A(new_n294), .B1(new_n290), .B2(new_n292), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n242), .B(KEYINPUT12), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n275), .A2(new_n276), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n275), .A2(new_n276), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n294), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n680), .B1(new_n683), .B2(KEYINPUT78), .ZN(new_n684));
  INV_X1    g498(.A(new_n289), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n679), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(G469), .B1(new_n686), .B2(G902), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n188), .A3(new_n298), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT99), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n687), .A2(KEYINPUT99), .A3(new_n188), .A4(new_n298), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n436), .A2(new_n620), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND4_X1  g508(.A1(new_n436), .A2(new_n626), .A3(new_n690), .A4(new_n691), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  INV_X1    g510(.A(new_n585), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n688), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n649), .A2(new_n698), .A3(new_n539), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  INV_X1    g514(.A(KEYINPUT100), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n615), .A2(new_n624), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n701), .B1(new_n615), .B2(new_n624), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n619), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n589), .A2(G472), .ZN(new_n705));
  INV_X1    g519(.A(new_n346), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n409), .B(new_n411), .C1(new_n391), .C2(new_n431), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n413), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n690), .A2(new_n704), .A3(new_n710), .A4(new_n691), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT101), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT100), .B1(new_n483), .B2(new_n532), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n615), .A2(new_n624), .A3(new_n701), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n585), .A3(new_n617), .A4(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n709), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(KEYINPUT101), .A3(new_n690), .A4(new_n691), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G122), .ZN(G24));
  AND2_X1   g534(.A1(new_n705), .A2(new_n708), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n721), .A2(new_n636), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n676), .A3(new_n698), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n298), .A2(new_n725), .A3(new_n301), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n725), .B1(new_n298), .B2(new_n301), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n188), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT103), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n412), .A2(new_n413), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT32), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n412), .A2(KEYINPUT32), .A3(new_n413), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n435), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n661), .A2(new_n540), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n735), .A2(new_n737), .A3(new_n706), .ZN(new_n738));
  OAI211_X1 g552(.A(KEYINPUT103), .B(new_n188), .C1(new_n726), .C2(new_n727), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n730), .A2(new_n738), .A3(new_n676), .A4(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT42), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  XNOR2_X1  g557(.A(new_n647), .B(KEYINPUT104), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n730), .A2(new_n744), .A3(new_n739), .A4(new_n738), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT105), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  NAND2_X1  g561(.A1(new_n609), .A2(new_n483), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT43), .B1(new_n483), .B2(KEYINPUT106), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n631), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n751), .A3(new_n636), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n736), .B1(new_n753), .B2(KEYINPUT44), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n300), .A2(KEYINPUT45), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n300), .A2(KEYINPUT45), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(G469), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(G469), .A2(G902), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT46), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n298), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n757), .A2(KEYINPUT46), .A3(new_n758), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n189), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n763), .A2(new_n653), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n754), .B(new_n764), .C1(KEYINPUT44), .C2(new_n753), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G137), .ZN(G39));
  XNOR2_X1  g580(.A(new_n763), .B(KEYINPUT47), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n675), .A2(new_n736), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n735), .A2(new_n706), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n772));
  INV_X1    g586(.A(new_n688), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n663), .A2(new_n541), .A3(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n750), .A2(new_n535), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n710), .ZN(new_n776));
  OR4_X1    g590(.A1(new_n772), .A2(new_n774), .A3(KEYINPUT50), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n688), .A2(new_n736), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n668), .A2(new_n778), .A3(new_n706), .A4(new_n535), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT114), .Z(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n483), .A3(new_n673), .ZN(new_n781));
  XNOR2_X1  g595(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(new_n774), .B2(new_n776), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n775), .A2(new_n722), .A3(new_n778), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n777), .A2(new_n781), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n767), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n687), .A2(new_n189), .A3(new_n298), .ZN(new_n787));
  AOI211_X1 g601(.A(new_n736), .B(new_n776), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n789), .A2(KEYINPUT51), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(KEYINPUT51), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n775), .A2(new_n436), .A3(new_n778), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT48), .Z(new_n793));
  NOR3_X1   g607(.A1(new_n776), .A2(new_n697), .A3(new_n688), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n794), .A2(KEYINPUT116), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(KEYINPUT116), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n534), .B(KEYINPUT115), .Z(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI211_X1 g612(.A(new_n793), .B(new_n798), .C1(new_n674), .C2(new_n780), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n790), .A2(new_n791), .A3(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n692), .A2(new_n695), .A3(new_n699), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n719), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n730), .A2(new_n721), .A3(new_n739), .A4(new_n768), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n736), .A2(new_n533), .A3(new_n646), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n304), .A2(new_n735), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n648), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n619), .B1(new_n616), .B2(new_n625), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n298), .A2(new_n301), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n303), .B1(new_n809), .B2(new_n188), .ZN(new_n810));
  AOI211_X1 g624(.A(KEYINPUT79), .B(new_n189), .C1(new_n298), .C2(new_n301), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n808), .B(new_n595), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n539), .B(new_n585), .C1(new_n810), .C2(new_n811), .ZN(new_n813));
  INV_X1    g627(.A(new_n436), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n813), .A2(new_n637), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT107), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT107), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n586), .A2(new_n639), .A3(new_n818), .A4(new_n812), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n807), .A2(new_n742), .A3(new_n746), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n636), .A2(new_n646), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n188), .B(new_n822), .C1(new_n726), .C2(new_n727), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT108), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n809), .A2(KEYINPUT102), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n298), .A2(new_n725), .A3(new_n301), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(KEYINPUT108), .A3(new_n188), .A4(new_n822), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n702), .A2(new_n703), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n585), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n668), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n825), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n650), .A3(new_n677), .A4(new_n723), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT109), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT109), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT52), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n834), .A2(KEYINPUT110), .A3(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n834), .A2(KEYINPUT110), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n837), .A3(KEYINPUT52), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n821), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n834), .B(KEYINPUT52), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n844), .B1(new_n821), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n843), .A2(KEYINPUT53), .B1(new_n846), .B2(KEYINPUT111), .ZN(new_n847));
  XOR2_X1   g661(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n848));
  INV_X1    g662(.A(KEYINPUT111), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n849), .B(new_n844), .C1(new_n821), .C2(new_n845), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  OR3_X1    g665(.A1(new_n821), .A2(new_n845), .A3(new_n844), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(KEYINPUT53), .B2(new_n843), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n800), .A2(new_n855), .B1(G952), .B2(G953), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n687), .A2(new_n298), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n857), .A2(KEYINPUT49), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(KEYINPUT49), .ZN(new_n859));
  INV_X1    g673(.A(new_n668), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n706), .A2(new_n188), .A3(new_n540), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n860), .A2(new_n748), .A3(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n663), .A2(new_n858), .A3(new_n859), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n856), .A2(new_n863), .ZN(G75));
  NOR2_X1   g678(.A1(new_n247), .A2(G952), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n577), .A2(new_n580), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(new_n578), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT55), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n846), .A2(KEYINPUT111), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n842), .A2(new_n836), .A3(new_n839), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n807), .A2(new_n742), .A3(new_n746), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT53), .A4(new_n820), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n869), .A2(new_n850), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(G210), .A3(G902), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT56), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n868), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n874), .B(KEYINPUT117), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n868), .A2(new_n875), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n865), .B(new_n876), .C1(new_n877), .C2(new_n878), .ZN(G51));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n873), .A2(G902), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(new_n757), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n758), .B(KEYINPUT57), .Z(new_n883));
  AOI21_X1  g697(.A(new_n848), .B1(new_n847), .B2(new_n850), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n848), .A2(new_n869), .A3(new_n850), .A4(new_n872), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n686), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n883), .ZN(new_n889));
  INV_X1    g703(.A(new_n848), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n873), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n889), .B1(new_n851), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT118), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n882), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n880), .B1(new_n894), .B2(new_n865), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n295), .B1(new_n892), .B2(KEYINPUT118), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n886), .A2(new_n887), .ZN(new_n897));
  OAI22_X1  g711(.A1(new_n896), .A2(new_n897), .B1(new_n757), .B2(new_n881), .ZN(new_n898));
  INV_X1    g712(.A(new_n865), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(KEYINPUT119), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n895), .A2(new_n900), .ZN(G54));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n881), .A2(new_n902), .A3(new_n614), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n899), .B1(new_n903), .B2(new_n473), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n473), .B2(new_n903), .ZN(G60));
  NAND2_X1  g719(.A1(G478), .A2(G902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT59), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n606), .B1(new_n855), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n606), .A2(new_n907), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n851), .B2(new_n891), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n908), .A2(new_n865), .A3(new_n910), .ZN(G63));
  NAND2_X1  g725(.A1(G217), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT60), .Z(new_n913));
  NAND3_X1  g727(.A1(new_n873), .A2(new_n634), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT120), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n343), .B1(new_n873), .B2(new_n913), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(new_n865), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g733(.A(G953), .B1(new_n537), .B2(new_n565), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT121), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n802), .B1(new_n819), .B2(new_n817), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(G953), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n866), .B1(G898), .B2(new_n247), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT122), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n923), .B(new_n925), .ZN(G69));
  NAND2_X1  g740(.A1(new_n418), .A2(new_n401), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT123), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n467), .B1(new_n464), .B2(new_n466), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n928), .B(new_n929), .Z(new_n930));
  NAND3_X1  g744(.A1(new_n650), .A2(new_n677), .A3(new_n723), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT124), .Z(new_n932));
  NAND2_X1  g746(.A1(new_n671), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n933), .A2(KEYINPUT62), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n770), .A2(new_n765), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n616), .A2(new_n625), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n656), .A2(new_n738), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n933), .B2(KEYINPUT62), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n930), .B1(new_n940), .B2(new_n247), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT125), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n764), .A2(new_n436), .A3(new_n585), .A4(new_n830), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n935), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(new_n742), .A3(new_n746), .A4(new_n932), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n247), .A3(new_n948), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n949), .B(new_n930), .C1(new_n642), .C2(new_n247), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n951));
  AOI21_X1  g765(.A(G953), .B1(new_n934), .B2(new_n939), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(new_n930), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n942), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n247), .B1(G227), .B2(G900), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n955), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n942), .A2(new_n957), .A3(new_n950), .A4(new_n953), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(G72));
  NOR2_X1   g773(.A1(new_n419), .A2(new_n420), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n392), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n947), .A2(new_n922), .A3(new_n948), .ZN(new_n962));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  NAND2_X1  g778(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n962), .A2(KEYINPUT127), .A3(new_n964), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n961), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n934), .A2(new_n922), .A3(new_n939), .ZN(new_n970));
  AOI211_X1 g784(.A(new_n392), .B(new_n960), .C1(new_n970), .C2(new_n964), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n422), .A2(new_n425), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n408), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n853), .A2(new_n964), .A3(new_n973), .ZN(new_n974));
  NOR4_X1   g788(.A1(new_n969), .A2(new_n865), .A3(new_n971), .A4(new_n974), .ZN(G57));
endmodule


