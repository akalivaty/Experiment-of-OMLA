

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(n749), .A2(n751), .ZN(n694) );
  NOR2_X1 U553 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U554 ( .A(n690), .B(KEYINPUT64), .ZN(n710) );
  NOR2_X1 U555 ( .A1(n790), .A2(n791), .ZN(n690) );
  BUF_X2 U556 ( .A(n896), .Z(n518) );
  NOR2_X1 U557 ( .A1(G2105), .A2(n525), .ZN(n896) );
  BUF_X2 U558 ( .A(n895), .Z(n519) );
  XNOR2_X1 U559 ( .A(n521), .B(KEYINPUT17), .ZN(n895) );
  INV_X1 U560 ( .A(G2105), .ZN(n520) );
  INV_X1 U561 ( .A(KEYINPUT95), .ZN(n734) );
  INV_X1 U562 ( .A(KEYINPUT99), .ZN(n745) );
  XNOR2_X1 U563 ( .A(n748), .B(KEYINPUT32), .ZN(n775) );
  INV_X1 U564 ( .A(n790), .ZN(n792) );
  NAND2_X1 U565 ( .A1(n520), .A2(n525), .ZN(n521) );
  AND2_X2 U566 ( .A1(n525), .A2(G2105), .ZN(n891) );
  NAND2_X1 U567 ( .A1(n519), .A2(G137), .ZN(n524) );
  INV_X1 U568 ( .A(G2104), .ZN(n525) );
  NAND2_X1 U569 ( .A1(G101), .A2(n518), .ZN(n522) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(n522), .Z(n523) );
  NAND2_X1 U571 ( .A1(n524), .A2(n523), .ZN(n529) );
  NAND2_X1 U572 ( .A1(G125), .A2(n891), .ZN(n527) );
  AND2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n892) );
  NAND2_X1 U574 ( .A1(G113), .A2(n892), .ZN(n526) );
  NAND2_X1 U575 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X2 U576 ( .A1(n529), .A2(n528), .ZN(G160) );
  NOR2_X2 U577 ( .A1(G543), .A2(G651), .ZN(n650) );
  NAND2_X1 U578 ( .A1(n650), .A2(G89), .ZN(n530) );
  XNOR2_X1 U579 ( .A(n530), .B(KEYINPUT4), .ZN(n532) );
  XOR2_X1 U580 ( .A(KEYINPUT0), .B(G543), .Z(n638) );
  INV_X1 U581 ( .A(G651), .ZN(n534) );
  NOR2_X1 U582 ( .A1(n638), .A2(n534), .ZN(n578) );
  BUF_X1 U583 ( .A(n578), .Z(n651) );
  NAND2_X1 U584 ( .A1(G76), .A2(n651), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U586 ( .A(n533), .B(KEYINPUT5), .ZN(n541) );
  NOR2_X1 U587 ( .A1(G543), .A2(n534), .ZN(n535) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n535), .Z(n576) );
  BUF_X1 U589 ( .A(n576), .Z(n649) );
  NAND2_X1 U590 ( .A1(G63), .A2(n649), .ZN(n538) );
  NOR2_X1 U591 ( .A1(n638), .A2(G651), .ZN(n536) );
  XNOR2_X1 U592 ( .A(KEYINPUT66), .B(n536), .ZN(n656) );
  NAND2_X1 U593 ( .A1(G51), .A2(n656), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U595 ( .A(KEYINPUT6), .B(n539), .Z(n540) );
  NAND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U597 ( .A(n542), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U598 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U599 ( .A(G2446), .B(G2451), .Z(n544) );
  XNOR2_X1 U600 ( .A(G2454), .B(KEYINPUT103), .ZN(n543) );
  XNOR2_X1 U601 ( .A(n544), .B(n543), .ZN(n551) );
  XOR2_X1 U602 ( .A(G2438), .B(G2430), .Z(n546) );
  XNOR2_X1 U603 ( .A(G2435), .B(G2443), .ZN(n545) );
  XNOR2_X1 U604 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U605 ( .A(n547), .B(G2427), .Z(n549) );
  XNOR2_X1 U606 ( .A(G1348), .B(G1341), .ZN(n548) );
  XNOR2_X1 U607 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U608 ( .A(n551), .B(n550), .ZN(n552) );
  AND2_X1 U609 ( .A1(n552), .A2(G14), .ZN(G401) );
  NAND2_X1 U610 ( .A1(G64), .A2(n649), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G52), .A2(n656), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n559) );
  NAND2_X1 U613 ( .A1(G90), .A2(n650), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G77), .A2(n651), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U616 ( .A(KEYINPUT9), .B(n557), .Z(n558) );
  NOR2_X1 U617 ( .A1(n559), .A2(n558), .ZN(G171) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G82), .ZN(G220) );
  INV_X1 U621 ( .A(G120), .ZN(G236) );
  INV_X1 U622 ( .A(G69), .ZN(G235) );
  INV_X1 U623 ( .A(G108), .ZN(G238) );
  AND2_X1 U624 ( .A1(n519), .A2(G138), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G102), .A2(n518), .ZN(n561) );
  NAND2_X1 U626 ( .A1(G114), .A2(n892), .ZN(n560) );
  AND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n891), .A2(G126), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT84), .ZN(n563) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n688) );
  BUF_X1 U632 ( .A(n688), .Z(G164) );
  NAND2_X1 U633 ( .A1(G62), .A2(n649), .ZN(n568) );
  NAND2_X1 U634 ( .A1(G50), .A2(n656), .ZN(n567) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U636 ( .A(KEYINPUT78), .B(n569), .Z(n573) );
  NAND2_X1 U637 ( .A1(G88), .A2(n650), .ZN(n571) );
  NAND2_X1 U638 ( .A1(G75), .A2(n651), .ZN(n570) );
  AND2_X1 U639 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(G303) );
  NAND2_X1 U641 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U643 ( .A(G223), .ZN(n841) );
  NAND2_X1 U644 ( .A1(n841), .A2(G567), .ZN(n575) );
  XOR2_X1 U645 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  INV_X1 U646 ( .A(G860), .ZN(n609) );
  NAND2_X1 U647 ( .A1(n576), .A2(G56), .ZN(n577) );
  XNOR2_X1 U648 ( .A(KEYINPUT14), .B(n577), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n578), .A2(G68), .ZN(n579) );
  XNOR2_X1 U650 ( .A(KEYINPUT68), .B(n579), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n650), .A2(G81), .ZN(n580) );
  XNOR2_X1 U652 ( .A(KEYINPUT12), .B(n580), .ZN(n581) );
  NAND2_X1 U653 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U654 ( .A(KEYINPUT13), .B(n583), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U656 ( .A(n586), .B(KEYINPUT69), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G43), .A2(n656), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U659 ( .A(KEYINPUT70), .B(n589), .ZN(n967) );
  OR2_X1 U660 ( .A1(n609), .A2(n967), .ZN(G153) );
  INV_X1 U661 ( .A(G868), .ZN(n669) );
  NOR2_X1 U662 ( .A1(n669), .A2(G171), .ZN(n590) );
  XNOR2_X1 U663 ( .A(n590), .B(KEYINPUT71), .ZN(n599) );
  NAND2_X1 U664 ( .A1(G66), .A2(n649), .ZN(n592) );
  NAND2_X1 U665 ( .A1(G92), .A2(n650), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U667 ( .A1(G79), .A2(n651), .ZN(n594) );
  NAND2_X1 U668 ( .A1(G54), .A2(n656), .ZN(n593) );
  NAND2_X1 U669 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U671 ( .A(KEYINPUT15), .B(n597), .Z(n945) );
  OR2_X1 U672 ( .A1(G868), .A2(n945), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U674 ( .A1(G65), .A2(n649), .ZN(n601) );
  NAND2_X1 U675 ( .A1(G53), .A2(n656), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U677 ( .A1(G91), .A2(n650), .ZN(n603) );
  NAND2_X1 U678 ( .A1(G78), .A2(n651), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n948) );
  XNOR2_X1 U681 ( .A(n948), .B(KEYINPUT67), .ZN(G299) );
  XNOR2_X1 U682 ( .A(KEYINPUT72), .B(n669), .ZN(n606) );
  NOR2_X1 U683 ( .A1(G286), .A2(n606), .ZN(n608) );
  NOR2_X1 U684 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U685 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U686 ( .A1(n609), .A2(G559), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n610), .A2(n945), .ZN(n611) );
  XNOR2_X1 U688 ( .A(n611), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U689 ( .A1(n967), .A2(G868), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G868), .A2(n945), .ZN(n612) );
  NOR2_X1 U691 ( .A1(G559), .A2(n612), .ZN(n613) );
  NOR2_X1 U692 ( .A1(n614), .A2(n613), .ZN(G282) );
  XOR2_X1 U693 ( .A(G2100), .B(KEYINPUT74), .Z(n624) );
  NAND2_X1 U694 ( .A1(G111), .A2(n892), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G135), .A2(n519), .ZN(n616) );
  NAND2_X1 U696 ( .A1(G99), .A2(n518), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U698 ( .A1(n891), .A2(G123), .ZN(n617) );
  XOR2_X1 U699 ( .A(KEYINPUT18), .B(n617), .Z(n618) );
  NOR2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U702 ( .A(n622), .B(KEYINPUT73), .ZN(n1011) );
  XNOR2_X1 U703 ( .A(n1011), .B(G2096), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(G156) );
  NAND2_X1 U705 ( .A1(G67), .A2(n649), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G93), .A2(n650), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G80), .A2(n651), .ZN(n628) );
  NAND2_X1 U709 ( .A1(G55), .A2(n656), .ZN(n627) );
  NAND2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n629) );
  OR2_X1 U711 ( .A1(n630), .A2(n629), .ZN(n668) );
  NAND2_X1 U712 ( .A1(n945), .A2(G559), .ZN(n666) );
  XOR2_X1 U713 ( .A(n967), .B(KEYINPUT75), .Z(n631) );
  XNOR2_X1 U714 ( .A(n666), .B(n631), .ZN(n632) );
  NOR2_X1 U715 ( .A1(G860), .A2(n632), .ZN(n633) );
  XNOR2_X1 U716 ( .A(n633), .B(KEYINPUT76), .ZN(n634) );
  XOR2_X1 U717 ( .A(n668), .B(n634), .Z(G145) );
  INV_X1 U718 ( .A(G303), .ZN(G166) );
  NAND2_X1 U719 ( .A1(G651), .A2(G74), .ZN(n636) );
  NAND2_X1 U720 ( .A1(G49), .A2(n656), .ZN(n635) );
  NAND2_X1 U721 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U722 ( .A1(n649), .A2(n637), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n638), .A2(G87), .ZN(n639) );
  NAND2_X1 U724 ( .A1(n640), .A2(n639), .ZN(G288) );
  NAND2_X1 U725 ( .A1(G73), .A2(n651), .ZN(n641) );
  XOR2_X1 U726 ( .A(KEYINPUT2), .B(n641), .Z(n646) );
  NAND2_X1 U727 ( .A1(G61), .A2(n649), .ZN(n643) );
  NAND2_X1 U728 ( .A1(G86), .A2(n650), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U730 ( .A(KEYINPUT77), .B(n644), .Z(n645) );
  NOR2_X1 U731 ( .A1(n646), .A2(n645), .ZN(n648) );
  NAND2_X1 U732 ( .A1(G48), .A2(n656), .ZN(n647) );
  NAND2_X1 U733 ( .A1(n648), .A2(n647), .ZN(G305) );
  AND2_X1 U734 ( .A1(n649), .A2(G60), .ZN(n655) );
  NAND2_X1 U735 ( .A1(G85), .A2(n650), .ZN(n653) );
  NAND2_X1 U736 ( .A1(G72), .A2(n651), .ZN(n652) );
  NAND2_X1 U737 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U738 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U739 ( .A1(G47), .A2(n656), .ZN(n657) );
  NAND2_X1 U740 ( .A1(n658), .A2(n657), .ZN(G290) );
  XNOR2_X1 U741 ( .A(n967), .B(G166), .ZN(n665) );
  XOR2_X1 U742 ( .A(KEYINPUT79), .B(KEYINPUT19), .Z(n659) );
  XNOR2_X1 U743 ( .A(G288), .B(n659), .ZN(n660) );
  XNOR2_X1 U744 ( .A(n660), .B(G305), .ZN(n663) );
  XNOR2_X1 U745 ( .A(n668), .B(G290), .ZN(n661) );
  XNOR2_X1 U746 ( .A(G299), .B(n661), .ZN(n662) );
  XNOR2_X1 U747 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U748 ( .A(n665), .B(n664), .ZN(n849) );
  XNOR2_X1 U749 ( .A(n666), .B(n849), .ZN(n667) );
  NAND2_X1 U750 ( .A1(n667), .A2(G868), .ZN(n671) );
  NAND2_X1 U751 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U753 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XOR2_X1 U754 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U755 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U757 ( .A1(n675), .A2(G2072), .ZN(n676) );
  XNOR2_X1 U758 ( .A(KEYINPUT80), .B(n676), .ZN(G158) );
  XNOR2_X1 U759 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U760 ( .A1(G235), .A2(G236), .ZN(n677) );
  XOR2_X1 U761 ( .A(KEYINPUT82), .B(n677), .Z(n678) );
  NOR2_X1 U762 ( .A1(G238), .A2(n678), .ZN(n679) );
  NAND2_X1 U763 ( .A1(G57), .A2(n679), .ZN(n846) );
  NAND2_X1 U764 ( .A1(G567), .A2(n846), .ZN(n680) );
  XNOR2_X1 U765 ( .A(n680), .B(KEYINPUT83), .ZN(n686) );
  NOR2_X1 U766 ( .A1(G220), .A2(G219), .ZN(n681) );
  XNOR2_X1 U767 ( .A(KEYINPUT22), .B(n681), .ZN(n682) );
  NAND2_X1 U768 ( .A1(n682), .A2(G96), .ZN(n683) );
  NOR2_X1 U769 ( .A1(G218), .A2(n683), .ZN(n684) );
  XNOR2_X1 U770 ( .A(KEYINPUT81), .B(n684), .ZN(n847) );
  AND2_X1 U771 ( .A1(G2106), .A2(n847), .ZN(n685) );
  NOR2_X1 U772 ( .A1(n686), .A2(n685), .ZN(G319) );
  INV_X1 U773 ( .A(G319), .ZN(n918) );
  NAND2_X1 U774 ( .A1(G483), .A2(G661), .ZN(n687) );
  NOR2_X1 U775 ( .A1(n918), .A2(n687), .ZN(n845) );
  NAND2_X1 U776 ( .A1(n845), .A2(G36), .ZN(G176) );
  NOR2_X1 U777 ( .A1(n688), .A2(G1384), .ZN(n689) );
  XNOR2_X1 U778 ( .A(n689), .B(KEYINPUT65), .ZN(n790) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n791) );
  INV_X1 U780 ( .A(n710), .ZN(n709) );
  NOR2_X1 U781 ( .A1(n709), .A2(G2084), .ZN(n749) );
  INV_X1 U782 ( .A(G8), .ZN(n691) );
  OR2_X1 U783 ( .A1(G1966), .A2(n691), .ZN(n692) );
  BUF_X1 U784 ( .A(n710), .Z(n704) );
  NOR2_X1 U785 ( .A1(n692), .A2(n704), .ZN(n693) );
  XNOR2_X1 U786 ( .A(n693), .B(KEYINPUT90), .ZN(n751) );
  XNOR2_X1 U787 ( .A(KEYINPUT96), .B(n694), .ZN(n695) );
  NAND2_X1 U788 ( .A1(n695), .A2(G8), .ZN(n696) );
  XNOR2_X1 U789 ( .A(KEYINPUT30), .B(n696), .ZN(n697) );
  NOR2_X1 U790 ( .A1(G168), .A2(n697), .ZN(n702) );
  NOR2_X1 U791 ( .A1(G1961), .A2(n704), .ZN(n699) );
  XOR2_X1 U792 ( .A(KEYINPUT25), .B(G2078), .Z(n931) );
  NOR2_X1 U793 ( .A1(n709), .A2(n931), .ZN(n698) );
  NOR2_X1 U794 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U795 ( .A(KEYINPUT91), .B(n700), .ZN(n730) );
  NOR2_X1 U796 ( .A1(G171), .A2(n730), .ZN(n701) );
  NOR2_X1 U797 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U798 ( .A(KEYINPUT31), .B(n703), .ZN(n737) );
  NAND2_X1 U799 ( .A1(G2072), .A2(n704), .ZN(n705) );
  XNOR2_X1 U800 ( .A(n705), .B(KEYINPUT27), .ZN(n707) );
  AND2_X1 U801 ( .A1(n709), .A2(G1956), .ZN(n706) );
  NOR2_X1 U802 ( .A1(n707), .A2(n706), .ZN(n723) );
  NOR2_X1 U803 ( .A1(n948), .A2(n723), .ZN(n708) );
  XOR2_X1 U804 ( .A(n708), .B(KEYINPUT28), .Z(n727) );
  NAND2_X1 U805 ( .A1(n709), .A2(G1341), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n710), .A2(G1996), .ZN(n711) );
  XNOR2_X1 U807 ( .A(n711), .B(KEYINPUT26), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U809 ( .A1(n714), .A2(n967), .ZN(n716) );
  NOR2_X1 U810 ( .A1(n716), .A2(n945), .ZN(n715) );
  XNOR2_X1 U811 ( .A(n715), .B(KEYINPUT93), .ZN(n722) );
  NAND2_X1 U812 ( .A1(n716), .A2(n945), .ZN(n720) );
  NOR2_X1 U813 ( .A1(G1348), .A2(n704), .ZN(n718) );
  NOR2_X1 U814 ( .A1(G2067), .A2(n709), .ZN(n717) );
  NOR2_X1 U815 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U816 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n948), .A2(n723), .ZN(n724) );
  NAND2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n727), .A2(n726), .ZN(n729) );
  XNOR2_X1 U821 ( .A(KEYINPUT29), .B(KEYINPUT94), .ZN(n728) );
  XNOR2_X1 U822 ( .A(n729), .B(n728), .ZN(n733) );
  AND2_X1 U823 ( .A1(n730), .A2(G171), .ZN(n731) );
  XNOR2_X1 U824 ( .A(n731), .B(KEYINPUT92), .ZN(n732) );
  NOR2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n735) );
  XNOR2_X1 U826 ( .A(n735), .B(n734), .ZN(n736) );
  XNOR2_X1 U827 ( .A(n738), .B(KEYINPUT97), .ZN(n750) );
  NAND2_X1 U828 ( .A1(n750), .A2(G286), .ZN(n739) );
  XNOR2_X1 U829 ( .A(n739), .B(KEYINPUT98), .ZN(n744) );
  NOR2_X1 U830 ( .A1(n709), .A2(G2090), .ZN(n741) );
  AND2_X1 U831 ( .A1(n709), .A2(G8), .ZN(n760) );
  INV_X1 U832 ( .A(n760), .ZN(n782) );
  NOR2_X1 U833 ( .A1(G1971), .A2(n782), .ZN(n740) );
  NOR2_X1 U834 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U835 ( .A1(n742), .A2(G303), .ZN(n743) );
  NAND2_X1 U836 ( .A1(n744), .A2(n743), .ZN(n746) );
  XNOR2_X1 U837 ( .A(n746), .B(n745), .ZN(n747) );
  NAND2_X1 U838 ( .A1(n747), .A2(G8), .ZN(n748) );
  NAND2_X1 U839 ( .A1(G8), .A2(n749), .ZN(n754) );
  INV_X1 U840 ( .A(n750), .ZN(n752) );
  NOR2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n773) );
  AND2_X1 U843 ( .A1(n773), .A2(n782), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n775), .A2(n755), .ZN(n759) );
  NOR2_X1 U845 ( .A1(G2090), .A2(G303), .ZN(n756) );
  NAND2_X1 U846 ( .A1(G8), .A2(n756), .ZN(n757) );
  OR2_X1 U847 ( .A1(n760), .A2(n757), .ZN(n758) );
  AND2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n788) );
  INV_X1 U849 ( .A(KEYINPUT33), .ZN(n763) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n956) );
  NAND2_X1 U851 ( .A1(n760), .A2(n956), .ZN(n761) );
  NOR2_X1 U852 ( .A1(n763), .A2(n761), .ZN(n762) );
  XNOR2_X1 U853 ( .A(n762), .B(KEYINPUT101), .ZN(n766) );
  INV_X1 U854 ( .A(n766), .ZN(n764) );
  OR2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n776) );
  INV_X1 U856 ( .A(n776), .ZN(n769) );
  NAND2_X1 U857 ( .A1(G288), .A2(G1976), .ZN(n765) );
  XOR2_X1 U858 ( .A(KEYINPUT100), .B(n765), .Z(n955) );
  NOR2_X1 U859 ( .A1(n782), .A2(n955), .ZN(n767) );
  AND2_X1 U860 ( .A1(n767), .A2(n766), .ZN(n768) );
  OR2_X1 U861 ( .A1(n769), .A2(n768), .ZN(n771) );
  XNOR2_X1 U862 ( .A(G1981), .B(G305), .ZN(n961) );
  INV_X1 U863 ( .A(n961), .ZN(n770) );
  NAND2_X1 U864 ( .A1(n771), .A2(n770), .ZN(n779) );
  INV_X1 U865 ( .A(n779), .ZN(n772) );
  AND2_X1 U866 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U867 ( .A1(n775), .A2(n774), .ZN(n786) );
  NOR2_X1 U868 ( .A1(G1971), .A2(G303), .ZN(n954) );
  NOR2_X1 U869 ( .A1(n956), .A2(n954), .ZN(n777) );
  AND2_X1 U870 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U871 ( .A1(n779), .A2(n778), .ZN(n784) );
  NOR2_X1 U872 ( .A1(G1981), .A2(G305), .ZN(n780) );
  XOR2_X1 U873 ( .A(n780), .B(KEYINPUT24), .Z(n781) );
  NOR2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n785) );
  AND2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n825) );
  XOR2_X1 U878 ( .A(G1986), .B(KEYINPUT85), .Z(n789) );
  XNOR2_X1 U879 ( .A(G290), .B(n789), .ZN(n953) );
  NOR2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n836) );
  NAND2_X1 U881 ( .A1(n953), .A2(n836), .ZN(n823) );
  NAND2_X1 U882 ( .A1(G105), .A2(n518), .ZN(n793) );
  XNOR2_X1 U883 ( .A(n793), .B(KEYINPUT38), .ZN(n800) );
  NAND2_X1 U884 ( .A1(G129), .A2(n891), .ZN(n795) );
  NAND2_X1 U885 ( .A1(G117), .A2(n892), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n798) );
  NAND2_X1 U887 ( .A1(G141), .A2(n519), .ZN(n796) );
  XNOR2_X1 U888 ( .A(KEYINPUT87), .B(n796), .ZN(n797) );
  NOR2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n800), .A2(n799), .ZN(n887) );
  NAND2_X1 U891 ( .A1(n887), .A2(G1996), .ZN(n808) );
  NAND2_X1 U892 ( .A1(G131), .A2(n519), .ZN(n802) );
  NAND2_X1 U893 ( .A1(G107), .A2(n892), .ZN(n801) );
  NAND2_X1 U894 ( .A1(n802), .A2(n801), .ZN(n806) );
  NAND2_X1 U895 ( .A1(G119), .A2(n891), .ZN(n804) );
  NAND2_X1 U896 ( .A1(G95), .A2(n518), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n805) );
  OR2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n910) );
  NAND2_X1 U899 ( .A1(G1991), .A2(n910), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U901 ( .A(n809), .B(KEYINPUT88), .ZN(n1004) );
  NAND2_X1 U902 ( .A1(n1004), .A2(n836), .ZN(n810) );
  XNOR2_X1 U903 ( .A(n810), .B(KEYINPUT89), .ZN(n829) );
  INV_X1 U904 ( .A(n829), .ZN(n821) );
  XNOR2_X1 U905 ( .A(G2067), .B(KEYINPUT37), .ZN(n834) );
  NAND2_X1 U906 ( .A1(G128), .A2(n891), .ZN(n812) );
  NAND2_X1 U907 ( .A1(G116), .A2(n892), .ZN(n811) );
  NAND2_X1 U908 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U909 ( .A(n813), .B(KEYINPUT35), .ZN(n818) );
  NAND2_X1 U910 ( .A1(G140), .A2(n519), .ZN(n815) );
  NAND2_X1 U911 ( .A1(G104), .A2(n518), .ZN(n814) );
  NAND2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U913 ( .A(KEYINPUT34), .B(n816), .Z(n817) );
  NAND2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n819) );
  XOR2_X1 U915 ( .A(n819), .B(KEYINPUT36), .Z(n888) );
  OR2_X1 U916 ( .A1(n834), .A2(n888), .ZN(n820) );
  XOR2_X1 U917 ( .A(KEYINPUT86), .B(n820), .Z(n1025) );
  NAND2_X1 U918 ( .A1(n836), .A2(n1025), .ZN(n832) );
  AND2_X1 U919 ( .A1(n821), .A2(n832), .ZN(n822) );
  AND2_X1 U920 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n839) );
  NOR2_X1 U922 ( .A1(G1996), .A2(n887), .ZN(n1007) );
  NOR2_X1 U923 ( .A1(G1991), .A2(n910), .ZN(n1012) );
  NOR2_X1 U924 ( .A1(G1986), .A2(G290), .ZN(n826) );
  XNOR2_X1 U925 ( .A(KEYINPUT102), .B(n826), .ZN(n827) );
  NOR2_X1 U926 ( .A1(n1012), .A2(n827), .ZN(n828) );
  NOR2_X1 U927 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U928 ( .A1(n1007), .A2(n830), .ZN(n831) );
  XNOR2_X1 U929 ( .A(n831), .B(KEYINPUT39), .ZN(n833) );
  NAND2_X1 U930 ( .A1(n833), .A2(n832), .ZN(n835) );
  NAND2_X1 U931 ( .A1(n888), .A2(n834), .ZN(n1003) );
  NAND2_X1 U932 ( .A1(n835), .A2(n1003), .ZN(n837) );
  NAND2_X1 U933 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U935 ( .A(KEYINPUT40), .B(n840), .ZN(G329) );
  NAND2_X1 U936 ( .A1(n841), .A2(G2106), .ZN(n842) );
  XNOR2_X1 U937 ( .A(n842), .B(KEYINPUT104), .ZN(G217) );
  AND2_X1 U938 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U939 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U940 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U941 ( .A1(n845), .A2(n844), .ZN(G188) );
  INV_X1 U943 ( .A(G96), .ZN(G221) );
  NOR2_X1 U944 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U945 ( .A(KEYINPUT105), .B(n848), .ZN(G261) );
  INV_X1 U946 ( .A(G261), .ZN(G325) );
  XOR2_X1 U947 ( .A(n849), .B(G286), .Z(n851) );
  XNOR2_X1 U948 ( .A(n945), .B(G171), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n852) );
  NOR2_X1 U950 ( .A1(G37), .A2(n852), .ZN(G397) );
  XOR2_X1 U951 ( .A(G2100), .B(KEYINPUT43), .Z(n854) );
  XNOR2_X1 U952 ( .A(G2090), .B(G2678), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U954 ( .A(n855), .B(KEYINPUT42), .Z(n857) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U957 ( .A(KEYINPUT106), .B(G2096), .Z(n859) );
  XNOR2_X1 U958 ( .A(G2078), .B(G2084), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(G227) );
  XOR2_X1 U961 ( .A(G1976), .B(G1961), .Z(n863) );
  XNOR2_X1 U962 ( .A(G1996), .B(G1956), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U964 ( .A(G1981), .B(G1971), .Z(n865) );
  XNOR2_X1 U965 ( .A(G1986), .B(G1966), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U967 ( .A(n867), .B(n866), .Z(n869) );
  XNOR2_X1 U968 ( .A(G2474), .B(KEYINPUT41), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n871) );
  XOR2_X1 U970 ( .A(G1991), .B(KEYINPUT107), .Z(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(G229) );
  NAND2_X1 U972 ( .A1(n891), .A2(G124), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n872), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G112), .A2(n892), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G136), .A2(n519), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G100), .A2(n518), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U979 ( .A1(n878), .A2(n877), .ZN(G162) );
  NAND2_X1 U980 ( .A1(G139), .A2(n519), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G103), .A2(n518), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G127), .A2(n891), .ZN(n882) );
  NAND2_X1 U984 ( .A1(G115), .A2(n892), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U986 ( .A(KEYINPUT47), .B(n883), .Z(n884) );
  NOR2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U988 ( .A(KEYINPUT109), .B(n886), .Z(n1016) );
  XNOR2_X1 U989 ( .A(n887), .B(n1016), .ZN(n890) );
  XOR2_X1 U990 ( .A(G160), .B(n888), .Z(n889) );
  XNOR2_X1 U991 ( .A(n890), .B(n889), .ZN(n904) );
  NAND2_X1 U992 ( .A1(G130), .A2(n891), .ZN(n894) );
  NAND2_X1 U993 ( .A1(G118), .A2(n892), .ZN(n893) );
  NAND2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n902) );
  NAND2_X1 U995 ( .A1(G142), .A2(n519), .ZN(n898) );
  NAND2_X1 U996 ( .A1(G106), .A2(n518), .ZN(n897) );
  NAND2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U998 ( .A(KEYINPUT108), .B(n899), .Z(n900) );
  XNOR2_X1 U999 ( .A(KEYINPUT45), .B(n900), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1001 ( .A(n904), .B(n903), .Z(n906) );
  XNOR2_X1 U1002 ( .A(G164), .B(G162), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n914) );
  XOR2_X1 U1004 ( .A(KEYINPUT112), .B(KEYINPUT111), .Z(n908) );
  XNOR2_X1 U1005 ( .A(n1011), .B(KEYINPUT110), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(KEYINPUT46), .B(n909), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n910), .B(KEYINPUT48), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n915), .ZN(G395) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(G397), .A2(n917), .ZN(n922) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n918), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(KEYINPUT113), .B(n919), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G395), .A2(n920), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1021 ( .A(KEYINPUT55), .B(KEYINPUT115), .ZN(n1027) );
  XNOR2_X1 U1022 ( .A(G2067), .B(G26), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(G1991), .B(G25), .ZN(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n930) );
  XOR2_X1 U1025 ( .A(G1996), .B(G32), .Z(n925) );
  NAND2_X1 U1026 ( .A1(n925), .A2(G28), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(KEYINPUT116), .B(G2072), .ZN(n926) );
  XNOR2_X1 U1028 ( .A(G33), .B(n926), .ZN(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(G27), .B(n931), .ZN(n932) );
  NOR2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1033 ( .A(KEYINPUT53), .B(n934), .Z(n937) );
  XOR2_X1 U1034 ( .A(KEYINPUT54), .B(G34), .Z(n935) );
  XNOR2_X1 U1035 ( .A(G2084), .B(n935), .ZN(n936) );
  NAND2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(G35), .B(G2090), .ZN(n938) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1039 ( .A(n1027), .B(n940), .Z(n942) );
  INV_X1 U1040 ( .A(G29), .ZN(n941) );
  NAND2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1042 ( .A1(n943), .A2(G11), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(n944), .B(KEYINPUT117), .ZN(n975) );
  XNOR2_X1 U1044 ( .A(G171), .B(G1961), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(G1348), .B(n945), .ZN(n946) );
  NAND2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(n948), .B(G1956), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(G1971), .A2(G303), .ZN(n949) );
  NAND2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n966) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n959) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n957), .B(KEYINPUT118), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n964) );
  XOR2_X1 U1055 ( .A(G1966), .B(G168), .Z(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n962), .B(KEYINPUT57), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n970) );
  XOR2_X1 U1060 ( .A(n967), .B(G1341), .Z(n968) );
  XNOR2_X1 U1061 ( .A(KEYINPUT119), .B(n968), .ZN(n969) );
  NOR2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1063 ( .A(KEYINPUT120), .B(n971), .Z(n973) );
  XNOR2_X1 U1064 ( .A(KEYINPUT56), .B(G16), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n1001) );
  XOR2_X1 U1067 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n998) );
  XNOR2_X1 U1068 ( .A(G1348), .B(KEYINPUT59), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(n976), .B(G4), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(G1341), .B(G19), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(G6), .B(G1981), .ZN(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n983) );
  XOR2_X1 U1074 ( .A(G20), .B(G1956), .Z(n981) );
  XNOR2_X1 U1075 ( .A(KEYINPUT121), .B(n981), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1077 ( .A(KEYINPUT60), .B(n984), .Z(n986) );
  XNOR2_X1 U1078 ( .A(G1966), .B(G21), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n996) );
  XNOR2_X1 U1080 ( .A(G1971), .B(G22), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(G23), .B(G1976), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1083 ( .A(KEYINPUT122), .B(n989), .Z(n991) );
  XNOR2_X1 U1084 ( .A(G1986), .B(G24), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1086 ( .A(KEYINPUT58), .B(n992), .Z(n994) );
  XNOR2_X1 U1087 ( .A(G1961), .B(G5), .ZN(n993) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(n998), .B(n997), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(G16), .A2(n999), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(KEYINPUT124), .B(n1002), .ZN(n1031) );
  INV_X1 U1094 ( .A(n1003), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1023) );
  XOR2_X1 U1096 ( .A(G160), .B(G2084), .Z(n1010) );
  XOR2_X1 U1097 ( .A(G2090), .B(G162), .Z(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1099 ( .A(KEYINPUT51), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(n1013), .B(KEYINPUT114), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1021) );
  XOR2_X1 U1104 ( .A(G2072), .B(n1016), .Z(n1018) );
  XOR2_X1 U1105 ( .A(G164), .B(G2078), .Z(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1107 ( .A(KEYINPUT50), .B(n1019), .Z(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1111 ( .A(KEYINPUT52), .B(n1026), .ZN(n1028) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(G29), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1115 ( .A(n1032), .B(KEYINPUT126), .ZN(n1034) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(KEYINPUT125), .Z(n1033) );
  XNOR2_X1 U1117 ( .A(n1034), .B(n1033), .ZN(G150) );
  INV_X1 U1118 ( .A(G150), .ZN(G311) );
  INV_X1 U1119 ( .A(G171), .ZN(G301) );
endmodule

