//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1222, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296, new_n1297;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  NAND2_X1  g0006(.A1(G116), .A2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  INV_X1    g0008(.A(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT68), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n213), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT66), .B(G68), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT67), .B(G238), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  AND3_X1   g0023(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n224));
  AOI21_X1  g0024(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G58), .ZN(new_n229));
  INV_X1    g0029(.A(G68), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT65), .Z(new_n233));
  AOI211_X1 g0033(.A(new_n206), .B(new_n223), .C1(new_n228), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(KEYINPUT69), .B(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n238), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT17), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(new_n224), .B2(new_n225), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n217), .A2(G1698), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n254), .B(new_n255), .C1(G223), .C2(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G87), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n257), .B(KEYINPUT80), .Z(new_n258));
  AOI21_X1  g0058(.A(new_n253), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT70), .B(G41), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n260), .B(G274), .C1(new_n261), .C2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n252), .A2(G1), .A3(G13), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G232), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n259), .A2(new_n263), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G190), .ZN(new_n270));
  XOR2_X1   g0070(.A(KEYINPUT8), .B(G58), .Z(new_n271));
  NAND2_X1  g0071(.A1(G1), .A2(G13), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT64), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n260), .A2(G20), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n271), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT79), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(KEYINPUT3), .ZN(new_n290));
  OAI211_X1 g0090(.A(KEYINPUT7), .B(new_n227), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(KEYINPUT3), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n287), .A2(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(KEYINPUT7), .B1(new_n295), .B2(new_n227), .ZN(new_n296));
  OAI21_X1  g0096(.A(G68), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n231), .B1(new_n219), .B2(new_n229), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n298), .A2(G20), .B1(G159), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n297), .A2(new_n300), .A3(KEYINPUT16), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n277), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT7), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n254), .B2(G20), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT78), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(new_n291), .ZN(new_n306));
  AND2_X1   g0106(.A1(KEYINPUT66), .A2(G68), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT66), .A2(G68), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n295), .A2(KEYINPUT78), .A3(KEYINPUT7), .A4(new_n227), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n306), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(KEYINPUT16), .B1(new_n311), .B2(new_n300), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n270), .B(new_n286), .C1(new_n302), .C2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G200), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n269), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n251), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n284), .B(KEYINPUT79), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n311), .A2(new_n300), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT16), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n277), .ZN(new_n321));
  INV_X1    g0121(.A(new_n231), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(new_n309), .B2(G58), .ZN(new_n323));
  INV_X1    g0123(.A(G159), .ZN(new_n324));
  INV_X1    g0124(.A(new_n299), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n323), .A2(new_n227), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n230), .B1(new_n304), .B2(new_n291), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n321), .B1(new_n328), .B2(KEYINPUT16), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n317), .B1(new_n320), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n315), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n330), .A2(KEYINPUT17), .A3(new_n331), .A4(new_n270), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n286), .B1(new_n302), .B2(new_n312), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT71), .B(G179), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NOR4_X1   g0135(.A1(new_n259), .A2(new_n263), .A3(new_n335), .A4(new_n268), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  OR3_X1    g0137(.A1(new_n259), .A2(new_n263), .A3(new_n268), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n333), .A2(KEYINPUT18), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT18), .B1(new_n333), .B2(new_n339), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n316), .B(new_n332), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT77), .ZN(new_n343));
  INV_X1    g0143(.A(G1698), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n217), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n267), .A2(G1698), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n254), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G97), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n253), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n264), .A2(G238), .A3(new_n265), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n262), .A2(new_n350), .ZN(new_n351));
  XOR2_X1   g0151(.A(KEYINPUT75), .B(KEYINPUT13), .Z(new_n352));
  NOR3_X1   g0152(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT13), .B1(new_n349), .B2(new_n351), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT76), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT76), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(KEYINPUT13), .C1(new_n349), .C2(new_n351), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n354), .A2(new_n356), .A3(G190), .A4(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n309), .A2(new_n227), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n227), .A2(G33), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n325), .A2(new_n216), .B1(new_n361), .B2(new_n208), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n277), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT11), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n363), .B(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n277), .A2(new_n279), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT12), .ZN(new_n367));
  OAI21_X1  g0167(.A(G68), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n282), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n219), .A2(new_n369), .A3(KEYINPUT12), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n368), .B(new_n370), .C1(KEYINPUT12), .C2(new_n369), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n352), .ZN(new_n373));
  INV_X1    g0173(.A(new_n349), .ZN(new_n374));
  INV_X1    g0174(.A(new_n351), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(G200), .B1(new_n376), .B2(new_n353), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n359), .A2(new_n372), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(G169), .B1(new_n376), .B2(new_n353), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT14), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n354), .A2(new_n356), .A3(G179), .A4(new_n358), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT14), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n382), .B(G169), .C1(new_n376), .C2(new_n353), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n372), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n378), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n342), .B1(new_n343), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n266), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n263), .B1(G244), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n344), .A2(G232), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n254), .B(new_n390), .C1(new_n220), .C2(new_n344), .ZN(new_n391));
  INV_X1    g0191(.A(new_n253), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n391), .B(new_n392), .C1(G107), .C2(new_n254), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G200), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n281), .A2(new_n325), .B1(new_n227), .B2(new_n208), .ZN(new_n396));
  XOR2_X1   g0196(.A(KEYINPUT15), .B(G87), .Z(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(new_n361), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n277), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n366), .A2(G77), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n369), .A2(new_n208), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT72), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n400), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G190), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n395), .B(new_n405), .C1(new_n406), .C2(new_n394), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n394), .A2(new_n337), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n408), .B(new_n404), .C1(new_n335), .C2(new_n394), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT73), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n344), .A2(G222), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G223), .A2(G1698), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n254), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n392), .B(new_n414), .C1(G77), .C2(new_n254), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n388), .A2(G226), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n262), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n334), .ZN(new_n419));
  OAI21_X1  g0219(.A(G20), .B1(new_n231), .B2(G50), .ZN(new_n420));
  INV_X1    g0220(.A(G150), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n420), .B1(new_n421), .B2(new_n325), .C1(new_n361), .C2(new_n281), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(new_n277), .B1(new_n366), .B2(G50), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(G50), .B2(new_n282), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n417), .A2(new_n337), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n419), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n424), .B(KEYINPUT9), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n417), .A2(G200), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n418), .A2(G190), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n428), .A2(KEYINPUT74), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT10), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT74), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n424), .A2(KEYINPUT9), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n424), .A2(KEYINPUT9), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT10), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n429), .A4(new_n430), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n427), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n387), .A2(new_n411), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n386), .A2(new_n343), .ZN(new_n441));
  OR3_X1    g0241(.A1(new_n440), .A2(KEYINPUT81), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT81), .B1(new_n440), .B2(new_n441), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n211), .B1(new_n445), .B2(G1), .ZN(new_n446));
  INV_X1    g0246(.A(G274), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n260), .A2(new_n447), .A3(G45), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n264), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  OR2_X1    g0249(.A1(G238), .A2(G1698), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n209), .A2(G1698), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n293), .A2(new_n450), .A3(new_n294), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G116), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n449), .B1(new_n454), .B2(new_n392), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(G169), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  INV_X1    g0257(.A(G107), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n210), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n348), .A2(new_n227), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT19), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n293), .A2(new_n294), .A3(new_n227), .A4(G68), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT19), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n348), .B2(G20), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n277), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n260), .A2(G33), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n321), .A2(new_n282), .A3(new_n397), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n398), .A2(new_n369), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT82), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT82), .A4(new_n469), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n456), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n455), .A2(new_n334), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n274), .A2(new_n275), .A3(new_n276), .A4(new_n467), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(new_n369), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G87), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n466), .A2(new_n478), .A3(new_n469), .ZN(new_n479));
  INV_X1    g0279(.A(new_n455), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n479), .B1(G200), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT83), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n455), .B2(G190), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n253), .B1(new_n453), .B2(new_n452), .ZN(new_n484));
  NOR4_X1   g0284(.A1(new_n484), .A2(KEYINPUT83), .A3(new_n406), .A4(new_n449), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n474), .A2(new_n475), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n306), .A2(G107), .A3(new_n310), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n458), .A2(KEYINPUT6), .A3(G97), .ZN(new_n489));
  XOR2_X1   g0289(.A(G97), .B(G107), .Z(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(KEYINPUT6), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(G20), .B1(G77), .B2(new_n299), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n277), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n369), .A2(new_n457), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n477), .A2(G97), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n293), .A2(new_n294), .A3(G244), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(G1698), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n254), .A2(G244), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G283), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n254), .A2(G250), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n344), .B1(new_n505), .B2(KEYINPUT4), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n392), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n264), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT5), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n260), .B(G45), .C1(new_n509), .C2(G41), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G41), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT70), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT70), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G41), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n515), .A3(new_n509), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n508), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n510), .B1(new_n261), .B2(new_n509), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n517), .A2(G257), .B1(G274), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n507), .A2(new_n335), .A3(new_n519), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n513), .A2(new_n515), .A3(new_n509), .ZN(new_n521));
  OAI211_X1 g0321(.A(G257), .B(new_n264), .C1(new_n521), .C2(new_n510), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n518), .A2(G274), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n498), .A2(new_n499), .B1(G33), .B2(G283), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n499), .B1(new_n254), .B2(G250), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n525), .B(new_n502), .C1(new_n344), .C2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n524), .B1(new_n392), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n520), .B1(new_n528), .B2(new_n337), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n497), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n507), .A2(new_n406), .A3(new_n519), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n528), .B2(G200), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n493), .A2(new_n277), .B1(new_n457), .B2(new_n369), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(new_n533), .A3(new_n496), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n487), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n293), .A2(new_n294), .A3(new_n227), .A4(G87), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT22), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT22), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n254), .A2(new_n538), .A3(new_n227), .A4(G87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n227), .A2(G107), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n541), .B(KEYINPUT23), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n227), .A2(G33), .A3(G116), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT24), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n540), .A2(KEYINPUT24), .A3(new_n542), .A4(new_n543), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(new_n277), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n477), .A2(G107), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n282), .A2(G107), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n550), .B(KEYINPUT25), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n517), .A2(G264), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT87), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n517), .A2(KEYINPUT87), .A3(G264), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n211), .A2(new_n344), .ZN(new_n558));
  INV_X1    g0358(.A(G257), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G1698), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n293), .A2(new_n558), .A3(new_n294), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G33), .A2(G294), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT85), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT85), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n561), .A2(new_n565), .A3(new_n562), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n392), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n557), .A2(new_n523), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n314), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n567), .A2(KEYINPUT86), .B1(G274), .B2(new_n518), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n561), .A2(new_n565), .A3(new_n562), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n565), .B1(new_n561), .B2(new_n562), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n571), .A2(new_n572), .A3(new_n253), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT86), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n570), .A2(new_n575), .A3(new_n406), .A4(new_n553), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n552), .B1(new_n569), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n535), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(G116), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n476), .A2(new_n579), .A3(new_n369), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(G20), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n503), .B(new_n227), .C1(G33), .C2(new_n457), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n277), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT20), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n277), .A2(KEYINPUT20), .A3(new_n581), .A4(new_n582), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n580), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G116), .B2(new_n282), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G264), .A2(G1698), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n254), .B(new_n589), .C1(new_n559), .C2(G1698), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n590), .B(new_n392), .C1(G303), .C2(new_n254), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n517), .A2(G270), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(G179), .A4(new_n523), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT84), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n588), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n282), .A2(G116), .ZN(new_n597));
  AOI211_X1 g0397(.A(new_n597), .B(new_n580), .C1(new_n585), .C2(new_n586), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT84), .B1(new_n598), .B2(new_n593), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT21), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n591), .A2(new_n523), .A3(new_n592), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G169), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n601), .B1(new_n603), .B2(new_n598), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n588), .A2(KEYINPUT21), .A3(G169), .A4(new_n602), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n602), .A2(G200), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n606), .B(new_n598), .C1(new_n406), .C2(new_n602), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n600), .A2(new_n604), .A3(new_n605), .A4(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n548), .A2(new_n551), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n523), .B1(new_n573), .B2(new_n574), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n553), .B1(new_n567), .B2(KEYINPUT86), .ZN(new_n611));
  OAI21_X1  g0411(.A(G169), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n557), .A2(G179), .A3(new_n523), .A4(new_n567), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n609), .A2(new_n549), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n444), .A2(new_n578), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n616), .B(KEYINPUT88), .ZN(G372));
  AND2_X1   g0417(.A1(new_n530), .A2(new_n534), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n569), .A2(new_n576), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(new_n549), .A3(new_n609), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT89), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n618), .A2(new_n620), .A3(new_n621), .A4(new_n487), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT89), .B1(new_n535), .B2(new_n577), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n612), .A2(new_n613), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n552), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n622), .A2(new_n623), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n474), .A2(new_n475), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  INV_X1    g0431(.A(new_n487), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n631), .B1(new_n632), .B2(new_n530), .ZN(new_n633));
  INV_X1    g0433(.A(new_n530), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(KEYINPUT26), .A3(new_n487), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n630), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n444), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT90), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n340), .B2(new_n341), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n333), .A2(new_n339), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT18), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n333), .A2(new_n339), .A3(KEYINPUT18), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(KEYINPUT90), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT91), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n409), .B(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n378), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n647), .A2(new_n648), .B1(new_n385), .B2(new_n384), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n332), .A2(new_n316), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n640), .B(new_n645), .C1(new_n649), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n432), .A2(new_n438), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n427), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n638), .A2(new_n654), .ZN(G369));
  INV_X1    g0455(.A(G13), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n656), .A2(G1), .A3(G20), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT27), .ZN(new_n658));
  OR3_X1    g0458(.A1(new_n657), .A2(KEYINPUT92), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G213), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n657), .B2(new_n658), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT92), .B1(new_n657), .B2(new_n658), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n552), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n627), .B1(new_n577), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n665), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n614), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n625), .A2(new_n665), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n598), .A2(new_n668), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n624), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n608), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n669), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n671), .B2(new_n667), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT93), .ZN(G399));
  INV_X1    g0481(.A(new_n204), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n261), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n459), .A2(G116), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G1), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n232), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT94), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n665), .B1(new_n629), .B2(new_n636), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT29), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT97), .B1(new_n614), .B2(new_n624), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT97), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n604), .A2(new_n605), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n627), .A2(new_n693), .A3(new_n694), .A4(new_n600), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(new_n578), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n636), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(KEYINPUT29), .A3(new_n668), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n691), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n578), .A2(new_n615), .A3(new_n668), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT96), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n594), .A2(new_n567), .A3(new_n557), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n528), .A2(new_n455), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT95), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OR3_X1    g0507(.A1(new_n703), .A2(new_n704), .A3(new_n702), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n602), .A2(new_n334), .ZN(new_n709));
  INV_X1    g0509(.A(new_n528), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n568), .A2(new_n709), .A3(new_n710), .A4(new_n480), .ZN(new_n711));
  OAI211_X1 g0511(.A(KEYINPUT95), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n707), .A2(new_n708), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n665), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT96), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n578), .A2(new_n615), .A3(new_n717), .A4(new_n668), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n708), .A2(new_n711), .A3(new_n705), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n701), .A2(new_n716), .A3(new_n718), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G330), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n699), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n689), .B1(new_n723), .B2(G1), .ZN(G364));
  OR2_X1    g0524(.A1(new_n675), .A2(G330), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n656), .A2(G20), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G45), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n684), .A2(G1), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n725), .A2(new_n676), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n226), .B1(G20), .B2(new_n337), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n227), .A2(G179), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G190), .A2(G200), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G329), .ZN(new_n736));
  INV_X1    g0536(.A(G303), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n732), .A2(G190), .A3(G200), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n334), .A2(new_n227), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G200), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G190), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(KEYINPUT33), .B(G317), .Z(new_n743));
  OAI221_X1 g0543(.A(new_n736), .B1(new_n737), .B2(new_n738), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n740), .A2(new_n406), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n744), .B1(G326), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G322), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n406), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n739), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n746), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  OR3_X1    g0550(.A1(new_n406), .A2(G179), .A3(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n254), .B(new_n750), .C1(G294), .C2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G283), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n732), .A2(new_n406), .A3(G200), .ZN(new_n755));
  INV_X1    g0555(.A(G311), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n739), .A2(new_n733), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n753), .B1(new_n754), .B2(new_n755), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n757), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n745), .A2(G50), .B1(new_n759), .B2(G77), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(new_n229), .B2(new_n749), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT98), .Z(new_n762));
  INV_X1    g0562(.A(new_n755), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G107), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n735), .A2(G159), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n741), .A2(G68), .B1(KEYINPUT32), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n752), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n766), .B1(KEYINPUT32), .B2(new_n765), .C1(new_n457), .C2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n738), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n768), .B1(G87), .B2(new_n769), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n762), .A2(new_n254), .A3(new_n764), .A4(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n731), .B1(new_n758), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n675), .A2(new_n776), .ZN(new_n777));
  OR3_X1    g0577(.A1(new_n772), .A2(new_n728), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n233), .A2(new_n445), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n682), .A2(new_n254), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n779), .B(new_n780), .C1(new_n246), .C2(new_n445), .ZN(new_n781));
  INV_X1    g0581(.A(G355), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n254), .A2(new_n204), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n781), .B1(G116), .B2(new_n204), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n730), .A2(new_n775), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n729), .B1(new_n778), .B2(new_n786), .ZN(G396));
  NAND2_X1  g0587(.A1(new_n404), .A2(new_n665), .ZN(new_n788));
  AND3_X1   g0588(.A1(new_n407), .A2(new_n409), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n788), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(new_n647), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n690), .B(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(new_n722), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n728), .ZN(new_n794));
  INV_X1    g0594(.A(new_n749), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G143), .A2(new_n795), .B1(new_n759), .B2(G159), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G137), .A2(new_n745), .B1(new_n741), .B2(G150), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n797), .A2(KEYINPUT100), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(KEYINPUT100), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n796), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT34), .ZN(new_n801));
  INV_X1    g0601(.A(G132), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n755), .A2(new_n230), .B1(new_n734), .B2(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n295), .B(new_n803), .C1(G50), .C2(new_n769), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n801), .B(new_n804), .C1(new_n229), .C2(new_n767), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n741), .A2(G283), .B1(G87), .B2(new_n763), .ZN(new_n806));
  INV_X1    g0606(.A(G294), .ZN(new_n807));
  INV_X1    g0607(.A(new_n745), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n806), .B1(new_n807), .B2(new_n749), .C1(new_n737), .C2(new_n808), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n767), .A2(new_n457), .B1(new_n738), .B2(new_n458), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n809), .A2(new_n254), .A3(new_n810), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n811), .B1(new_n579), .B2(new_n757), .C1(new_n756), .C2(new_n734), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n731), .B1(new_n805), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n791), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n774), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n813), .A2(new_n815), .A3(new_n728), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n731), .A2(new_n774), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT99), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n816), .B1(G77), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n794), .A2(new_n819), .ZN(G384));
  NAND2_X1  g0620(.A1(new_n384), .A2(new_n385), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n665), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n328), .A2(KEYINPUT16), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n284), .B1(new_n302), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n663), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n342), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n824), .B1(new_n339), .B2(new_n825), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n320), .A2(new_n329), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n829), .A2(new_n331), .A3(new_n270), .A4(new_n286), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n828), .A2(new_n830), .A3(KEYINPUT37), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n333), .A2(new_n825), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n830), .A2(new_n641), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT37), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n827), .A2(new_n831), .A3(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT38), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n827), .A2(KEYINPUT38), .A3(new_n831), .A4(new_n835), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n838), .A2(KEYINPUT39), .A3(new_n839), .ZN(new_n840));
  AND4_X1   g0640(.A1(KEYINPUT38), .A2(new_n827), .A3(new_n831), .A4(new_n835), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n650), .A2(new_n640), .A3(new_n645), .ZN(new_n842));
  INV_X1    g0642(.A(new_n832), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT105), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n833), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n830), .A2(new_n641), .A3(new_n832), .A4(KEYINPUT105), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n830), .A2(new_n639), .A3(new_n832), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n846), .A2(KEYINPUT37), .A3(new_n849), .A4(new_n847), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n844), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n841), .B1(new_n853), .B2(new_n837), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n822), .B(new_n840), .C1(new_n854), .C2(KEYINPUT39), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n640), .A2(new_n645), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n663), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n637), .A2(new_n668), .A3(new_n814), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n409), .A2(new_n665), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT103), .B1(new_n372), .B2(new_n668), .ZN(new_n862));
  OR3_X1    g0662(.A1(new_n372), .A2(KEYINPUT103), .A3(new_n668), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n821), .A2(new_n648), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT104), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT104), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n386), .A2(new_n866), .A3(new_n862), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n384), .A2(new_n385), .A3(new_n665), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n838), .A2(new_n839), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n861), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n855), .A2(new_n857), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n444), .A2(new_n691), .A3(new_n698), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n654), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n874), .B(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n701), .A2(new_n716), .A3(new_n718), .A4(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n880), .A2(new_n814), .A3(new_n870), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n853), .A2(new_n837), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n839), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n878), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT40), .B1(new_n838), .B2(new_n839), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n880), .A2(new_n814), .A3(new_n870), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(G330), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n444), .A2(G330), .A3(new_n880), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT40), .B1(new_n887), .B2(new_n854), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n885), .A2(new_n814), .A3(new_n880), .A4(new_n870), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(new_n444), .A3(new_n880), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n877), .B(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n260), .B2(new_n726), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n208), .B(new_n232), .C1(new_n309), .C2(G58), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n216), .A2(G68), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT102), .ZN(new_n901));
  OAI211_X1 g0701(.A(G1), .B(new_n656), .C1(new_n899), .C2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n579), .B1(new_n491), .B2(KEYINPUT35), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n903), .B(new_n228), .C1(KEYINPUT35), .C2(new_n491), .ZN(new_n904));
  XOR2_X1   g0704(.A(KEYINPUT101), .B(KEYINPUT36), .Z(new_n905));
  XNOR2_X1  g0705(.A(new_n904), .B(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n898), .A2(new_n902), .A3(new_n906), .ZN(G367));
  OAI21_X1  g0707(.A(new_n295), .B1(new_n749), .B2(new_n737), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n808), .A2(new_n756), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT46), .B1(new_n769), .B2(G116), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n769), .A2(KEYINPUT46), .A3(G116), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n763), .A2(G97), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n911), .B(new_n912), .C1(new_n757), .C2(new_n754), .ZN(new_n913));
  OR3_X1    g0713(.A1(new_n909), .A2(new_n910), .A3(new_n913), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n908), .B(new_n914), .C1(G294), .C2(new_n741), .ZN(new_n915));
  INV_X1    g0715(.A(G317), .ZN(new_n916));
  OAI221_X1 g0716(.A(new_n915), .B1(new_n458), .B2(new_n767), .C1(new_n916), .C2(new_n734), .ZN(new_n917));
  INV_X1    g0717(.A(G143), .ZN(new_n918));
  OAI221_X1 g0718(.A(new_n254), .B1(new_n229), .B2(new_n738), .C1(new_n808), .C2(new_n918), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n749), .A2(new_n421), .B1(new_n767), .B2(new_n230), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n735), .A2(G137), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n755), .A2(new_n208), .ZN(new_n922));
  NOR4_X1   g0722(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  OAI221_X1 g0723(.A(new_n923), .B1(new_n216), .B2(new_n757), .C1(new_n324), .C2(new_n742), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT47), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n238), .A2(new_n780), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n775), .B(new_n730), .C1(new_n682), .C2(new_n397), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n926), .A2(new_n730), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n728), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT106), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n479), .A2(new_n665), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n931), .B1(new_n632), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n487), .A2(KEYINPUT106), .A3(new_n932), .ZN(new_n935));
  INV_X1    g0735(.A(new_n630), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n934), .B(new_n935), .C1(new_n936), .C2(new_n932), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n929), .B(new_n930), .C1(new_n776), .C2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n670), .A2(new_n671), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n497), .A2(new_n665), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n618), .A2(new_n941), .ZN(new_n942));
  OR3_X1    g0742(.A1(new_n940), .A2(KEYINPUT42), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n678), .A2(new_n618), .A3(new_n941), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n634), .A2(new_n668), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT42), .B1(new_n940), .B2(new_n942), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n943), .A2(new_n944), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(KEYINPUT107), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(KEYINPUT107), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n953));
  INV_X1    g0753(.A(new_n951), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n948), .A2(new_n953), .A3(new_n949), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n634), .A2(new_n665), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n942), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n956), .B1(new_n677), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n677), .A2(new_n959), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n952), .A2(new_n961), .A3(new_n955), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n727), .A2(G1), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n679), .A2(new_n958), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT45), .Z(new_n967));
  NOR2_X1   g0767(.A1(new_n679), .A2(new_n958), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT44), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n677), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n672), .A2(new_n676), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n677), .A2(new_n940), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n974), .A2(new_n722), .A3(new_n699), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n976), .A2(new_n723), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n683), .B(KEYINPUT41), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n965), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n939), .B1(new_n963), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(G387));
  NAND2_X1  g0782(.A1(new_n752), .A2(new_n397), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n757), .B2(new_n230), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n295), .B(new_n984), .C1(G50), .C2(new_n795), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n745), .A2(G159), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n734), .A2(new_n421), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n738), .A2(new_n208), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(new_n741), .C2(new_n271), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n985), .A2(new_n912), .A3(new_n986), .A4(new_n989), .ZN(new_n990));
  AOI22_X1  g0790(.A1(G294), .A2(new_n769), .B1(new_n752), .B2(G283), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n737), .A2(new_n757), .B1(new_n749), .B2(new_n916), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT109), .Z(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(new_n756), .B2(new_n742), .C1(new_n747), .C2(new_n808), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT48), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n991), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT110), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n995), .B2(new_n994), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(KEYINPUT49), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n763), .A2(G116), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n735), .A2(G326), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n999), .A2(new_n295), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n998), .A2(KEYINPUT49), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n990), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n730), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n670), .A2(new_n776), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n685), .B(new_n445), .C1(new_n230), .C2(new_n208), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT108), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n271), .A2(new_n216), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT50), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n780), .B1(new_n1008), .B2(new_n1010), .C1(new_n242), .C2(new_n445), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(G107), .B2(new_n204), .C1(new_n685), .C2(new_n783), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n785), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1005), .A2(new_n930), .A3(new_n1006), .A4(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n683), .B1(new_n723), .B2(new_n974), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1014), .B1(new_n965), .B2(new_n973), .C1(new_n975), .C2(new_n1015), .ZN(G393));
  INV_X1    g0816(.A(new_n971), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n970), .A2(new_n677), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n683), .B(new_n976), .C1(new_n1019), .C2(new_n975), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n964), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n780), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n785), .B1(new_n457), .B2(new_n204), .C1(new_n249), .C2(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n808), .A2(new_n421), .B1(new_n749), .B2(new_n324), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT51), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n295), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n755), .A2(new_n210), .B1(new_n734), .B2(new_n918), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n757), .A2(new_n281), .B1(new_n219), .B2(new_n738), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(G77), .C2(new_n752), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1026), .B(new_n1029), .C1(new_n1025), .C2(new_n1024), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G50), .B2(new_n741), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n745), .A2(G317), .B1(new_n795), .B2(G311), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT52), .Z(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n295), .C1(new_n807), .C2(new_n757), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n738), .A2(new_n754), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n734), .A2(new_n747), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n764), .B1(new_n742), .B2(new_n737), .ZN(new_n1037));
  NOR4_X1   g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n752), .A2(G116), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1031), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n930), .B(new_n1023), .C1(new_n1040), .C2(new_n731), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT111), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1041), .A2(new_n1042), .B1(new_n775), .B2(new_n959), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1020), .A2(new_n1021), .A3(new_n1044), .ZN(G390));
  NAND4_X1  g0845(.A1(new_n721), .A2(new_n870), .A3(G330), .A4(new_n814), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n665), .B(new_n791), .C1(new_n696), .C2(new_n636), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n870), .B1(new_n1047), .B2(new_n859), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n822), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n883), .A3(new_n1049), .ZN(new_n1050));
  AND3_X1   g0850(.A1(new_n838), .A2(KEYINPUT39), .A3(new_n839), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT39), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1051), .B1(new_n883), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n822), .B1(new_n861), .B2(new_n870), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1046), .B(new_n1050), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n840), .B1(new_n854), .B2(KEYINPUT39), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n859), .B1(new_n690), .B2(new_n814), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n870), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1049), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n854), .A2(new_n822), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1056), .A2(new_n1059), .B1(new_n1060), .B2(new_n1048), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n880), .A2(new_n870), .A3(G330), .A4(new_n814), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1055), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n880), .A2(G330), .A3(new_n814), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n1058), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1047), .A2(new_n859), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n1046), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n721), .A2(G330), .A3(new_n814), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n881), .A2(G330), .B1(new_n1069), .B2(new_n1058), .ZN(new_n1070));
  OAI21_X1  g0870(.A(KEYINPUT112), .B1(new_n1070), .B2(new_n1057), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1058), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n1062), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT112), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(new_n1074), .A3(new_n861), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1068), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n890), .A2(new_n875), .A3(new_n654), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1063), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1074), .B1(new_n1073), .B2(new_n861), .ZN(new_n1079));
  AOI211_X1 g0879(.A(KEYINPUT112), .B(new_n1057), .C1(new_n1072), .C2(new_n1062), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1067), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1050), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1062), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1077), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1081), .A2(new_n1055), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1078), .A2(new_n1086), .A3(new_n683), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1063), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n295), .B1(new_n767), .B2(new_n208), .C1(new_n749), .C2(new_n579), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n741), .A2(G107), .B1(G87), .B2(new_n769), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n755), .A2(new_n230), .B1(new_n734), .B2(new_n807), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1090), .B(new_n1092), .C1(new_n754), .C2(new_n808), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1089), .B(new_n1093), .C1(G97), .C2(new_n759), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n735), .A2(G125), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n745), .A2(G128), .B1(G50), .B2(new_n763), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n752), .A2(G159), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n738), .A2(new_n421), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT53), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n741), .A2(G137), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n749), .A2(new_n802), .ZN(new_n1102));
  XOR2_X1   g0902(.A(KEYINPUT54), .B(G143), .Z(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n254), .B1(new_n757), .B2(new_n1104), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1101), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1094), .B1(new_n1095), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(new_n731), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n728), .B(new_n1108), .C1(new_n1056), .C2(new_n773), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n818), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n281), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1088), .A2(new_n964), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1087), .A2(new_n1112), .ZN(G378));
  XOR2_X1   g0913(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OR2_X1    g0915(.A1(new_n439), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n439), .A2(new_n1115), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1116), .A2(new_n1117), .B1(new_n424), .B2(new_n825), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n439), .A2(new_n1115), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n427), .B(new_n1114), .C1(new_n432), .C2(new_n438), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n424), .A2(new_n825), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n889), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1123), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n894), .A2(G330), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1124), .A2(new_n873), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1125), .B1(new_n894), .B2(G330), .ZN(new_n1128));
  INV_X1    g0928(.A(G330), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1129), .B(new_n1123), .C1(new_n892), .C2(new_n893), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n874), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(KEYINPUT117), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT117), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n873), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n964), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n745), .A2(G116), .B1(G58), .B2(new_n763), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1137), .B1(new_n754), .B2(new_n734), .C1(new_n398), .C2(new_n757), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G97), .B2(new_n741), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n749), .A2(new_n458), .ZN(new_n1140));
  NOR4_X1   g0940(.A1(new_n1140), .A2(new_n254), .A3(new_n261), .A4(new_n988), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1139), .B(new_n1141), .C1(new_n230), .C2(new_n767), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT58), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n216), .B1(G33), .B2(G41), .C1(new_n254), .C2(new_n261), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n745), .A2(G125), .B1(G150), .B2(new_n752), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT113), .ZN(new_n1146));
  INV_X1    g0946(.A(G128), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n749), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n741), .A2(G132), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n759), .A2(G137), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n769), .A2(new_n1103), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT59), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(G33), .A2(G41), .ZN(new_n1155));
  INV_X1    g0955(.A(G124), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1155), .B1(new_n734), .B2(new_n1156), .C1(new_n324), .C2(new_n755), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1143), .B(new_n1144), .C1(new_n1154), .C2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT114), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n731), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT115), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1123), .A2(new_n774), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n930), .B1(new_n818), .B2(G50), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT116), .Z(new_n1166));
  NOR3_X1   g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1136), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1085), .B1(new_n1076), .B2(new_n1063), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n684), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT118), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1175));
  AND4_X1   g0975(.A1(new_n1174), .A2(new_n1175), .A3(new_n1170), .A4(KEYINPUT57), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1172), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1174), .B1(new_n1177), .B2(new_n1170), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1169), .B1(new_n1173), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(G375));
  OAI21_X1  g0981(.A(KEYINPUT119), .B1(new_n1076), .B2(new_n965), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G159), .A2(new_n769), .B1(new_n752), .B2(G50), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n254), .C1(new_n742), .C2(new_n1104), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n808), .A2(new_n802), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n795), .A2(G137), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n763), .A2(G58), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n1147), .B2(new_n734), .C1(new_n757), .C2(new_n421), .ZN(new_n1188));
  NOR4_X1   g0988(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n983), .B1(new_n757), .B2(new_n458), .C1(new_n754), .C2(new_n749), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT120), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n295), .B1(new_n755), .B2(new_n208), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n745), .A2(G294), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n1191), .B2(new_n1192), .C1(new_n579), .C2(new_n742), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1190), .B(new_n1194), .C1(G97), .C2(new_n769), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n735), .A2(G303), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1189), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT121), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1198), .A2(new_n730), .B1(new_n230), .B2(new_n1110), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1199), .B(new_n930), .C1(new_n774), .C2(new_n870), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT119), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1081), .A2(new_n1201), .A3(new_n964), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1182), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1077), .B(new_n1067), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n978), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1204), .A2(new_n1207), .ZN(G381));
  INV_X1    g1008(.A(KEYINPUT123), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(G378), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1087), .A2(KEYINPUT123), .A3(new_n1112), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1180), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(G390), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n980), .A2(new_n960), .A3(new_n962), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1214), .A2(new_n1215), .A3(new_n938), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1216), .A2(G381), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT122), .Z(new_n1219));
  NAND3_X1  g1019(.A1(new_n1213), .A2(new_n1217), .A3(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT124), .ZN(G407));
  NAND2_X1  g1021(.A1(new_n1213), .A2(new_n664), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(G407), .A2(G213), .A3(new_n1222), .ZN(G409));
  NAND3_X1  g1023(.A1(new_n1076), .A2(KEYINPUT60), .A3(new_n1077), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT60), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1206), .A2(new_n1225), .ZN(new_n1226));
  AND4_X1   g1026(.A1(new_n683), .A2(new_n1224), .A3(new_n1226), .A4(new_n1205), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n794), .B(new_n819), .C1(new_n1227), .C2(new_n1203), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1224), .A2(new_n1226), .A3(new_n683), .A4(new_n1205), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1204), .A2(G384), .A3(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n660), .A2(G343), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(G2897), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1228), .A2(new_n1230), .A3(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1232), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1167), .B1(new_n1175), .B2(new_n964), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n978), .B(new_n1170), .C1(new_n1132), .C2(new_n1135), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1210), .A2(new_n1211), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1180), .B2(G378), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1235), .B1(new_n1239), .B2(new_n1231), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1169), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1170), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n873), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1128), .A2(new_n1130), .A3(new_n874), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1133), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1127), .A2(KEYINPUT117), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1242), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n683), .B1(new_n1247), .B2(KEYINPUT57), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1177), .A2(new_n1170), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(KEYINPUT118), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1177), .A2(new_n1174), .A3(new_n1170), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(G378), .B(new_n1241), .C1(new_n1248), .C2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1237), .A2(new_n1236), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1212), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1231), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1240), .A2(KEYINPUT63), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1231), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1260), .A2(KEYINPUT63), .A3(new_n1258), .A4(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT125), .B1(new_n981), .B2(new_n1214), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(G393), .B(G396), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1263), .B(new_n1264), .C1(new_n981), .C2(new_n1214), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1264), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT125), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1216), .A2(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n981), .A2(new_n1214), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1266), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1265), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1262), .A2(new_n1271), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1259), .A2(KEYINPUT61), .A3(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1260), .A2(new_n1261), .A3(new_n1258), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1274), .A2(KEYINPUT62), .B1(new_n1275), .B2(new_n1235), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1231), .B(new_n1257), .C1(new_n1253), .C2(new_n1255), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT61), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1271), .B1(new_n1276), .B2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT126), .B1(new_n1273), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1240), .A2(KEYINPUT63), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1274), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1272), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT126), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1265), .A2(new_n1270), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1240), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1285), .B1(new_n1274), .B2(KEYINPUT62), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1288), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1286), .A2(new_n1287), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1281), .A2(new_n1292), .ZN(G405));
  NAND2_X1  g1093(.A1(new_n1257), .A2(KEYINPUT127), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1288), .B(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G375), .A2(new_n1212), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1296), .B(new_n1253), .C1(KEYINPUT127), .C2(new_n1257), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(new_n1295), .B(new_n1297), .ZN(G402));
endmodule


