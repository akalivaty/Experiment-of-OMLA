

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740;

  INV_X1 U371 ( .A(G953), .ZN(n712) );
  NOR2_X2 U372 ( .A1(n592), .A2(n350), .ZN(n422) );
  XNOR2_X2 U373 ( .A(n488), .B(KEYINPUT33), .ZN(n673) );
  XNOR2_X2 U374 ( .A(n477), .B(n478), .ZN(n540) );
  NOR2_X1 U375 ( .A1(n653), .A2(n654), .ZN(n525) );
  XNOR2_X1 U376 ( .A(n462), .B(G472), .ZN(n554) );
  AND2_X1 U377 ( .A1(n678), .A2(n607), .ZN(n605) );
  XNOR2_X1 U378 ( .A(n509), .B(KEYINPUT35), .ZN(n734) );
  XNOR2_X1 U379 ( .A(n554), .B(KEYINPUT6), .ZN(n573) );
  XNOR2_X1 U380 ( .A(n695), .B(n424), .ZN(n696) );
  XNOR2_X1 U381 ( .A(n430), .B(n389), .ZN(n716) );
  XOR2_X1 U382 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n436) );
  XOR2_X1 U383 ( .A(KEYINPUT67), .B(G101), .Z(n456) );
  XNOR2_X2 U384 ( .A(n722), .B(n423), .ZN(n487) );
  XNOR2_X2 U385 ( .A(n372), .B(n395), .ZN(n722) );
  OR2_X1 U386 ( .A1(n689), .A2(G902), .ZN(n404) );
  INV_X1 U387 ( .A(KEYINPUT74), .ZN(n420) );
  XNOR2_X1 U388 ( .A(n497), .B(n370), .ZN(n372) );
  XNOR2_X1 U389 ( .A(n371), .B(G137), .ZN(n370) );
  INV_X1 U390 ( .A(KEYINPUT4), .ZN(n371) );
  XNOR2_X1 U391 ( .A(n438), .B(G125), .ZN(n467) );
  INV_X1 U392 ( .A(G146), .ZN(n438) );
  NAND2_X1 U393 ( .A1(n651), .A2(n553), .ZN(n576) );
  AND2_X1 U394 ( .A1(n630), .A2(n573), .ZN(n574) );
  XNOR2_X1 U395 ( .A(n445), .B(n357), .ZN(n580) );
  INV_X1 U396 ( .A(KEYINPUT19), .ZN(n357) );
  NOR2_X1 U397 ( .A1(G902), .A2(n611), .ZN(n462) );
  NOR2_X1 U398 ( .A1(G953), .A2(G237), .ZN(n500) );
  XNOR2_X1 U399 ( .A(n356), .B(n355), .ZN(n492) );
  INV_X1 U400 ( .A(KEYINPUT8), .ZN(n355) );
  NAND2_X1 U401 ( .A1(n712), .A2(G234), .ZN(n356) );
  XNOR2_X1 U402 ( .A(n467), .B(n419), .ZN(n721) );
  XNOR2_X1 U403 ( .A(G140), .B(KEYINPUT10), .ZN(n419) );
  XNOR2_X1 U404 ( .A(n392), .B(n716), .ZN(n686) );
  XNOR2_X1 U405 ( .A(n394), .B(n393), .ZN(n392) );
  XNOR2_X1 U406 ( .A(n433), .B(n434), .ZN(n393) );
  XNOR2_X1 U407 ( .A(n439), .B(n437), .ZN(n394) );
  XNOR2_X1 U408 ( .A(n366), .B(KEYINPUT39), .ZN(n601) );
  INV_X1 U409 ( .A(n641), .ZN(n373) );
  INV_X1 U410 ( .A(KEYINPUT1), .ZN(n403) );
  XNOR2_X1 U411 ( .A(n409), .B(KEYINPUT100), .ZN(n642) );
  NOR2_X1 U412 ( .A1(n630), .A2(n634), .ZN(n409) );
  NOR2_X1 U413 ( .A1(n740), .A2(n739), .ZN(n572) );
  XOR2_X1 U414 ( .A(KEYINPUT76), .B(KEYINPUT24), .Z(n469) );
  XNOR2_X1 U415 ( .A(n456), .B(G146), .ZN(n423) );
  XNOR2_X1 U416 ( .A(n458), .B(n415), .ZN(n414) );
  INV_X1 U417 ( .A(KEYINPUT94), .ZN(n415) );
  XNOR2_X1 U418 ( .A(n416), .B(n429), .ZN(n457) );
  XNOR2_X1 U419 ( .A(n428), .B(KEYINPUT3), .ZN(n416) );
  XNOR2_X1 U420 ( .A(G116), .B(G113), .ZN(n428) );
  INV_X1 U421 ( .A(KEYINPUT16), .ZN(n391) );
  XNOR2_X1 U422 ( .A(G104), .B(G110), .ZN(n426) );
  XNOR2_X1 U423 ( .A(G116), .B(G107), .ZN(n489) );
  XOR2_X1 U424 ( .A(KEYINPUT99), .B(G122), .Z(n490) );
  INV_X1 U425 ( .A(G134), .ZN(n454) );
  XOR2_X1 U426 ( .A(KEYINPUT98), .B(G104), .Z(n496) );
  XNOR2_X1 U427 ( .A(G143), .B(G113), .ZN(n495) );
  XNOR2_X1 U428 ( .A(G122), .B(KEYINPUT96), .ZN(n498) );
  NAND2_X1 U429 ( .A1(n379), .A2(n378), .ZN(n377) );
  INV_X1 U430 ( .A(n382), .ZN(n379) );
  AND2_X1 U431 ( .A1(n381), .A2(n380), .ZN(n376) );
  NAND2_X1 U432 ( .A1(n399), .A2(n585), .ZN(n398) );
  NAND2_X1 U433 ( .A1(n526), .A2(KEYINPUT34), .ZN(n399) );
  AND2_X1 U434 ( .A1(n573), .A2(n525), .ZN(n488) );
  XNOR2_X1 U435 ( .A(n516), .B(n515), .ZN(n534) );
  XNOR2_X1 U436 ( .A(n514), .B(KEYINPUT65), .ZN(n515) );
  AND2_X1 U437 ( .A1(n535), .A2(n388), .ZN(n387) );
  INV_X1 U438 ( .A(n573), .ZN(n388) );
  NAND2_X1 U439 ( .A1(n565), .A2(n566), .ZN(n374) );
  NOR2_X1 U440 ( .A1(n686), .A2(n607), .ZN(n443) );
  NOR2_X1 U441 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U442 ( .A(n507), .B(n506), .ZN(n521) );
  XOR2_X1 U443 ( .A(n494), .B(G478), .Z(n519) );
  NOR2_X1 U444 ( .A1(n699), .A2(G902), .ZN(n494) );
  XNOR2_X1 U445 ( .A(n363), .B(n418), .ZN(n706) );
  XNOR2_X1 U446 ( .A(n721), .B(n475), .ZN(n418) );
  XNOR2_X1 U447 ( .A(n472), .B(n476), .ZN(n363) );
  XNOR2_X1 U448 ( .A(n584), .B(KEYINPUT80), .ZN(n421) );
  INV_X1 U449 ( .A(KEYINPUT70), .ZN(n405) );
  INV_X1 U450 ( .A(KEYINPUT48), .ZN(n369) );
  XNOR2_X1 U451 ( .A(n510), .B(KEYINPUT101), .ZN(n640) );
  NOR2_X1 U452 ( .A1(n519), .A2(n521), .ZN(n510) );
  XOR2_X1 U453 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n499) );
  XNOR2_X1 U454 ( .A(KEYINPUT4), .B(KEYINPUT83), .ZN(n435) );
  XNOR2_X1 U455 ( .A(n432), .B(KEYINPUT84), .ZN(n433) );
  NAND2_X1 U456 ( .A1(G224), .A2(n712), .ZN(n432) );
  NAND2_X1 U457 ( .A1(G234), .A2(G237), .ZN(n446) );
  XOR2_X1 U458 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n447) );
  NOR2_X1 U459 ( .A1(n531), .A2(n530), .ZN(n532) );
  OR2_X1 U460 ( .A1(n576), .A2(n383), .ZN(n382) );
  XNOR2_X1 U461 ( .A(KEYINPUT66), .B(KEYINPUT0), .ZN(n452) );
  NOR2_X1 U462 ( .A1(n580), .A2(n451), .ZN(n453) );
  XNOR2_X1 U463 ( .A(G137), .B(G128), .ZN(n474) );
  XOR2_X1 U464 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n470) );
  XNOR2_X1 U465 ( .A(G119), .B(G110), .ZN(n468) );
  XNOR2_X1 U466 ( .A(n486), .B(n487), .ZN(n689) );
  NAND2_X1 U467 ( .A1(n540), .A2(n417), .ZN(n653) );
  INV_X1 U468 ( .A(n650), .ZN(n417) );
  XNOR2_X1 U469 ( .A(n487), .B(n461), .ZN(n611) );
  XNOR2_X1 U470 ( .A(n457), .B(n414), .ZN(n459) );
  XNOR2_X1 U471 ( .A(n481), .B(n390), .ZN(n389) );
  XNOR2_X1 U472 ( .A(n427), .B(n391), .ZN(n390) );
  XNOR2_X1 U473 ( .A(n412), .B(n493), .ZN(n699) );
  XNOR2_X1 U474 ( .A(n503), .B(n364), .ZN(n695) );
  XNOR2_X1 U475 ( .A(n504), .B(n505), .ZN(n364) );
  AND2_X1 U476 ( .A1(n601), .A2(n630), .ZN(n571) );
  AND2_X1 U477 ( .A1(n375), .A2(n384), .ZN(n578) );
  INV_X1 U478 ( .A(n654), .ZN(n384) );
  NOR2_X1 U479 ( .A1(n400), .A2(n398), .ZN(n397) );
  XNOR2_X1 U480 ( .A(n386), .B(n385), .ZN(n536) );
  INV_X1 U481 ( .A(KEYINPUT32), .ZN(n385) );
  INV_X1 U482 ( .A(n519), .ZN(n520) );
  NAND2_X1 U483 ( .A1(n374), .A2(n570), .ZN(n587) );
  INV_X1 U484 ( .A(n521), .ZN(n411) );
  XNOR2_X1 U485 ( .A(n537), .B(n359), .ZN(n358) );
  INV_X1 U486 ( .A(KEYINPUT104), .ZN(n359) );
  XNOR2_X1 U487 ( .A(n704), .B(n367), .ZN(n707) );
  XNOR2_X1 U488 ( .A(n706), .B(n705), .ZN(n367) );
  INV_X1 U489 ( .A(KEYINPUT56), .ZN(n361) );
  XNOR2_X1 U490 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n349) );
  AND2_X1 U491 ( .A1(n642), .A2(KEYINPUT47), .ZN(n350) );
  AND2_X1 U492 ( .A1(n570), .A2(n373), .ZN(n351) );
  OR2_X1 U493 ( .A1(n575), .A2(n377), .ZN(n352) );
  INV_X1 U494 ( .A(KEYINPUT34), .ZN(n402) );
  XOR2_X1 U495 ( .A(n686), .B(n685), .Z(n353) );
  XOR2_X1 U496 ( .A(n611), .B(KEYINPUT62), .Z(n354) );
  INV_X1 U497 ( .A(n410), .ZN(n634) );
  NAND2_X1 U498 ( .A1(n519), .A2(n411), .ZN(n410) );
  NAND2_X1 U499 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U500 ( .A1(n673), .A2(n401), .ZN(n400) );
  NAND2_X1 U501 ( .A1(n397), .A2(n396), .ZN(n509) );
  NAND2_X1 U502 ( .A1(n358), .A2(n538), .ZN(n539) );
  XNOR2_X1 U503 ( .A(n365), .B(n369), .ZN(n604) );
  NAND2_X1 U504 ( .A1(n360), .A2(n613), .ZN(n614) );
  XNOR2_X1 U505 ( .A(n612), .B(n354), .ZN(n360) );
  XNOR2_X1 U506 ( .A(n362), .B(n361), .ZN(G51) );
  NAND2_X1 U507 ( .A1(n688), .A2(n613), .ZN(n362) );
  NOR2_X1 U508 ( .A1(n650), .A2(n640), .ZN(n511) );
  NAND2_X1 U509 ( .A1(n595), .A2(n594), .ZN(n365) );
  NOR2_X2 U510 ( .A1(n724), .A2(KEYINPUT2), .ZN(n679) );
  NAND2_X1 U511 ( .A1(n351), .A2(n374), .ZN(n366) );
  NAND2_X1 U512 ( .A1(n534), .A2(n654), .ZN(n537) );
  XNOR2_X1 U513 ( .A(n491), .B(n349), .ZN(n413) );
  NOR2_X1 U514 ( .A1(n554), .A2(n576), .ZN(n556) );
  XNOR2_X1 U515 ( .A(n368), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U516 ( .A1(n698), .A2(n708), .ZN(n368) );
  XNOR2_X2 U517 ( .A(n455), .B(n454), .ZN(n395) );
  XNOR2_X2 U518 ( .A(n431), .B(G128), .ZN(n455) );
  NAND2_X1 U519 ( .A1(n352), .A2(n376), .ZN(n375) );
  INV_X1 U520 ( .A(n577), .ZN(n378) );
  NAND2_X1 U521 ( .A1(n382), .A2(n577), .ZN(n380) );
  NAND2_X1 U522 ( .A1(n575), .A2(n577), .ZN(n381) );
  NOR2_X1 U523 ( .A1(n575), .A2(n576), .ZN(n596) );
  INV_X1 U524 ( .A(n599), .ZN(n383) );
  NAND2_X1 U525 ( .A1(n534), .A2(n387), .ZN(n386) );
  XNOR2_X1 U526 ( .A(n413), .B(n395), .ZN(n412) );
  NAND2_X1 U527 ( .A1(n673), .A2(KEYINPUT34), .ZN(n396) );
  NAND2_X1 U528 ( .A1(n512), .A2(n402), .ZN(n401) );
  XNOR2_X2 U529 ( .A(n557), .B(n403), .ZN(n654) );
  XNOR2_X2 U530 ( .A(n404), .B(G469), .ZN(n557) );
  XNOR2_X1 U531 ( .A(n406), .B(n405), .ZN(n594) );
  NOR2_X1 U532 ( .A1(n622), .A2(n642), .ZN(n590) );
  XNOR2_X1 U533 ( .A(n408), .B(n420), .ZN(n407) );
  NAND2_X1 U534 ( .A1(n407), .A2(n593), .ZN(n406) );
  XNOR2_X1 U535 ( .A(n501), .B(n425), .ZN(n502) );
  NAND2_X1 U536 ( .A1(n422), .A2(n421), .ZN(n408) );
  INV_X1 U537 ( .A(n540), .ZN(n651) );
  NAND2_X1 U538 ( .A1(n605), .A2(n679), .ZN(n610) );
  XNOR2_X2 U539 ( .A(n606), .B(KEYINPUT81), .ZN(n724) );
  XNOR2_X1 U540 ( .A(KEYINPUT119), .B(KEYINPUT59), .ZN(n424) );
  AND2_X1 U541 ( .A1(G214), .A2(n500), .ZN(n425) );
  NOR2_X1 U542 ( .A1(G952), .A2(n712), .ZN(n708) );
  INV_X1 U543 ( .A(n640), .ZN(n644) );
  INV_X1 U544 ( .A(KEYINPUT44), .ZN(n541) );
  INV_X1 U545 ( .A(n637), .ZN(n602) );
  NOR2_X1 U546 ( .A1(n638), .A2(n602), .ZN(n603) );
  XNOR2_X1 U547 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U548 ( .A(n453), .B(n452), .ZN(n512) );
  XNOR2_X1 U549 ( .A(n474), .B(n473), .ZN(n475) );
  INV_X1 U550 ( .A(n708), .ZN(n613) );
  XNOR2_X1 U551 ( .A(n697), .B(n696), .ZN(n698) );
  XOR2_X1 U552 ( .A(KEYINPUT73), .B(G122), .Z(n427) );
  XNOR2_X1 U553 ( .A(n426), .B(G107), .ZN(n481) );
  XOR2_X1 U554 ( .A(KEYINPUT71), .B(G119), .Z(n429) );
  INV_X1 U555 ( .A(n457), .ZN(n430) );
  XNOR2_X2 U556 ( .A(G143), .B(KEYINPUT79), .ZN(n431) );
  INV_X1 U557 ( .A(n455), .ZN(n434) );
  XOR2_X1 U558 ( .A(n436), .B(n435), .Z(n437) );
  XNOR2_X1 U559 ( .A(n467), .B(n456), .ZN(n439) );
  XNOR2_X1 U560 ( .A(G902), .B(KEYINPUT15), .ZN(n463) );
  INV_X1 U561 ( .A(n463), .ZN(n607) );
  XOR2_X1 U562 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n441) );
  OR2_X1 U563 ( .A1(G237), .A2(G902), .ZN(n444) );
  NAND2_X1 U564 ( .A1(G210), .A2(n444), .ZN(n440) );
  XNOR2_X1 U565 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X2 U566 ( .A(n443), .B(n442), .ZN(n599) );
  NAND2_X1 U567 ( .A1(G214), .A2(n444), .ZN(n639) );
  NAND2_X1 U568 ( .A1(n599), .A2(n639), .ZN(n445) );
  XNOR2_X1 U569 ( .A(n447), .B(n446), .ZN(n448) );
  NAND2_X1 U570 ( .A1(G952), .A2(n448), .ZN(n671) );
  NOR2_X1 U571 ( .A1(G953), .A2(n671), .ZN(n552) );
  NAND2_X1 U572 ( .A1(n448), .A2(G902), .ZN(n449) );
  XOR2_X1 U573 ( .A(n449), .B(KEYINPUT89), .Z(n549) );
  XOR2_X1 U574 ( .A(G898), .B(KEYINPUT88), .Z(n711) );
  NAND2_X1 U575 ( .A1(G953), .A2(n711), .ZN(n717) );
  NOR2_X1 U576 ( .A1(n549), .A2(n717), .ZN(n450) );
  NOR2_X1 U577 ( .A1(n552), .A2(n450), .ZN(n451) );
  INV_X1 U578 ( .A(n512), .ZN(n526) );
  XOR2_X1 U579 ( .A(KEYINPUT69), .B(G131), .Z(n497) );
  NAND2_X1 U580 ( .A1(n500), .A2(G210), .ZN(n460) );
  XOR2_X1 U581 ( .A(KEYINPUT5), .B(KEYINPUT75), .Z(n458) );
  XNOR2_X1 U582 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U583 ( .A(KEYINPUT25), .B(KEYINPUT93), .Z(n466) );
  NAND2_X1 U584 ( .A1(G234), .A2(n463), .ZN(n464) );
  XNOR2_X1 U585 ( .A(KEYINPUT20), .B(n464), .ZN(n479) );
  NAND2_X1 U586 ( .A1(n479), .A2(G217), .ZN(n465) );
  XNOR2_X1 U587 ( .A(n466), .B(n465), .ZN(n478) );
  XNOR2_X1 U588 ( .A(n469), .B(n468), .ZN(n471) );
  INV_X1 U589 ( .A(KEYINPUT23), .ZN(n473) );
  AND2_X1 U590 ( .A1(n492), .A2(G221), .ZN(n476) );
  NOR2_X1 U591 ( .A1(G902), .A2(n706), .ZN(n477) );
  NAND2_X1 U592 ( .A1(n479), .A2(G221), .ZN(n480) );
  XNOR2_X1 U593 ( .A(n480), .B(KEYINPUT21), .ZN(n650) );
  XNOR2_X1 U594 ( .A(G140), .B(KEYINPUT90), .ZN(n485) );
  XOR2_X1 U595 ( .A(n481), .B(KEYINPUT77), .Z(n483) );
  NAND2_X1 U596 ( .A1(G227), .A2(n712), .ZN(n482) );
  XNOR2_X1 U597 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U598 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U599 ( .A(n490), .B(n489), .ZN(n491) );
  NAND2_X1 U600 ( .A1(G217), .A2(n492), .ZN(n493) );
  XNOR2_X1 U601 ( .A(n496), .B(n495), .ZN(n505) );
  XNOR2_X1 U602 ( .A(n497), .B(KEYINPUT12), .ZN(n504) );
  XNOR2_X1 U603 ( .A(n499), .B(n498), .ZN(n501) );
  XNOR2_X1 U604 ( .A(n721), .B(n502), .ZN(n503) );
  NOR2_X1 U605 ( .A1(G902), .A2(n695), .ZN(n507) );
  XNOR2_X1 U606 ( .A(KEYINPUT13), .B(G475), .ZN(n506) );
  NAND2_X1 U607 ( .A1(n519), .A2(n521), .ZN(n508) );
  XNOR2_X1 U608 ( .A(KEYINPUT105), .B(n508), .ZN(n585) );
  NAND2_X1 U609 ( .A1(n734), .A2(KEYINPUT44), .ZN(n518) );
  XNOR2_X1 U610 ( .A(n511), .B(KEYINPUT102), .ZN(n513) );
  NAND2_X1 U611 ( .A1(n513), .A2(n512), .ZN(n516) );
  XNOR2_X1 U612 ( .A(KEYINPUT72), .B(KEYINPUT22), .ZN(n514) );
  NOR2_X1 U613 ( .A1(n573), .A2(n537), .ZN(n517) );
  NAND2_X1 U614 ( .A1(n517), .A2(n540), .ZN(n615) );
  NAND2_X1 U615 ( .A1(n518), .A2(n615), .ZN(n531) );
  NAND2_X1 U616 ( .A1(n521), .A2(n520), .ZN(n628) );
  INV_X1 U617 ( .A(n628), .ZN(n630) );
  INV_X1 U618 ( .A(n557), .ZN(n569) );
  NOR2_X1 U619 ( .A1(n653), .A2(n526), .ZN(n523) );
  INV_X1 U620 ( .A(n554), .ZN(n560) );
  BUF_X1 U621 ( .A(n560), .Z(n522) );
  INV_X1 U622 ( .A(n522), .ZN(n538) );
  NAND2_X1 U623 ( .A1(n523), .A2(n538), .ZN(n524) );
  NOR2_X1 U624 ( .A1(n569), .A2(n524), .ZN(n617) );
  NAND2_X1 U625 ( .A1(n522), .A2(n525), .ZN(n662) );
  NOR2_X1 U626 ( .A1(n526), .A2(n662), .ZN(n528) );
  XNOR2_X1 U627 ( .A(KEYINPUT95), .B(KEYINPUT31), .ZN(n527) );
  XNOR2_X1 U628 ( .A(n528), .B(n527), .ZN(n635) );
  NOR2_X1 U629 ( .A1(n617), .A2(n635), .ZN(n529) );
  NOR2_X1 U630 ( .A1(n642), .A2(n529), .ZN(n530) );
  XNOR2_X1 U631 ( .A(n532), .B(KEYINPUT82), .ZN(n546) );
  OR2_X1 U632 ( .A1(n540), .A2(n654), .ZN(n533) );
  XNOR2_X1 U633 ( .A(KEYINPUT103), .B(n533), .ZN(n535) );
  XNOR2_X1 U634 ( .A(n536), .B(KEYINPUT64), .ZN(n736) );
  NOR2_X1 U635 ( .A1(n540), .A2(n539), .ZN(n621) );
  NOR2_X1 U636 ( .A1(n736), .A2(n621), .ZN(n542) );
  XNOR2_X1 U637 ( .A(n542), .B(n541), .ZN(n544) );
  NAND2_X1 U638 ( .A1(n542), .A2(n734), .ZN(n543) );
  NAND2_X1 U639 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X2 U640 ( .A(n547), .B(KEYINPUT45), .ZN(n678) );
  XNOR2_X1 U641 ( .A(KEYINPUT38), .B(n599), .ZN(n641) );
  NOR2_X1 U642 ( .A1(n641), .A2(n640), .ZN(n648) );
  NAND2_X1 U643 ( .A1(n639), .A2(n648), .ZN(n548) );
  XOR2_X1 U644 ( .A(KEYINPUT41), .B(n548), .Z(n672) );
  OR2_X1 U645 ( .A1(n712), .A2(n549), .ZN(n550) );
  NOR2_X1 U646 ( .A1(G900), .A2(n550), .ZN(n551) );
  NOR2_X1 U647 ( .A1(n552), .A2(n551), .ZN(n567) );
  NOR2_X1 U648 ( .A1(n567), .A2(n650), .ZN(n553) );
  XNOR2_X1 U649 ( .A(KEYINPUT108), .B(KEYINPUT28), .ZN(n555) );
  XNOR2_X1 U650 ( .A(n556), .B(n555), .ZN(n558) );
  NAND2_X1 U651 ( .A1(n558), .A2(n557), .ZN(n579) );
  NOR2_X1 U652 ( .A1(n672), .A2(n579), .ZN(n559) );
  XNOR2_X1 U653 ( .A(n559), .B(KEYINPUT42), .ZN(n740) );
  NAND2_X1 U654 ( .A1(n560), .A2(n639), .ZN(n561) );
  XNOR2_X1 U655 ( .A(n561), .B(KEYINPUT30), .ZN(n562) );
  NAND2_X1 U656 ( .A1(KEYINPUT107), .A2(n562), .ZN(n566) );
  INV_X1 U657 ( .A(KEYINPUT107), .ZN(n564) );
  INV_X1 U658 ( .A(n562), .ZN(n563) );
  NAND2_X1 U659 ( .A1(n564), .A2(n563), .ZN(n565) );
  OR2_X1 U660 ( .A1(n653), .A2(n567), .ZN(n568) );
  XNOR2_X1 U661 ( .A(n571), .B(KEYINPUT40), .ZN(n739) );
  XNOR2_X1 U662 ( .A(n572), .B(KEYINPUT46), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n574), .A2(n639), .ZN(n575) );
  XNOR2_X1 U664 ( .A(KEYINPUT109), .B(KEYINPUT36), .ZN(n577) );
  XNOR2_X1 U665 ( .A(n578), .B(KEYINPUT110), .ZN(n737) );
  INV_X1 U666 ( .A(n737), .ZN(n593) );
  INV_X1 U667 ( .A(n579), .ZN(n582) );
  INV_X1 U668 ( .A(n580), .ZN(n581) );
  NAND2_X1 U669 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X2 U670 ( .A(n583), .B(KEYINPUT78), .ZN(n622) );
  NAND2_X1 U671 ( .A1(n622), .A2(KEYINPUT47), .ZN(n584) );
  INV_X1 U672 ( .A(n585), .ZN(n586) );
  NOR2_X1 U673 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U674 ( .A1(n588), .A2(n599), .ZN(n627) );
  XOR2_X1 U675 ( .A(KEYINPUT47), .B(KEYINPUT68), .Z(n589) );
  NAND2_X1 U676 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U677 ( .A1(n627), .A2(n591), .ZN(n592) );
  XOR2_X1 U678 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n598) );
  NAND2_X1 U679 ( .A1(n596), .A2(n654), .ZN(n597) );
  XNOR2_X1 U680 ( .A(n598), .B(n597), .ZN(n600) );
  NOR2_X1 U681 ( .A1(n600), .A2(n599), .ZN(n638) );
  NAND2_X1 U682 ( .A1(n634), .A2(n601), .ZN(n637) );
  AND2_X2 U683 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n606), .A2(n678), .ZN(n677) );
  AND2_X1 U685 ( .A1(KEYINPUT2), .A2(n607), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n677), .A2(n608), .ZN(n609) );
  NAND2_X2 U687 ( .A1(n610), .A2(n609), .ZN(n703) );
  NAND2_X1 U688 ( .A1(n703), .A2(G472), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n614), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U690 ( .A(G101), .B(n615), .ZN(G3) );
  NAND2_X1 U691 ( .A1(n617), .A2(n630), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n616), .B(G104), .ZN(G6) );
  XOR2_X1 U693 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n619) );
  NAND2_X1 U694 ( .A1(n617), .A2(n634), .ZN(n618) );
  XNOR2_X1 U695 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U696 ( .A(G107), .B(n620), .ZN(G9) );
  XOR2_X1 U697 ( .A(n621), .B(G110), .Z(G12) );
  BUF_X1 U698 ( .A(n622), .Z(n623) );
  NOR2_X1 U699 ( .A1(n623), .A2(n410), .ZN(n625) );
  XNOR2_X1 U700 ( .A(G128), .B(KEYINPUT29), .ZN(n624) );
  XNOR2_X1 U701 ( .A(n625), .B(n624), .ZN(G30) );
  XOR2_X1 U702 ( .A(G143), .B(KEYINPUT111), .Z(n626) );
  XNOR2_X1 U703 ( .A(n627), .B(n626), .ZN(G45) );
  NOR2_X1 U704 ( .A1(n623), .A2(n628), .ZN(n629) );
  XOR2_X1 U705 ( .A(G146), .B(n629), .Z(G48) );
  XOR2_X1 U706 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n632) );
  NAND2_X1 U707 ( .A1(n635), .A2(n630), .ZN(n631) );
  XNOR2_X1 U708 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U709 ( .A(G113), .B(n633), .ZN(G15) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n636), .B(G116), .ZN(G18) );
  XNOR2_X1 U712 ( .A(G134), .B(n637), .ZN(G36) );
  XOR2_X1 U713 ( .A(G140), .B(n638), .Z(G42) );
  INV_X1 U714 ( .A(n639), .ZN(n646) );
  NOR2_X1 U715 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U717 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U718 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U719 ( .A1(n673), .A2(n649), .ZN(n667) );
  NAND2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U721 ( .A(KEYINPUT49), .B(n652), .Z(n660) );
  XOR2_X1 U722 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n656) );
  NAND2_X1 U723 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U724 ( .A(n656), .B(n655), .ZN(n657) );
  XOR2_X1 U725 ( .A(KEYINPUT114), .B(n657), .Z(n658) );
  NOR2_X1 U726 ( .A1(n658), .A2(n522), .ZN(n659) );
  NAND2_X1 U727 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U729 ( .A(KEYINPUT51), .B(n663), .ZN(n664) );
  NOR2_X1 U730 ( .A1(n672), .A2(n664), .ZN(n665) );
  XNOR2_X1 U731 ( .A(n665), .B(KEYINPUT116), .ZN(n666) );
  NOR2_X1 U732 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U733 ( .A(n668), .B(KEYINPUT52), .Z(n669) );
  XNOR2_X1 U734 ( .A(KEYINPUT117), .B(n669), .ZN(n670) );
  NOR2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n675) );
  NOR2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U738 ( .A1(n676), .A2(n712), .ZN(n683) );
  NAND2_X1 U739 ( .A1(n677), .A2(KEYINPUT2), .ZN(n681) );
  NAND2_X1 U740 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U741 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U742 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U743 ( .A(n684), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U744 ( .A1(n703), .A2(G210), .ZN(n687) );
  XOR2_X1 U745 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n685) );
  XNOR2_X1 U746 ( .A(n687), .B(n353), .ZN(n688) );
  XNOR2_X1 U747 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n691) );
  XNOR2_X1 U748 ( .A(n689), .B(KEYINPUT57), .ZN(n690) );
  XNOR2_X1 U749 ( .A(n691), .B(n690), .ZN(n693) );
  NAND2_X1 U750 ( .A1(n703), .A2(G469), .ZN(n692) );
  XOR2_X1 U751 ( .A(n693), .B(n692), .Z(n694) );
  NOR2_X1 U752 ( .A1(n708), .A2(n694), .ZN(G54) );
  NAND2_X1 U753 ( .A1(n703), .A2(G475), .ZN(n697) );
  XNOR2_X1 U754 ( .A(n699), .B(KEYINPUT120), .ZN(n701) );
  NAND2_X1 U755 ( .A1(G478), .A2(n703), .ZN(n700) );
  XNOR2_X1 U756 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U757 ( .A1(n708), .A2(n702), .ZN(G63) );
  XOR2_X1 U758 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n705) );
  NAND2_X1 U759 ( .A1(n703), .A2(G217), .ZN(n704) );
  NOR2_X1 U760 ( .A1(n708), .A2(n707), .ZN(G66) );
  NAND2_X1 U761 ( .A1(G953), .A2(G224), .ZN(n709) );
  XOR2_X1 U762 ( .A(KEYINPUT61), .B(n709), .Z(n710) );
  NOR2_X1 U763 ( .A1(n711), .A2(n710), .ZN(n714) );
  AND2_X1 U764 ( .A1(n712), .A2(n678), .ZN(n713) );
  NOR2_X1 U765 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U766 ( .A(n715), .B(KEYINPUT123), .Z(n720) );
  XOR2_X1 U767 ( .A(G101), .B(n716), .Z(n718) );
  NAND2_X1 U768 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U769 ( .A(n720), .B(n719), .ZN(G69) );
  XOR2_X1 U770 ( .A(n722), .B(n721), .Z(n723) );
  XOR2_X1 U771 ( .A(KEYINPUT124), .B(n723), .Z(n728) );
  INV_X1 U772 ( .A(n728), .ZN(n725) );
  XOR2_X1 U773 ( .A(n725), .B(n724), .Z(n726) );
  NOR2_X1 U774 ( .A1(G953), .A2(n726), .ZN(n727) );
  XNOR2_X1 U775 ( .A(KEYINPUT125), .B(n727), .ZN(n733) );
  XOR2_X1 U776 ( .A(G227), .B(n728), .Z(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(G900), .ZN(n730) );
  XNOR2_X1 U778 ( .A(KEYINPUT126), .B(n730), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n731), .A2(G953), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n733), .A2(n732), .ZN(G72) );
  XNOR2_X1 U781 ( .A(n734), .B(G122), .ZN(n735) );
  XNOR2_X1 U782 ( .A(n735), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U783 ( .A(G119), .B(n736), .Z(G21) );
  XNOR2_X1 U784 ( .A(G125), .B(KEYINPUT37), .ZN(n738) );
  XNOR2_X1 U785 ( .A(n738), .B(n737), .ZN(G27) );
  XOR2_X1 U786 ( .A(n739), .B(G131), .Z(G33) );
  XOR2_X1 U787 ( .A(G137), .B(n740), .Z(G39) );
endmodule

