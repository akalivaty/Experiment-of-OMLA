

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739;

  INV_X1 U372 ( .A(n659), .ZN(n397) );
  OR2_X1 U373 ( .A1(n703), .A2(G902), .ZN(n394) );
  NOR2_X1 U374 ( .A1(n681), .A2(n715), .ZN(n676) );
  XOR2_X2 U375 ( .A(n470), .B(n469), .Z(n721) );
  OR2_X2 U376 ( .A1(n604), .A2(G902), .ZN(n386) );
  AND2_X2 U377 ( .A1(n516), .A2(n387), .ZN(n520) );
  AND2_X2 U378 ( .A1(n539), .A2(n554), .ZN(n540) );
  XNOR2_X2 U379 ( .A(n452), .B(n451), .ZN(n549) );
  AND2_X2 U380 ( .A1(n610), .A2(n596), .ZN(n452) );
  AND2_X2 U381 ( .A1(n603), .A2(n602), .ZN(n418) );
  NAND2_X1 U382 ( .A1(n365), .A2(n359), .ZN(n603) );
  INV_X1 U383 ( .A(n676), .ZN(n602) );
  NOR2_X1 U384 ( .A1(n586), .A2(n569), .ZN(n627) );
  OR2_X2 U385 ( .A1(n377), .A2(n373), .ZN(n581) );
  XNOR2_X1 U386 ( .A(n519), .B(n518), .ZN(n559) );
  XNOR2_X1 U387 ( .A(n481), .B(n355), .ZN(n393) );
  XNOR2_X1 U388 ( .A(n434), .B(G128), .ZN(n447) );
  OR2_X1 U389 ( .A1(n572), .A2(n397), .ZN(n586) );
  XNOR2_X1 U390 ( .A(n372), .B(n371), .ZN(n592) );
  INV_X1 U391 ( .A(KEYINPUT44), .ZN(n371) );
  NAND2_X1 U392 ( .A1(n353), .A2(n370), .ZN(n372) );
  XNOR2_X1 U393 ( .A(n722), .B(G146), .ZN(n495) );
  XNOR2_X1 U394 ( .A(n447), .B(KEYINPUT4), .ZN(n460) );
  XNOR2_X1 U395 ( .A(n431), .B(G475), .ZN(n529) );
  XNOR2_X1 U396 ( .A(n662), .B(KEYINPUT6), .ZN(n396) );
  AND2_X1 U397 ( .A1(n404), .A2(n526), .ZN(n368) );
  XOR2_X1 U398 ( .A(G137), .B(G140), .Z(n469) );
  XOR2_X1 U399 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n443) );
  XNOR2_X1 U400 ( .A(G902), .B(KEYINPUT15), .ZN(n596) );
  INV_X1 U401 ( .A(n529), .ZN(n453) );
  INV_X1 U402 ( .A(KEYINPUT0), .ZN(n375) );
  NAND2_X1 U403 ( .A1(n558), .A2(KEYINPUT0), .ZN(n378) );
  XNOR2_X1 U404 ( .A(n495), .B(n412), .ZN(n604) );
  XNOR2_X1 U405 ( .A(n413), .B(n492), .ZN(n412) );
  XNOR2_X1 U406 ( .A(n496), .B(n414), .ZN(n413) );
  NOR2_X1 U407 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U408 ( .A(n441), .B(n352), .ZN(n380) );
  XNOR2_X1 U409 ( .A(n442), .B(n382), .ZN(n381) );
  XNOR2_X1 U410 ( .A(n493), .B(KEYINPUT16), .ZN(n382) );
  INV_X1 U411 ( .A(G143), .ZN(n434) );
  XNOR2_X1 U412 ( .A(n436), .B(n354), .ZN(n369) );
  XNOR2_X1 U413 ( .A(G134), .B(G122), .ZN(n432) );
  XNOR2_X1 U414 ( .A(KEYINPUT41), .B(n532), .ZN(n668) );
  NOR2_X1 U415 ( .A1(n634), .A2(n530), .ZN(n409) );
  XNOR2_X1 U416 ( .A(n360), .B(KEYINPUT34), .ZN(n561) );
  NOR2_X1 U417 ( .A1(n653), .A2(n581), .ZN(n360) );
  NOR2_X1 U418 ( .A1(n581), .A2(n566), .ZN(n568) );
  XNOR2_X1 U419 ( .A(n468), .B(n467), .ZN(n515) );
  NAND2_X1 U420 ( .A1(n517), .A2(n646), .ZN(n519) );
  INV_X1 U421 ( .A(n396), .ZN(n587) );
  INV_X1 U422 ( .A(G953), .ZN(n730) );
  NOR2_X1 U423 ( .A1(G952), .A2(n730), .ZN(n707) );
  INV_X1 U424 ( .A(KEYINPUT66), .ZN(n392) );
  AND2_X1 U425 ( .A1(n632), .A2(KEYINPUT78), .ZN(n362) );
  AND2_X1 U426 ( .A1(n527), .A2(n368), .ZN(n403) );
  XNOR2_X1 U427 ( .A(n494), .B(KEYINPUT5), .ZN(n414) );
  XNOR2_X1 U428 ( .A(G101), .B(G113), .ZN(n487) );
  XOR2_X1 U429 ( .A(G137), .B(G116), .Z(n488) );
  XNOR2_X1 U430 ( .A(n460), .B(n461), .ZN(n722) );
  XNOR2_X1 U431 ( .A(G131), .B(G134), .ZN(n461) );
  INV_X1 U432 ( .A(n618), .ZN(n589) );
  XNOR2_X1 U433 ( .A(G119), .B(KEYINPUT3), .ZN(n493) );
  NOR2_X1 U434 ( .A1(G953), .A2(G237), .ZN(n489) );
  XOR2_X1 U435 ( .A(G107), .B(G104), .Z(n462) );
  NAND2_X1 U436 ( .A1(G234), .A2(G237), .ZN(n454) );
  XOR2_X1 U437 ( .A(KEYINPUT14), .B(KEYINPUT86), .Z(n455) );
  NOR2_X1 U438 ( .A1(G902), .A2(G237), .ZN(n450) );
  XNOR2_X1 U439 ( .A(n363), .B(n472), .ZN(n476) );
  XNOR2_X1 U440 ( .A(n471), .B(n364), .ZN(n363) );
  INV_X1 U441 ( .A(KEYINPUT91), .ZN(n364) );
  XNOR2_X1 U442 ( .A(G128), .B(KEYINPUT23), .ZN(n473) );
  XOR2_X1 U443 ( .A(KEYINPUT89), .B(KEYINPUT24), .Z(n474) );
  XOR2_X1 U444 ( .A(G140), .B(G131), .Z(n420) );
  INV_X1 U445 ( .A(KEYINPUT10), .ZN(n425) );
  XNOR2_X1 U446 ( .A(G113), .B(G104), .ZN(n426) );
  XNOR2_X1 U447 ( .A(G143), .B(KEYINPUT12), .ZN(n421) );
  XOR2_X1 U448 ( .A(KEYINPUT11), .B(KEYINPUT98), .Z(n422) );
  INV_X1 U449 ( .A(n596), .ZN(n408) );
  XNOR2_X1 U450 ( .A(n495), .B(n398), .ZN(n687) );
  XNOR2_X1 U451 ( .A(n466), .B(n399), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U453 ( .A(n463), .B(n352), .ZN(n399) );
  XNOR2_X1 U454 ( .A(n405), .B(n708), .ZN(n610) );
  XNOR2_X1 U455 ( .A(n449), .B(n406), .ZN(n405) );
  XNOR2_X1 U456 ( .A(n445), .B(n446), .ZN(n406) );
  XNOR2_X1 U457 ( .A(n384), .B(n383), .ZN(n653) );
  INV_X1 U458 ( .A(KEYINPUT33), .ZN(n383) );
  NOR2_X1 U459 ( .A1(n658), .A2(n396), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n367), .B(n366), .ZN(n539) );
  INV_X1 U461 ( .A(KEYINPUT102), .ZN(n366) );
  NAND2_X1 U462 ( .A1(n379), .A2(n378), .ZN(n377) );
  NAND2_X1 U463 ( .A1(n376), .A2(n375), .ZN(n374) );
  XNOR2_X1 U464 ( .A(n435), .B(n369), .ZN(n439) );
  NOR2_X1 U465 ( .A1(n389), .A2(n668), .ZN(n533) );
  NAND2_X1 U466 ( .A1(n511), .A2(n397), .ZN(n640) );
  NOR2_X1 U467 ( .A1(n549), .A2(n547), .ZN(n509) );
  XNOR2_X1 U468 ( .A(n564), .B(n563), .ZN(n736) );
  XNOR2_X1 U469 ( .A(n575), .B(KEYINPUT32), .ZN(n739) );
  NOR2_X1 U470 ( .A1(n607), .A2(n707), .ZN(n609) );
  XNOR2_X1 U471 ( .A(n693), .B(n416), .ZN(n694) );
  NOR2_X1 U472 ( .A1(n615), .A2(n707), .ZN(n617) );
  XNOR2_X1 U473 ( .A(G101), .B(G110), .ZN(n352) );
  AND2_X1 U474 ( .A1(n385), .A2(n739), .ZN(n353) );
  XNOR2_X1 U475 ( .A(KEYINPUT100), .B(KEYINPUT7), .ZN(n354) );
  XNOR2_X1 U476 ( .A(n515), .B(n510), .ZN(n659) );
  XOR2_X1 U477 ( .A(n479), .B(KEYINPUT92), .Z(n355) );
  AND2_X1 U478 ( .A1(n601), .A2(n641), .ZN(n356) );
  AND2_X1 U479 ( .A1(n478), .A2(G221), .ZN(n357) );
  AND2_X1 U480 ( .A1(n641), .A2(n408), .ZN(n358) );
  XOR2_X1 U481 ( .A(n598), .B(KEYINPUT65), .Z(n359) );
  XNOR2_X1 U482 ( .A(n381), .B(n380), .ZN(n708) );
  NAND2_X1 U483 ( .A1(n601), .A2(n600), .ZN(n681) );
  XNOR2_X2 U484 ( .A(n553), .B(KEYINPUT81), .ZN(n601) );
  XNOR2_X1 U485 ( .A(n411), .B(KEYINPUT105), .ZN(n410) );
  INV_X1 U486 ( .A(n715), .ZN(n595) );
  NOR2_X1 U487 ( .A1(n696), .A2(n707), .ZN(n697) );
  XNOR2_X1 U488 ( .A(n361), .B(n357), .ZN(n703) );
  XNOR2_X1 U489 ( .A(n477), .B(n721), .ZN(n361) );
  XNOR2_X1 U490 ( .A(n514), .B(KEYINPUT28), .ZN(n516) );
  NOR2_X1 U491 ( .A1(n545), .A2(n362), .ZN(n390) );
  NAND2_X1 U492 ( .A1(n407), .A2(n595), .ZN(n365) );
  NAND2_X1 U493 ( .A1(n640), .A2(n512), .ZN(n522) );
  NAND2_X1 U494 ( .A1(n410), .A2(n409), .ZN(n547) );
  NAND2_X1 U495 ( .A1(n528), .A2(n453), .ZN(n367) );
  NAND2_X1 U496 ( .A1(n403), .A2(n402), .ZN(n401) );
  NOR2_X2 U497 ( .A1(n506), .A2(n580), .ZN(n536) );
  XNOR2_X2 U498 ( .A(n425), .B(n444), .ZN(n470) );
  INV_X1 U499 ( .A(n736), .ZN(n370) );
  NOR2_X1 U500 ( .A1(n559), .A2(n374), .ZN(n373) );
  INV_X1 U501 ( .A(n558), .ZN(n376) );
  NAND2_X1 U502 ( .A1(n559), .A2(KEYINPUT0), .ZN(n379) );
  NAND2_X1 U503 ( .A1(n395), .A2(n397), .ZN(n384) );
  INV_X1 U504 ( .A(n627), .ZN(n385) );
  XNOR2_X2 U505 ( .A(n386), .B(G472), .ZN(n662) );
  NAND2_X1 U506 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U507 ( .A1(n516), .A2(n515), .ZN(n389) );
  NOR2_X1 U508 ( .A1(n559), .A2(n388), .ZN(n387) );
  INV_X1 U509 ( .A(n515), .ZN(n388) );
  NAND2_X1 U510 ( .A1(n391), .A2(n390), .ZN(n546) );
  NAND2_X1 U511 ( .A1(n543), .A2(n392), .ZN(n391) );
  XNOR2_X2 U512 ( .A(n394), .B(n393), .ZN(n654) );
  NOR2_X1 U513 ( .A1(n659), .A2(n658), .ZN(n576) );
  XNOR2_X1 U514 ( .A(n401), .B(n400), .ZN(n552) );
  INV_X1 U515 ( .A(KEYINPUT48), .ZN(n400) );
  XNOR2_X1 U516 ( .A(n542), .B(n541), .ZN(n402) );
  NAND2_X1 U517 ( .A1(n546), .A2(KEYINPUT47), .ZN(n404) );
  AND2_X1 U518 ( .A1(n601), .A2(n358), .ZN(n407) );
  NAND2_X1 U519 ( .A1(n356), .A2(n595), .ZN(n682) );
  NAND2_X1 U520 ( .A1(n587), .A2(n513), .ZN(n411) );
  XNOR2_X1 U521 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U522 ( .A(KEYINPUT84), .B(KEYINPUT39), .ZN(n415) );
  XNOR2_X1 U523 ( .A(KEYINPUT59), .B(KEYINPUT117), .ZN(n416) );
  XNOR2_X1 U524 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n417) );
  XNOR2_X1 U525 ( .A(KEYINPUT46), .B(KEYINPUT83), .ZN(n541) );
  XNOR2_X1 U526 ( .A(n444), .B(n443), .ZN(n445) );
  INV_X1 U527 ( .A(n493), .ZN(n494) );
  XNOR2_X1 U528 ( .A(n460), .B(n448), .ZN(n449) );
  XNOR2_X1 U529 ( .A(n476), .B(n475), .ZN(n477) );
  INV_X1 U530 ( .A(KEYINPUT19), .ZN(n518) );
  INV_X1 U531 ( .A(KEYINPUT119), .ZN(n702) );
  XNOR2_X1 U532 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U533 ( .A(n562), .B(KEYINPUT80), .ZN(n563) );
  INV_X1 U534 ( .A(KEYINPUT63), .ZN(n608) );
  XNOR2_X1 U535 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U536 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n430) );
  NAND2_X1 U537 ( .A1(G214), .A2(n489), .ZN(n419) );
  XNOR2_X1 U538 ( .A(n420), .B(n419), .ZN(n424) );
  XNOR2_X1 U539 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U540 ( .A(n424), .B(n423), .Z(n428) );
  XOR2_X2 U541 ( .A(G146), .B(G125), .Z(n444) );
  XNOR2_X1 U542 ( .A(n426), .B(G122), .ZN(n442) );
  XNOR2_X1 U543 ( .A(n470), .B(n442), .ZN(n427) );
  XNOR2_X1 U544 ( .A(n428), .B(n427), .ZN(n693) );
  NOR2_X1 U545 ( .A1(G902), .A2(n693), .ZN(n429) );
  XNOR2_X1 U546 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U547 ( .A(KEYINPUT101), .B(KEYINPUT9), .Z(n433) );
  XNOR2_X1 U548 ( .A(n433), .B(n432), .ZN(n436) );
  XOR2_X1 U549 ( .A(G116), .B(G107), .Z(n441) );
  XNOR2_X1 U550 ( .A(n447), .B(n441), .ZN(n435) );
  NAND2_X1 U551 ( .A1(G234), .A2(n730), .ZN(n437) );
  XOR2_X1 U552 ( .A(KEYINPUT8), .B(n437), .Z(n478) );
  NAND2_X1 U553 ( .A1(G217), .A2(n478), .ZN(n438) );
  XNOR2_X1 U554 ( .A(n439), .B(n438), .ZN(n699) );
  NOR2_X1 U555 ( .A1(G902), .A2(n699), .ZN(n440) );
  XNOR2_X1 U556 ( .A(G478), .B(n440), .ZN(n528) );
  NOR2_X1 U557 ( .A1(n453), .A2(n528), .ZN(n623) );
  NOR2_X1 U558 ( .A1(n623), .A2(n539), .ZN(n649) );
  NAND2_X1 U559 ( .A1(n649), .A2(KEYINPUT47), .ZN(n502) );
  INV_X1 U560 ( .A(KEYINPUT72), .ZN(n446) );
  NAND2_X1 U561 ( .A1(G224), .A2(n730), .ZN(n448) );
  XNOR2_X1 U562 ( .A(n450), .B(KEYINPUT69), .ZN(n486) );
  AND2_X1 U563 ( .A1(G210), .A2(n486), .ZN(n451) );
  INV_X1 U564 ( .A(n549), .ZN(n517) );
  NOR2_X1 U565 ( .A1(n529), .A2(n528), .ZN(n560) );
  XOR2_X1 U566 ( .A(n455), .B(n454), .Z(n456) );
  NAND2_X1 U567 ( .A1(G952), .A2(n456), .ZN(n674) );
  NOR2_X1 U568 ( .A1(G953), .A2(n674), .ZN(n556) );
  AND2_X1 U569 ( .A1(n456), .A2(G953), .ZN(n457) );
  NAND2_X1 U570 ( .A1(G902), .A2(n457), .ZN(n555) );
  XNOR2_X1 U571 ( .A(n555), .B(KEYINPUT104), .ZN(n458) );
  NOR2_X1 U572 ( .A1(G900), .A2(n458), .ZN(n459) );
  NOR2_X1 U573 ( .A1(n556), .A2(n459), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n469), .B(n462), .ZN(n463) );
  XOR2_X1 U575 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n465) );
  NAND2_X1 U576 ( .A1(G227), .A2(n730), .ZN(n464) );
  NOR2_X1 U577 ( .A1(n687), .A2(G902), .ZN(n468) );
  INV_X1 U578 ( .A(G469), .ZN(n467) );
  XOR2_X1 U579 ( .A(G110), .B(KEYINPUT90), .Z(n472) );
  XNOR2_X1 U580 ( .A(G119), .B(KEYINPUT68), .ZN(n471) );
  XNOR2_X1 U581 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U582 ( .A(KEYINPUT25), .B(KEYINPUT71), .ZN(n479) );
  NAND2_X1 U583 ( .A1(G234), .A2(n596), .ZN(n480) );
  XNOR2_X1 U584 ( .A(KEYINPUT20), .B(n480), .ZN(n482) );
  AND2_X1 U585 ( .A1(n482), .A2(G217), .ZN(n481) );
  NAND2_X1 U586 ( .A1(n482), .A2(G221), .ZN(n483) );
  XNOR2_X1 U587 ( .A(n483), .B(KEYINPUT21), .ZN(n484) );
  XNOR2_X1 U588 ( .A(KEYINPUT93), .B(n484), .ZN(n655) );
  AND2_X1 U589 ( .A1(n654), .A2(n655), .ZN(n485) );
  NAND2_X1 U590 ( .A1(n515), .A2(n485), .ZN(n580) );
  NAND2_X1 U591 ( .A1(G214), .A2(n486), .ZN(n646) );
  XNOR2_X1 U592 ( .A(n488), .B(n487), .ZN(n496) );
  XOR2_X1 U593 ( .A(KEYINPUT70), .B(KEYINPUT94), .Z(n491) );
  NAND2_X1 U594 ( .A1(n489), .A2(G210), .ZN(n490) );
  XNOR2_X1 U595 ( .A(n491), .B(n490), .ZN(n492) );
  NAND2_X1 U596 ( .A1(n646), .A2(n662), .ZN(n499) );
  XNOR2_X1 U597 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n497) );
  XNOR2_X1 U598 ( .A(n497), .B(KEYINPUT30), .ZN(n498) );
  XNOR2_X1 U599 ( .A(n499), .B(n498), .ZN(n535) );
  AND2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n500) );
  AND2_X1 U601 ( .A1(n560), .A2(n500), .ZN(n501) );
  NAND2_X1 U602 ( .A1(n517), .A2(n501), .ZN(n631) );
  NAND2_X1 U603 ( .A1(n502), .A2(n631), .ZN(n503) );
  NAND2_X1 U604 ( .A1(n503), .A2(KEYINPUT77), .ZN(n505) );
  INV_X1 U605 ( .A(KEYINPUT77), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n544), .A2(n631), .ZN(n504) );
  NAND2_X1 U607 ( .A1(n505), .A2(n504), .ZN(n512) );
  INV_X1 U608 ( .A(n539), .ZN(n634) );
  INV_X1 U609 ( .A(n655), .ZN(n565) );
  NOR2_X1 U610 ( .A1(n565), .A2(n506), .ZN(n507) );
  XNOR2_X1 U611 ( .A(n507), .B(KEYINPUT67), .ZN(n508) );
  NOR2_X1 U612 ( .A1(n654), .A2(n508), .ZN(n513) );
  XNOR2_X1 U613 ( .A(n509), .B(KEYINPUT36), .ZN(n511) );
  INV_X1 U614 ( .A(KEYINPUT1), .ZN(n510) );
  AND2_X1 U615 ( .A1(n662), .A2(n513), .ZN(n514) );
  XNOR2_X2 U616 ( .A(n520), .B(KEYINPUT75), .ZN(n632) );
  NOR2_X1 U617 ( .A1(KEYINPUT78), .A2(n632), .ZN(n521) );
  NOR2_X1 U618 ( .A1(n522), .A2(n521), .ZN(n527) );
  NOR2_X1 U619 ( .A1(n649), .A2(n632), .ZN(n543) );
  NAND2_X1 U620 ( .A1(KEYINPUT66), .A2(n543), .ZN(n523) );
  NAND2_X1 U621 ( .A1(n523), .A2(KEYINPUT78), .ZN(n525) );
  INV_X1 U622 ( .A(KEYINPUT47), .ZN(n524) );
  NAND2_X1 U623 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U624 ( .A(KEYINPUT38), .B(n549), .ZN(n647) );
  NAND2_X1 U625 ( .A1(n529), .A2(n528), .ZN(n644) );
  INV_X1 U626 ( .A(n646), .ZN(n530) );
  NOR2_X1 U627 ( .A1(n644), .A2(n530), .ZN(n531) );
  AND2_X1 U628 ( .A1(n647), .A2(n531), .ZN(n532) );
  XNOR2_X1 U629 ( .A(n533), .B(KEYINPUT42), .ZN(n534) );
  XNOR2_X1 U630 ( .A(n534), .B(KEYINPUT109), .ZN(n734) );
  AND2_X1 U631 ( .A1(n647), .A2(n535), .ZN(n537) );
  NAND2_X1 U632 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X2 U633 ( .A(n538), .B(n415), .ZN(n554) );
  XOR2_X1 U634 ( .A(KEYINPUT40), .B(n540), .Z(n735) );
  NAND2_X1 U635 ( .A1(n734), .A2(n735), .ZN(n542) );
  AND2_X1 U636 ( .A1(n544), .A2(n649), .ZN(n545) );
  OR2_X1 U637 ( .A1(n397), .A2(n547), .ZN(n548) );
  XNOR2_X1 U638 ( .A(n548), .B(KEYINPUT43), .ZN(n550) );
  NAND2_X1 U639 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U640 ( .A(KEYINPUT106), .B(n551), .ZN(n738) );
  NAND2_X1 U641 ( .A1(n552), .A2(n738), .ZN(n553) );
  NAND2_X1 U642 ( .A1(n623), .A2(n554), .ZN(n641) );
  NOR2_X1 U643 ( .A1(G898), .A2(n555), .ZN(n557) );
  NOR2_X1 U644 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U645 ( .A1(n654), .A2(n655), .ZN(n658) );
  NAND2_X1 U646 ( .A1(n561), .A2(n560), .ZN(n564) );
  XOR2_X1 U647 ( .A(KEYINPUT73), .B(KEYINPUT35), .Z(n562) );
  OR2_X1 U648 ( .A1(n644), .A2(n565), .ZN(n566) );
  INV_X1 U649 ( .A(KEYINPUT22), .ZN(n567) );
  XNOR2_X1 U650 ( .A(n568), .B(n567), .ZN(n572) );
  OR2_X1 U651 ( .A1(n654), .A2(n662), .ZN(n569) );
  XOR2_X1 U652 ( .A(n587), .B(KEYINPUT74), .Z(n574) );
  NOR2_X1 U653 ( .A1(n654), .A2(n659), .ZN(n570) );
  XNOR2_X1 U654 ( .A(KEYINPUT103), .B(n570), .ZN(n571) );
  NOR2_X1 U655 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U656 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U657 ( .A1(n662), .A2(n576), .ZN(n577) );
  XOR2_X1 U658 ( .A(KEYINPUT95), .B(n577), .Z(n665) );
  NOR2_X1 U659 ( .A1(n581), .A2(n665), .ZN(n579) );
  XNOR2_X1 U660 ( .A(KEYINPUT96), .B(KEYINPUT31), .ZN(n578) );
  XNOR2_X1 U661 ( .A(n579), .B(n578), .ZN(n637) );
  INV_X1 U662 ( .A(n580), .ZN(n583) );
  NOR2_X1 U663 ( .A1(n662), .A2(n581), .ZN(n582) );
  NAND2_X1 U664 ( .A1(n583), .A2(n582), .ZN(n624) );
  NAND2_X1 U665 ( .A1(n637), .A2(n624), .ZN(n584) );
  XNOR2_X1 U666 ( .A(KEYINPUT97), .B(n584), .ZN(n585) );
  NOR2_X1 U667 ( .A1(n585), .A2(n649), .ZN(n590) );
  NOR2_X1 U668 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U669 ( .A1(n654), .A2(n588), .ZN(n618) );
  XOR2_X1 U670 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n593) );
  XNOR2_X2 U671 ( .A(n594), .B(n593), .ZN(n715) );
  XNOR2_X1 U672 ( .A(KEYINPUT79), .B(n596), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n597), .A2(KEYINPUT2), .ZN(n598) );
  NAND2_X1 U674 ( .A1(KEYINPUT2), .A2(n641), .ZN(n599) );
  XOR2_X1 U675 ( .A(KEYINPUT76), .B(n599), .Z(n600) );
  NAND2_X1 U676 ( .A1(n418), .A2(G472), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n604), .B(n417), .ZN(n605) );
  XNOR2_X1 U678 ( .A(n606), .B(n605), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n609), .B(n608), .ZN(G57) );
  XOR2_X1 U680 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n612) );
  XNOR2_X1 U681 ( .A(n610), .B(KEYINPUT85), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n612), .B(n611), .ZN(n614) );
  NAND2_X1 U683 ( .A1(n418), .A2(G210), .ZN(n613) );
  XNOR2_X1 U684 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U685 ( .A(KEYINPUT82), .B(KEYINPUT56), .ZN(n616) );
  XNOR2_X1 U686 ( .A(n617), .B(n616), .ZN(G51) );
  XNOR2_X1 U687 ( .A(G101), .B(n618), .ZN(G3) );
  NOR2_X1 U688 ( .A1(n634), .A2(n624), .ZN(n620) );
  XNOR2_X1 U689 ( .A(G104), .B(KEYINPUT111), .ZN(n619) );
  XNOR2_X1 U690 ( .A(n620), .B(n619), .ZN(G6) );
  XOR2_X1 U691 ( .A(KEYINPUT112), .B(KEYINPUT26), .Z(n622) );
  XNOR2_X1 U692 ( .A(G107), .B(KEYINPUT27), .ZN(n621) );
  XNOR2_X1 U693 ( .A(n622), .B(n621), .ZN(n626) );
  INV_X1 U694 ( .A(n623), .ZN(n636) );
  NOR2_X1 U695 ( .A1(n636), .A2(n624), .ZN(n625) );
  XOR2_X1 U696 ( .A(n626), .B(n625), .Z(G9) );
  XOR2_X1 U697 ( .A(G110), .B(n627), .Z(G12) );
  NOR2_X1 U698 ( .A1(n636), .A2(n632), .ZN(n629) );
  XNOR2_X1 U699 ( .A(KEYINPUT113), .B(KEYINPUT29), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n629), .B(n628), .ZN(n630) );
  XOR2_X1 U701 ( .A(G128), .B(n630), .Z(G30) );
  XNOR2_X1 U702 ( .A(G143), .B(n631), .ZN(G45) );
  NOR2_X1 U703 ( .A1(n634), .A2(n632), .ZN(n633) );
  XOR2_X1 U704 ( .A(G146), .B(n633), .Z(G48) );
  NOR2_X1 U705 ( .A1(n634), .A2(n637), .ZN(n635) );
  XOR2_X1 U706 ( .A(G113), .B(n635), .Z(G15) );
  NOR2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U708 ( .A(G116), .B(n638), .Z(G18) );
  XOR2_X1 U709 ( .A(G125), .B(KEYINPUT37), .Z(n639) );
  XNOR2_X1 U710 ( .A(n640), .B(n639), .ZN(G27) );
  XNOR2_X1 U711 ( .A(G134), .B(n641), .ZN(G36) );
  NOR2_X1 U712 ( .A1(n653), .A2(n668), .ZN(n642) );
  NOR2_X1 U713 ( .A1(G953), .A2(n642), .ZN(n680) );
  NOR2_X1 U714 ( .A1(n647), .A2(n646), .ZN(n643) );
  NOR2_X1 U715 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U716 ( .A(KEYINPUT115), .B(n645), .Z(n651) );
  NAND2_X1 U717 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U719 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U720 ( .A1(n653), .A2(n652), .ZN(n671) );
  NOR2_X1 U721 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U722 ( .A(n656), .B(KEYINPUT49), .ZN(n657) );
  XNOR2_X1 U723 ( .A(n657), .B(KEYINPUT114), .ZN(n664) );
  NAND2_X1 U724 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U725 ( .A(KEYINPUT50), .B(n660), .Z(n661) );
  NOR2_X1 U726 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U727 ( .A1(n664), .A2(n663), .ZN(n666) );
  NAND2_X1 U728 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U729 ( .A(KEYINPUT51), .B(n667), .ZN(n669) );
  NOR2_X1 U730 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U731 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U732 ( .A(n672), .B(KEYINPUT52), .ZN(n673) );
  NOR2_X1 U733 ( .A1(n674), .A2(n673), .ZN(n678) );
  INV_X1 U734 ( .A(KEYINPUT2), .ZN(n675) );
  NOR2_X1 U735 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U736 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U737 ( .A1(n680), .A2(n679), .ZN(n685) );
  INV_X1 U738 ( .A(n681), .ZN(n683) );
  NOR2_X1 U739 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U740 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U741 ( .A(KEYINPUT53), .B(n686), .ZN(G75) );
  XNOR2_X1 U742 ( .A(KEYINPUT58), .B(KEYINPUT116), .ZN(n689) );
  XNOR2_X1 U743 ( .A(n687), .B(KEYINPUT57), .ZN(n688) );
  XNOR2_X1 U744 ( .A(n689), .B(n688), .ZN(n691) );
  NAND2_X1 U745 ( .A1(n418), .A2(G469), .ZN(n690) );
  XOR2_X1 U746 ( .A(n691), .B(n690), .Z(n692) );
  NOR2_X1 U747 ( .A1(n707), .A2(n692), .ZN(G54) );
  NAND2_X1 U748 ( .A1(n418), .A2(G475), .ZN(n695) );
  XNOR2_X1 U749 ( .A(KEYINPUT60), .B(n697), .ZN(G60) );
  NAND2_X1 U750 ( .A1(n418), .A2(G478), .ZN(n698) );
  XNOR2_X1 U751 ( .A(n698), .B(KEYINPUT118), .ZN(n700) );
  XNOR2_X1 U752 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U753 ( .A1(n707), .A2(n701), .ZN(G63) );
  NAND2_X1 U754 ( .A1(n418), .A2(G217), .ZN(n705) );
  NOR2_X1 U755 ( .A1(n707), .A2(n706), .ZN(G66) );
  XNOR2_X1 U756 ( .A(KEYINPUT123), .B(n708), .ZN(n710) );
  NOR2_X1 U757 ( .A1(n730), .A2(G898), .ZN(n709) );
  NOR2_X1 U758 ( .A1(n710), .A2(n709), .ZN(n720) );
  NAND2_X1 U759 ( .A1(G224), .A2(G953), .ZN(n711) );
  XNOR2_X1 U760 ( .A(n711), .B(KEYINPUT120), .ZN(n712) );
  XNOR2_X1 U761 ( .A(KEYINPUT61), .B(n712), .ZN(n713) );
  NAND2_X1 U762 ( .A1(n713), .A2(G898), .ZN(n714) );
  XNOR2_X1 U763 ( .A(n714), .B(KEYINPUT121), .ZN(n717) );
  NOR2_X1 U764 ( .A1(G953), .A2(n715), .ZN(n716) );
  NOR2_X1 U765 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U766 ( .A(n718), .B(KEYINPUT122), .Z(n719) );
  XNOR2_X1 U767 ( .A(n720), .B(n719), .ZN(G69) );
  XNOR2_X1 U768 ( .A(KEYINPUT87), .B(KEYINPUT124), .ZN(n724) );
  XNOR2_X1 U769 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U770 ( .A(n724), .B(n723), .ZN(n729) );
  XNOR2_X1 U771 ( .A(n729), .B(G227), .ZN(n725) );
  XNOR2_X1 U772 ( .A(n725), .B(KEYINPUT125), .ZN(n726) );
  NAND2_X1 U773 ( .A1(n726), .A2(G900), .ZN(n727) );
  XNOR2_X1 U774 ( .A(KEYINPUT126), .B(n727), .ZN(n728) );
  NAND2_X1 U775 ( .A1(n728), .A2(G953), .ZN(n733) );
  XNOR2_X1 U776 ( .A(n356), .B(n729), .ZN(n731) );
  NAND2_X1 U777 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U778 ( .A1(n733), .A2(n732), .ZN(G72) );
  XNOR2_X1 U779 ( .A(n734), .B(G137), .ZN(G39) );
  XNOR2_X1 U780 ( .A(G131), .B(n735), .ZN(G33) );
  XNOR2_X1 U781 ( .A(G122), .B(KEYINPUT127), .ZN(n737) );
  XNOR2_X1 U782 ( .A(n737), .B(n736), .ZN(G24) );
  XNOR2_X1 U783 ( .A(G140), .B(n738), .ZN(G42) );
  XNOR2_X1 U784 ( .A(n739), .B(G119), .ZN(G21) );
endmodule

