//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1259, new_n1260, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n209), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n209), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n206), .A2(G50), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g0024(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G20), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n221), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n217), .A2(new_n220), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n216), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n202), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n242), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G232), .A3(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G97), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  OAI211_X1 g0059(.A(G226), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n255), .A2(new_n256), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n226), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  AND2_X1   g0066(.A1(G1), .A2(G13), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(new_n262), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G238), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n262), .A2(G1), .A3(G13), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n270), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n272), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n265), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n278), .B1(new_n265), .B2(new_n277), .ZN(new_n281));
  OAI21_X1  g0081(.A(G200), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n265), .A2(new_n277), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT13), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(G190), .A3(new_n279), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n224), .A2(new_n225), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT69), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n224), .A2(KEYINPUT69), .A3(new_n225), .A4(new_n286), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n292), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n293));
  INV_X1    g0093(.A(G77), .ZN(new_n294));
  INV_X1    g0094(.A(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G33), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n293), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n291), .A2(KEYINPUT11), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G13), .ZN(new_n299));
  NOR3_X1   g0099(.A1(new_n299), .A2(new_n295), .A3(G1), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(new_n289), .B2(new_n290), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n269), .A2(G20), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(G68), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n297), .A2(new_n289), .A3(new_n290), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT11), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n300), .A2(new_n202), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT12), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n298), .A2(new_n303), .A3(new_n306), .A4(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n282), .A2(new_n285), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT13), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n276), .B1(new_n264), .B2(new_n261), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n279), .B(G179), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT74), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n284), .A2(KEYINPUT74), .A3(G179), .A4(new_n279), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(G169), .B1(new_n280), .B2(new_n281), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT14), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT14), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n322), .B(G169), .C1(new_n280), .C2(new_n281), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n319), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n312), .B1(new_n324), .B2(new_n309), .ZN(new_n325));
  OR2_X1    g0125(.A1(KEYINPUT8), .A2(G58), .ZN(new_n326));
  NAND2_X1  g0126(.A1(KEYINPUT8), .A2(G58), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n302), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT77), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n301), .ZN(new_n332));
  INV_X1    g0132(.A(new_n300), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n331), .A2(new_n332), .B1(new_n333), .B2(new_n328), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT16), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G58), .A2(G68), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n203), .A2(new_n205), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G20), .ZN(new_n338));
  INV_X1    g0138(.A(G159), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n339), .A2(G20), .A3(G33), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT75), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT75), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n338), .A2(new_n344), .A3(new_n341), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT76), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n258), .A2(new_n259), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT7), .B1(new_n348), .B2(new_n295), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n295), .A4(new_n253), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n347), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n252), .A2(new_n295), .A3(new_n253), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n347), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n202), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n335), .B1(new_n346), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n289), .A2(new_n290), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n344), .B1(new_n338), .B2(new_n341), .ZN(new_n360));
  AOI211_X1 g0160(.A(KEYINPUT75), .B(new_n340), .C1(new_n337), .C2(G20), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n353), .A2(new_n354), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n202), .B1(new_n363), .B2(new_n350), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n335), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n359), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n334), .B1(new_n358), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n272), .B1(new_n232), .B2(new_n275), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n254), .A2(G223), .A3(new_n257), .ZN(new_n369));
  OAI211_X1 g0169(.A(G226), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G87), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n368), .B1(new_n264), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G179), .ZN(new_n374));
  INV_X1    g0174(.A(G169), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(new_n373), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT18), .B1(new_n367), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n329), .B(KEYINPUT77), .ZN(new_n379));
  INV_X1    g0179(.A(new_n328), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n379), .A2(new_n301), .B1(new_n300), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(G68), .B1(new_n349), .B2(new_n351), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT16), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n291), .B1(new_n346), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT76), .B1(new_n363), .B2(new_n350), .ZN(new_n385));
  OAI21_X1  g0185(.A(G68), .B1(new_n385), .B2(new_n355), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT16), .B1(new_n362), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n381), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT18), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(new_n376), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n378), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n372), .A2(new_n264), .ZN(new_n393));
  INV_X1    g0193(.A(new_n368), .ZN(new_n394));
  INV_X1    g0194(.A(G190), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(G200), .B2(new_n373), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n381), .B(new_n397), .C1(new_n384), .C2(new_n387), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT17), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n358), .A2(new_n366), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n401), .A2(KEYINPUT17), .A3(new_n381), .A4(new_n397), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n325), .A2(new_n392), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n406));
  INV_X1    g0206(.A(G150), .ZN(new_n407));
  INV_X1    g0207(.A(new_n292), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n406), .B1(new_n407), .B2(new_n408), .C1(new_n380), .C2(new_n296), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n409), .A2(new_n291), .B1(new_n243), .B2(new_n300), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n301), .A2(G50), .A3(new_n302), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n410), .A2(KEYINPUT9), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT9), .B1(new_n410), .B2(new_n411), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G223), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT67), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(new_n348), .B2(new_n257), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n254), .A2(KEYINPUT67), .A3(G1698), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(G1698), .B1(new_n252), .B2(new_n253), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G222), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n294), .B2(new_n254), .ZN(new_n422));
  OR3_X1    g0222(.A1(new_n419), .A2(new_n422), .A3(KEYINPUT68), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT68), .B1(new_n419), .B2(new_n422), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n264), .ZN(new_n425));
  INV_X1    g0225(.A(new_n272), .ZN(new_n426));
  INV_X1    g0226(.A(new_n275), .ZN(new_n427));
  XOR2_X1   g0227(.A(KEYINPUT66), .B(G226), .Z(new_n428));
  AOI21_X1  g0228(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n425), .A2(G190), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n425), .A2(new_n429), .ZN(new_n431));
  XOR2_X1   g0231(.A(KEYINPUT71), .B(G200), .Z(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n414), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT10), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT10), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n414), .A2(new_n437), .A3(new_n434), .A4(new_n430), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n431), .A2(G179), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT70), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n410), .A2(new_n411), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n431), .B2(new_n375), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  OAI22_X1  g0244(.A1(new_n380), .A2(new_n408), .B1(new_n295), .B2(new_n294), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT15), .B(G87), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(new_n296), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n291), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n301), .A2(G77), .A3(new_n302), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n300), .A2(new_n294), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n273), .B1(new_n417), .B2(new_n418), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n254), .A2(G232), .A3(new_n257), .ZN(new_n453));
  INV_X1    g0253(.A(G107), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(new_n254), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n264), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n426), .B1(G244), .B2(new_n427), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n451), .B1(new_n375), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n458), .ZN(new_n460));
  INV_X1    g0260(.A(G179), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n451), .B1(new_n458), .B2(new_n395), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(new_n433), .B2(new_n458), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n439), .A2(new_n444), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT72), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT72), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n439), .A2(new_n444), .A3(new_n470), .A4(new_n467), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n405), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n295), .B(G87), .C1(new_n258), .C2(new_n259), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT22), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT22), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n254), .A2(new_n475), .A3(new_n295), .A4(G87), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT86), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n251), .A2(new_n479), .A3(G20), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT23), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n295), .B2(G107), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n454), .A2(KEYINPUT23), .A3(G20), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n477), .A2(new_n478), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n478), .B1(new_n477), .B2(new_n484), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT24), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT24), .ZN(new_n488));
  AOI21_X1  g0288(.A(G20), .B1(new_n252), .B2(new_n253), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n475), .B1(new_n489), .B2(G87), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n473), .A2(KEYINPUT22), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n484), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT86), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n477), .A2(new_n478), .A3(new_n484), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n488), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n291), .B1(new_n487), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n251), .A2(G1), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n301), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(new_n454), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n300), .A2(new_n454), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n501), .B(KEYINPUT25), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n496), .A2(KEYINPUT87), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT87), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT24), .B1(new_n485), .B2(new_n486), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n493), .A2(new_n488), .A3(new_n494), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n359), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n503), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT79), .ZN(new_n511));
  INV_X1    g0311(.A(G41), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT5), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT5), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(KEYINPUT79), .B2(G41), .ZN(new_n515));
  INV_X1    g0315(.A(G45), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(G1), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n268), .A2(new_n513), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n513), .A2(new_n515), .A3(new_n517), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n519), .A2(new_n274), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G264), .ZN(new_n521));
  OAI211_X1 g0321(.A(G257), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n522));
  INV_X1    g0322(.A(G294), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n522), .B1(new_n251), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT88), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n420), .A2(new_n525), .A3(G250), .ZN(new_n526));
  OAI211_X1 g0326(.A(G250), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT88), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n524), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n518), .B(new_n521), .C1(new_n529), .C2(new_n263), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G169), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n526), .A2(new_n528), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n264), .B1(new_n532), .B2(new_n524), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n533), .A2(G179), .A3(new_n518), .A4(new_n521), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n504), .A2(new_n510), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(G200), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n533), .A2(new_n395), .A3(new_n518), .A4(new_n521), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n496), .A2(new_n503), .A3(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G238), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n542));
  OAI211_X1 g0342(.A(G244), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n543), .C1(new_n251), .C2(new_n479), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n264), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n274), .A2(G274), .A3(new_n517), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n269), .A2(G45), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n274), .A2(G250), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n545), .A2(new_n461), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n549), .B1(new_n544), .B2(new_n264), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(G169), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n446), .ZN(new_n554));
  AND4_X1   g0354(.A1(new_n359), .A2(new_n333), .A3(new_n554), .A4(new_n498), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n295), .B1(new_n256), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(G97), .A2(G107), .ZN(new_n558));
  INV_X1    g0358(.A(G87), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n295), .B(G68), .C1(new_n258), .C2(new_n259), .ZN(new_n562));
  INV_X1    g0362(.A(G97), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n556), .B1(new_n296), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(new_n289), .A3(new_n290), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n554), .A2(new_n333), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(KEYINPUT81), .B1(new_n555), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n567), .B1(new_n291), .B2(new_n565), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT81), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n301), .A2(new_n554), .A3(new_n498), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n553), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n552), .A2(G190), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n359), .A2(G87), .A3(new_n333), .A4(new_n498), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n578), .A2(new_n566), .A3(new_n568), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n552), .A2(new_n432), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n577), .B1(new_n581), .B2(KEYINPUT82), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT82), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n579), .B2(new_n580), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n575), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(G244), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT4), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(KEYINPUT78), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G283), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(KEYINPUT78), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n254), .A2(G244), .A3(new_n257), .A4(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n254), .A2(G250), .A3(G1698), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n588), .A2(new_n589), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n264), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n519), .A2(G257), .A3(new_n274), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n518), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT80), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n594), .A2(KEYINPUT80), .A3(new_n597), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(G190), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(G107), .B1(new_n385), .B2(new_n355), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT6), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n563), .A2(new_n454), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n604), .B1(new_n605), .B2(new_n558), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n454), .A2(KEYINPUT6), .A3(G97), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n608), .A2(G20), .B1(G77), .B2(new_n292), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n359), .B1(new_n603), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n499), .A2(new_n563), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n333), .A2(G97), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n598), .A2(G200), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n602), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI211_X1 g0415(.A(G179), .B(new_n596), .C1(new_n593), .C2(new_n264), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n454), .B1(new_n352), .B2(new_n356), .ZN(new_n617));
  INV_X1    g0417(.A(new_n609), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n291), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI211_X1 g0419(.A(new_n300), .B(new_n497), .C1(new_n289), .C2(new_n290), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n612), .B1(new_n620), .B2(G97), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n616), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  AOI211_X1 g0422(.A(new_n599), .B(new_n596), .C1(new_n593), .C2(new_n264), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT80), .B1(new_n594), .B2(new_n597), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n375), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n585), .A2(new_n615), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(G20), .B1(G33), .B2(G283), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n251), .A2(G97), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n628), .A2(new_n629), .B1(G20), .B2(new_n479), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n630), .A2(new_n287), .A3(KEYINPUT20), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT20), .B1(new_n630), .B2(new_n287), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n631), .A2(new_n632), .B1(G116), .B2(new_n333), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n301), .A2(G116), .A3(new_n498), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT85), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT85), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n620), .A2(new_n636), .A3(G116), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n633), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(G257), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n639));
  OAI211_X1 g0439(.A(G264), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n640));
  XNOR2_X1  g0440(.A(KEYINPUT83), .B(G303), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n639), .B(new_n640), .C1(new_n254), .C2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT84), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n641), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n348), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n646), .A2(KEYINPUT84), .A3(new_n639), .A4(new_n640), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n644), .A2(new_n647), .A3(new_n264), .ZN(new_n648));
  INV_X1    g0448(.A(new_n518), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n520), .B2(G270), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G200), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n638), .B(new_n652), .C1(new_n395), .C2(new_n651), .ZN(new_n653));
  INV_X1    g0453(.A(new_n633), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n634), .A2(KEYINPUT85), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n636), .B1(new_n620), .B2(G116), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n375), .B1(new_n648), .B2(new_n650), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(KEYINPUT21), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT21), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n651), .A2(G169), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n638), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n651), .A2(new_n461), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n653), .A2(new_n659), .A3(new_n662), .A4(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n627), .A2(new_n665), .ZN(new_n666));
  AND4_X1   g0466(.A1(new_n472), .A2(new_n536), .A3(new_n541), .A4(new_n666), .ZN(G372));
  NAND3_X1  g0467(.A1(new_n659), .A2(new_n662), .A3(new_n664), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n496), .A2(new_n503), .B1(new_n531), .B2(new_n534), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n575), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n541), .A2(new_n672), .A3(new_n615), .A4(new_n626), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT89), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n541), .A2(new_n615), .A3(new_n626), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT89), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n535), .B1(new_n508), .B2(new_n509), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n677), .A2(new_n662), .A3(new_n664), .A4(new_n659), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n675), .A2(new_n676), .A3(new_n678), .A4(new_n672), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n622), .A2(new_n625), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n680), .B1(new_n585), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n552), .A2(G169), .ZN(new_n683));
  AOI211_X1 g0483(.A(G179), .B(new_n549), .C1(new_n264), .C2(new_n544), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n555), .A2(new_n569), .A3(KEYINPUT81), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n572), .B1(new_n571), .B2(new_n573), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n581), .A2(new_n576), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n688), .A2(new_n622), .A3(new_n625), .A4(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(new_n690), .B2(KEYINPUT26), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n682), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n674), .A2(new_n679), .A3(new_n692), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n472), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n324), .A2(new_n309), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n463), .B2(new_n312), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n391), .B1(new_n696), .B2(new_n404), .ZN(new_n697));
  INV_X1    g0497(.A(new_n439), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n444), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n694), .A2(new_n699), .ZN(G369));
  NAND3_X1  g0500(.A1(new_n269), .A2(new_n295), .A3(G13), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G213), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G343), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n638), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n665), .B2(KEYINPUT90), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(KEYINPUT90), .B2(new_n665), .ZN(new_n710));
  INV_X1    g0510(.A(new_n668), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n708), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G330), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n536), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n706), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n504), .A2(new_n510), .A3(new_n706), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n536), .A2(new_n718), .A3(new_n541), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n669), .A2(new_n707), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n711), .A2(new_n706), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(new_n536), .A3(new_n541), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(G399));
  INV_X1    g0525(.A(new_n218), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G41), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n560), .A2(G116), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(G1), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n221), .B2(new_n728), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT28), .Z(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n693), .A2(new_n733), .A3(new_n707), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT26), .B1(new_n585), .B2(new_n681), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT92), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n681), .A2(KEYINPUT26), .A3(new_n672), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(KEYINPUT92), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n673), .B1(new_n536), .B2(new_n711), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n575), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n706), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n734), .B1(new_n742), .B2(new_n733), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n666), .A2(new_n536), .A3(new_n541), .A4(new_n707), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n623), .A2(new_n624), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT91), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(new_n651), .B2(new_n461), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n648), .A2(KEYINPUT91), .A3(new_n650), .A4(G179), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n533), .A2(new_n521), .A3(new_n552), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n745), .A2(new_n747), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT30), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n749), .A2(new_n623), .A3(new_n624), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n754), .A2(KEYINPUT30), .A3(new_n748), .A4(new_n747), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n552), .A2(G179), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n651), .A2(new_n530), .A3(new_n598), .A4(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n753), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n706), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT31), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n744), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G330), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n743), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n732), .B1(new_n767), .B2(new_n269), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT93), .ZN(G364));
  OR2_X1    g0569(.A1(new_n715), .A2(KEYINPUT94), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n715), .A2(KEYINPUT94), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n299), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n269), .B1(new_n773), .B2(G45), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n727), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n713), .B2(new_n714), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G13), .A2(G33), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n713), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n226), .B1(new_n295), .B2(G169), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(G20), .A2(G179), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT96), .ZN(new_n785));
  AOI21_X1  g0585(.A(G200), .B1(new_n784), .B2(KEYINPUT96), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n395), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n784), .A2(new_n395), .A3(new_n537), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n789), .A2(new_n201), .B1(new_n243), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT97), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n787), .B2(G190), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n785), .A2(new_n786), .A3(KEYINPUT97), .A4(new_n395), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n792), .B1(new_n796), .B2(G77), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT98), .Z(new_n798));
  NOR2_X1   g0598(.A1(new_n295), .A2(G190), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G179), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n801), .A2(KEYINPUT32), .A3(new_n339), .ZN(new_n802));
  OAI21_X1  g0602(.A(KEYINPUT32), .B1(new_n801), .B2(new_n339), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n295), .B1(new_n800), .B2(G190), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n563), .B2(new_n804), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n784), .A2(new_n537), .A3(G190), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n348), .B1(new_n806), .B2(G68), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n295), .A2(new_n395), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n433), .A2(new_n461), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n433), .A2(new_n461), .A3(new_n799), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n807), .B1(new_n809), .B2(new_n559), .C1(new_n454), .C2(new_n810), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n798), .A2(new_n802), .A3(new_n805), .A4(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G326), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n791), .A2(new_n813), .B1(new_n804), .B2(new_n523), .ZN(new_n814));
  AOI22_X1  g0614(.A1(KEYINPUT99), .A2(new_n814), .B1(new_n788), .B2(G322), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(KEYINPUT99), .B2(new_n814), .ZN(new_n816));
  INV_X1    g0616(.A(G317), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT33), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n817), .A2(KEYINPUT33), .ZN(new_n819));
  AND3_X1   g0619(.A1(new_n806), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n801), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n254), .B(new_n820), .C1(G329), .C2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  INV_X1    g0623(.A(G303), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n822), .B1(new_n823), .B2(new_n810), .C1(new_n824), .C2(new_n809), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n816), .B(new_n825), .C1(G311), .C2(new_n796), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n783), .B1(new_n812), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n776), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n254), .A2(new_n218), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT95), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n830), .A2(G355), .B1(new_n479), .B2(new_n726), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n248), .A2(new_n516), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n726), .A2(new_n254), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n221), .B2(G45), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n831), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n783), .A2(new_n780), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n828), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n827), .A2(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n772), .A2(new_n777), .B1(new_n781), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G396));
  NAND2_X1  g0640(.A1(new_n782), .A2(new_n779), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n776), .B1(new_n841), .B2(G77), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n559), .A2(new_n810), .B1(new_n809), .B2(new_n454), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n804), .A2(new_n563), .ZN(new_n844));
  INV_X1    g0644(.A(G311), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n348), .B1(new_n801), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n806), .ZN(new_n847));
  XOR2_X1   g0647(.A(KEYINPUT100), .B(G283), .Z(new_n848));
  OAI22_X1  g0648(.A1(new_n791), .A2(new_n824), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR4_X1   g0649(.A1(new_n843), .A2(new_n844), .A3(new_n846), .A4(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n796), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n479), .B2(new_n851), .C1(new_n523), .C2(new_n789), .ZN(new_n852));
  INV_X1    g0652(.A(G132), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n254), .B1(new_n801), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n810), .A2(new_n202), .ZN(new_n855));
  INV_X1    g0655(.A(new_n809), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(G50), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT102), .Z(new_n858));
  INV_X1    g0658(.A(new_n804), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n854), .B(new_n858), .C1(G58), .C2(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G137), .A2(new_n790), .B1(new_n806), .B2(G150), .ZN(new_n861));
  INV_X1    g0661(.A(G143), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n861), .B1(new_n862), .B2(new_n789), .C1(new_n851), .C2(new_n339), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT101), .Z(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT34), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n864), .A2(KEYINPUT34), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n852), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n842), .B1(new_n868), .B2(new_n783), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT103), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n451), .A2(new_n707), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n463), .B1(new_n466), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n464), .A2(new_n707), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n869), .A2(new_n870), .B1(new_n778), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n870), .B2(new_n869), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT104), .Z(new_n877));
  NAND2_X1  g0677(.A1(new_n693), .A2(new_n707), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n874), .ZN(new_n879));
  INV_X1    g0679(.A(new_n874), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n693), .A2(new_n707), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n765), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT105), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n765), .A2(new_n879), .A3(new_n881), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n884), .A2(new_n828), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n877), .A2(new_n887), .ZN(G384));
  AND2_X1   g0688(.A1(new_n608), .A2(KEYINPUT35), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n608), .A2(KEYINPUT35), .ZN(new_n890));
  NOR4_X1   g0690(.A1(new_n889), .A2(new_n890), .A3(new_n479), .A4(new_n227), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT36), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n206), .A2(G50), .A3(G77), .A4(new_n336), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n269), .B(G13), .C1(new_n893), .C2(new_n244), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n695), .A2(new_n706), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n335), .B1(new_n346), .B2(new_n364), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n334), .B1(new_n898), .B2(new_n366), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n398), .B1(new_n899), .B2(new_n704), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n377), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT37), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n704), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n388), .B1(new_n376), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(KEYINPUT107), .B(KEYINPUT37), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(new_n398), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n378), .A2(new_n400), .A3(new_n390), .A4(new_n402), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n899), .A2(new_n704), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n907), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT108), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n907), .B2(new_n910), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n907), .A2(new_n910), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT38), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(KEYINPUT108), .A3(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT39), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n908), .A2(new_n388), .A3(new_n903), .ZN(new_n921));
  INV_X1    g0721(.A(new_n905), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n904), .A2(KEYINPUT109), .A3(new_n398), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT109), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n905), .B1(new_n904), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n398), .B2(new_n904), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n917), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT39), .B1(new_n928), .B2(new_n911), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT110), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n920), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n916), .A2(new_n917), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n912), .A3(new_n911), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n935), .B2(new_n918), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT110), .B1(new_n936), .B2(new_n929), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n897), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n319), .A2(new_n311), .A3(new_n321), .A4(new_n323), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n310), .A2(new_n707), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT106), .ZN(new_n942));
  INV_X1    g0742(.A(new_n940), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n941), .A2(new_n942), .B1(new_n325), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n939), .A2(new_n940), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(KEYINPUT106), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n881), .B2(new_n873), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n915), .A2(new_n919), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n949), .A2(new_n950), .B1(new_n391), .B2(new_n704), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n938), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n699), .B1(new_n743), .B2(new_n472), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n874), .B1(new_n944), .B2(new_n946), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n935), .A2(new_n763), .A3(new_n956), .A4(new_n918), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT40), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n956), .A2(new_n763), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n958), .B1(new_n928), .B2(new_n911), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n957), .A2(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n961), .A2(new_n472), .A3(new_n763), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n961), .B1(new_n472), .B2(new_n763), .ZN(new_n963));
  OR3_X1    g0763(.A1(new_n962), .A2(new_n963), .A3(new_n714), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n955), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n269), .B2(new_n773), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n955), .A2(new_n964), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n895), .B1(new_n966), .B2(new_n967), .ZN(G367));
  NAND3_X1  g0768(.A1(new_n575), .A2(new_n579), .A3(new_n706), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n579), .A2(new_n706), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n970), .B1(new_n672), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT43), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n615), .A2(new_n626), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n613), .A2(new_n707), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n681), .B2(new_n706), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n724), .A2(new_n978), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(KEYINPUT42), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n716), .A2(new_n615), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n706), .B1(new_n981), .B2(new_n626), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n979), .B2(KEYINPUT42), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n974), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n972), .A2(new_n973), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n984), .A2(new_n985), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n721), .A2(new_n978), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n727), .B(new_n992), .Z(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n724), .B1(new_n720), .B2(new_n723), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n770), .A2(new_n771), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n715), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n997), .B2(new_n995), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n999), .A2(new_n766), .A3(KEYINPUT112), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n978), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n722), .B2(new_n724), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT44), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n724), .A2(new_n722), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1004), .A2(new_n978), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT45), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(new_n721), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT112), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n998), .B2(new_n767), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1000), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n994), .B1(new_n1011), .B2(new_n766), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n774), .B(KEYINPUT113), .Z(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n991), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n972), .A2(new_n780), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n836), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n726), .B2(new_n554), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n238), .A2(new_n833), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n828), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT46), .B1(new_n856), .B2(G116), .ZN(new_n1021));
  AND3_X1   g0821(.A1(new_n856), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(new_n645), .C2(new_n788), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n847), .A2(new_n523), .B1(new_n804), .B2(new_n454), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n348), .B1(new_n801), .B2(new_n817), .C1(new_n791), .C2(new_n845), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n810), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1024), .B(new_n1025), .C1(G97), .C2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1023), .B(new_n1027), .C1(new_n851), .C2(new_n848), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT114), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n201), .A2(new_n809), .B1(new_n810), .B2(new_n294), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n804), .A2(new_n202), .ZN(new_n1031));
  INV_X1    g0831(.A(G137), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n254), .B1(new_n801), .B2(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n791), .A2(new_n862), .B1(new_n847), .B2(new_n339), .ZN(new_n1034));
  NOR4_X1   g0834(.A1(new_n1030), .A2(new_n1031), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n243), .B2(new_n851), .C1(new_n407), .C2(new_n789), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1029), .A2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT47), .Z(new_n1038));
  OAI211_X1 g0838(.A(new_n1016), .B(new_n1020), .C1(new_n1038), .C2(new_n782), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1015), .A2(new_n1039), .ZN(G387));
  NAND3_X1  g0840(.A1(new_n717), .A2(new_n719), .A3(new_n780), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n729), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n830), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(G107), .B2(new_n218), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n235), .A2(G45), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT115), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n328), .A2(new_n243), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT50), .Z(new_n1048));
  AOI211_X1 g0848(.A(G45), .B(new_n1042), .C1(G68), .C2(G77), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n726), .B(new_n254), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1044), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n776), .B1(new_n1051), .B2(new_n1017), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT116), .Z(new_n1053));
  AOI22_X1  g0853(.A1(new_n796), .A2(G68), .B1(new_n328), .B2(new_n806), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT117), .Z(new_n1055));
  OAI22_X1  g0855(.A1(new_n294), .A2(new_n809), .B1(new_n810), .B2(new_n563), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n348), .B1(new_n821), .B2(G150), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n339), .B2(new_n791), .C1(new_n446), .C2(new_n804), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1056), .B(new_n1058), .C1(G50), .C2(new_n788), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G322), .A2(new_n790), .B1(new_n806), .B2(G311), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n817), .B2(new_n789), .C1(new_n851), .C2(new_n641), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1063), .A2(KEYINPUT48), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(KEYINPUT48), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n809), .A2(new_n523), .B1(new_n804), .B2(new_n848), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(KEYINPUT49), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n348), .B1(new_n813), .B2(new_n801), .C1(new_n810), .C2(new_n479), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT118), .Z(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1067), .A2(KEYINPUT49), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1060), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1053), .B1(new_n783), .B2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n999), .A2(new_n1014), .B1(new_n1041), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n999), .A2(new_n766), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n727), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n999), .A2(new_n766), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(G393));
  INV_X1    g0879(.A(new_n721), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1007), .B(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT119), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1013), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n728), .B1(new_n1081), .B2(new_n1076), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n1011), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n978), .A2(new_n780), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1017), .B1(G97), .B2(new_n726), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n242), .A2(new_n833), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n828), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n847), .A2(new_n641), .B1(new_n479), .B2(new_n804), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT120), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n254), .B1(new_n821), .B2(G322), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n809), .B2(new_n848), .C1(new_n454), .C2(new_n810), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1092), .B(new_n1094), .C1(G294), .C2(new_n796), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n788), .A2(G311), .B1(G317), .B2(new_n790), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT52), .Z(new_n1097));
  AOI22_X1  g0897(.A1(new_n788), .A2(G159), .B1(G150), .B2(new_n790), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT51), .Z(new_n1099));
  OAI22_X1  g0899(.A1(new_n202), .A2(new_n809), .B1(new_n810), .B2(new_n559), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n348), .B1(new_n821), .B2(G143), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1101), .B1(new_n243), .B2(new_n847), .C1(new_n294), .C2(new_n804), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1100), .B(new_n1102), .C1(new_n328), .C2(new_n796), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1095), .A2(new_n1097), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1087), .B(new_n1090), .C1(new_n782), .C2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1084), .A2(new_n1086), .A3(new_n1105), .ZN(G390));
  NAND2_X1  g0906(.A1(new_n765), .A2(new_n472), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n742), .A2(new_n872), .B1(new_n464), .B2(new_n707), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n763), .A2(G330), .A3(new_n880), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n948), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n763), .A2(G330), .A3(new_n880), .A4(new_n947), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1108), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1110), .A2(new_n1111), .B1(new_n873), .B2(new_n881), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n954), .B(new_n1107), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n881), .A2(new_n873), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n947), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n897), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n932), .A2(new_n937), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n896), .B1(new_n928), .B2(new_n911), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n1108), .B2(new_n948), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1118), .A2(new_n1120), .A3(new_n1111), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1111), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1114), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1111), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1118), .A2(new_n1120), .A3(new_n1111), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n954), .A2(new_n1107), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1113), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1108), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1126), .A2(new_n1127), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1123), .A2(new_n1132), .A3(new_n727), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n809), .A2(new_n559), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n348), .B1(new_n804), .B2(new_n294), .C1(new_n523), .C2(new_n801), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n791), .A2(new_n823), .B1(new_n847), .B2(new_n454), .ZN(new_n1136));
  NOR4_X1   g0936(.A1(new_n1134), .A2(new_n855), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1137), .B1(new_n563), .B2(new_n851), .C1(new_n479), .C2(new_n789), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT122), .Z(new_n1139));
  NAND2_X1  g0939(.A1(new_n1026), .A2(G50), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n859), .A2(G159), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n348), .B1(new_n821), .B2(G125), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(G128), .A2(new_n790), .B1(new_n806), .B2(G137), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT54), .B(G143), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n851), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(KEYINPUT53), .B1(new_n809), .B2(new_n407), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n853), .B2(new_n789), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n809), .A2(KEYINPUT53), .A3(new_n407), .ZN(new_n1149));
  NOR4_X1   g0949(.A1(new_n1144), .A2(new_n1146), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT121), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n783), .B1(new_n1139), .B2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1152), .B(new_n776), .C1(new_n328), .C2(new_n841), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n931), .B1(new_n920), .B2(new_n930), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n936), .A2(KEYINPUT110), .A3(new_n929), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1153), .B1(new_n1156), .B2(new_n778), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n1014), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT123), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1133), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1160), .B1(new_n1133), .B2(new_n1159), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(G378));
  XOR2_X1   g0963(.A(KEYINPUT124), .B(KEYINPUT56), .Z(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n442), .A2(new_n704), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT55), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n439), .A2(new_n444), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1167), .B1(new_n439), .B2(new_n444), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1165), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n439), .A2(new_n444), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1167), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(new_n1164), .A3(new_n1168), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT125), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1171), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n961), .B2(G330), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n957), .A2(new_n958), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n959), .A2(new_n960), .ZN(new_n1180));
  AND4_X1   g0980(.A1(G330), .A2(new_n1179), .A3(new_n1180), .A4(new_n1177), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n1178), .A2(new_n1181), .B1(new_n938), .B2(new_n952), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n896), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1179), .A2(G330), .A3(new_n1180), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1177), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n961), .A2(G330), .A3(new_n1177), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1183), .A2(new_n1186), .A3(new_n951), .A4(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1182), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1014), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1171), .A2(new_n1175), .A3(new_n778), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n776), .B1(new_n841), .B2(G50), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n201), .A2(new_n810), .B1(new_n809), .B2(new_n294), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n791), .A2(new_n479), .B1(new_n847), .B2(new_n563), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n512), .B(new_n348), .C1(new_n801), .C2(new_n823), .ZN(new_n1195));
  NOR4_X1   g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1031), .A4(new_n1195), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n454), .B2(new_n789), .C1(new_n446), .C2(new_n851), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT58), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(G50), .B1(new_n251), .B2(new_n512), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n254), .B2(G41), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n790), .A2(G125), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n407), .B2(new_n804), .C1(new_n853), .C2(new_n847), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n809), .A2(new_n1145), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(G128), .C2(new_n788), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1032), .B2(new_n851), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1026), .A2(G159), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G33), .B(G41), .C1(new_n821), .C2(G124), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1202), .B1(new_n1198), .B2(new_n1197), .C1(new_n1208), .C2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1192), .B1(new_n1213), .B2(new_n783), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1191), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1190), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT57), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1182), .B2(new_n1188), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1121), .A2(new_n1122), .A3(new_n1114), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1219), .B1(new_n1220), .B2(new_n1128), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n727), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1128), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1132), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT57), .B1(new_n1224), .B2(new_n1189), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1217), .B1(new_n1222), .B2(new_n1225), .ZN(G375));
  NAND2_X1  g1026(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n948), .A2(new_n778), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n776), .B1(new_n841), .B2(G68), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n348), .B1(new_n801), .B2(new_n824), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n791), .A2(new_n523), .B1(new_n847), .B2(new_n479), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n554), .C2(new_n859), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G77), .A2(new_n1026), .B1(new_n856), .B2(G97), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(new_n823), .C2(new_n789), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n851), .A2(new_n454), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G58), .A2(new_n1026), .B1(new_n856), .B2(G159), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n348), .B1(new_n821), .B2(G128), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n847), .B2(new_n1145), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n791), .A2(new_n853), .B1(new_n804), .B2(new_n243), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1236), .B(new_n1240), .C1(new_n1032), .C2(new_n789), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n851), .A2(new_n407), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n1234), .A2(new_n1235), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1229), .B1(new_n1243), .B2(new_n783), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1227), .A2(new_n1014), .B1(new_n1228), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1114), .A2(new_n993), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1227), .A2(new_n1223), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1245), .B1(new_n1246), .B2(new_n1247), .ZN(G381));
  OR2_X1    g1048(.A1(G384), .A2(G381), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(G390), .A2(new_n1249), .A3(G396), .A4(G393), .ZN(new_n1250));
  INV_X1    g1050(.A(G387), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1133), .A2(new_n1159), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1225), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n728), .B1(new_n1224), .B2(new_n1219), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1216), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1250), .A2(new_n1251), .A3(new_n1253), .A4(new_n1256), .ZN(G407));
  NAND2_X1  g1057(.A1(new_n705), .A2(G213), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1256), .A2(new_n1253), .A3(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(G407), .A2(new_n1260), .A3(G213), .ZN(G409));
  NAND2_X1  g1061(.A1(new_n1189), .A2(KEYINPUT126), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT126), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1182), .A2(new_n1188), .A3(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(new_n1014), .A3(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n993), .B(new_n1189), .C1(new_n1220), .C2(new_n1128), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(new_n1215), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1253), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1252), .A2(KEYINPUT123), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1133), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1268), .B1(new_n1271), .B2(G375), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1247), .B1(KEYINPUT60), .B2(new_n1114), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1128), .A2(new_n1129), .A3(KEYINPUT60), .A4(new_n1130), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n727), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1245), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n877), .A3(new_n887), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G384), .B(new_n1245), .C1(new_n1273), .C2(new_n1275), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1272), .A2(new_n1258), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT62), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT61), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1259), .A2(G2897), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1277), .A2(new_n1278), .A3(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1284), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1256), .A2(G378), .B1(new_n1253), .B2(new_n1267), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1287), .B1(new_n1288), .B2(new_n1259), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT62), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1272), .A2(new_n1290), .A3(new_n1258), .A4(new_n1280), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1282), .A2(new_n1283), .A3(new_n1289), .A4(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(G390), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G387), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1015), .A2(G390), .A3(new_n1039), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(G393), .B(G396), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G390), .B1(new_n1015), .B2(new_n1039), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT127), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1297), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1294), .A2(new_n1297), .A3(new_n1295), .A4(new_n1299), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1292), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1272), .A2(new_n1258), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT61), .B1(new_n1305), .B2(new_n1287), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT63), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1281), .A2(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1272), .A2(KEYINPUT63), .A3(new_n1258), .A4(new_n1280), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1306), .A2(new_n1307), .A3(new_n1309), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1304), .A2(new_n1311), .ZN(G405));
  NAND2_X1  g1112(.A1(new_n1256), .A2(G378), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G375), .A2(new_n1253), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1280), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1313), .A2(new_n1279), .A3(new_n1314), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1303), .B(new_n1318), .ZN(G402));
endmodule


